
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire _43812_;
  wire _43813_;
  wire _43814_;
  wire _43815_;
  wire _43816_;
  wire _43817_;
  wire _43818_;
  wire _43819_;
  wire _43820_;
  wire _43821_;
  wire _43822_;
  wire _43823_;
  wire _43824_;
  wire _43825_;
  wire _43826_;
  wire _43827_;
  wire _43828_;
  wire _43829_;
  wire _43830_;
  wire _43831_;
  wire _43832_;
  wire _43833_;
  wire _43834_;
  wire _43835_;
  wire _43836_;
  wire _43837_;
  wire _43838_;
  wire _43839_;
  wire _43840_;
  wire _43841_;
  wire _43842_;
  wire _43843_;
  wire _43844_;
  wire _43845_;
  wire _43846_;
  wire _43847_;
  wire _43848_;
  wire _43849_;
  wire _43850_;
  wire _43851_;
  wire _43852_;
  wire _43853_;
  wire _43854_;
  wire _43855_;
  wire _43856_;
  wire _43857_;
  wire _43858_;
  wire _43859_;
  wire _43860_;
  wire _43861_;
  wire _43862_;
  wire _43863_;
  wire _43864_;
  wire _43865_;
  wire _43866_;
  wire _43867_;
  wire _43868_;
  wire _43869_;
  wire _43870_;
  wire _43871_;
  wire _43872_;
  wire _43873_;
  wire _43874_;
  wire _43875_;
  wire _43876_;
  wire _43877_;
  wire _43878_;
  wire _43879_;
  wire _43880_;
  wire _43881_;
  wire _43882_;
  wire _43883_;
  wire _43884_;
  wire _43885_;
  wire _43886_;
  wire _43887_;
  wire _43888_;
  wire _43889_;
  wire _43890_;
  wire _43891_;
  wire _43892_;
  wire _43893_;
  wire _43894_;
  wire _43895_;
  wire _43896_;
  wire _43897_;
  wire _43898_;
  wire _43899_;
  wire _43900_;
  wire _43901_;
  wire _43902_;
  wire _43903_;
  wire _43904_;
  wire _43905_;
  wire _43906_;
  wire _43907_;
  wire _43908_;
  wire _43909_;
  wire _43910_;
  wire _43911_;
  wire _43912_;
  wire _43913_;
  wire _43914_;
  wire _43915_;
  wire _43916_;
  wire _43917_;
  wire _43918_;
  wire _43919_;
  wire _43920_;
  wire _43921_;
  wire _43922_;
  wire _43923_;
  wire _43924_;
  wire _43925_;
  wire _43926_;
  wire _43927_;
  wire _43928_;
  wire _43929_;
  wire _43930_;
  wire _43931_;
  wire _43932_;
  wire _43933_;
  wire _43934_;
  wire _43935_;
  wire _43936_;
  wire _43937_;
  wire _43938_;
  wire _43939_;
  wire _43940_;
  wire _43941_;
  wire _43942_;
  wire _43943_;
  wire _43944_;
  wire _43945_;
  wire _43946_;
  wire _43947_;
  wire _43948_;
  wire _43949_;
  wire _43950_;
  wire _43951_;
  wire _43952_;
  wire _43953_;
  wire _43954_;
  wire _43955_;
  wire _43956_;
  wire _43957_;
  wire _43958_;
  wire _43959_;
  wire _43960_;
  wire _43961_;
  wire _43962_;
  wire _43963_;
  wire _43964_;
  wire _43965_;
  wire _43966_;
  wire _43967_;
  wire _43968_;
  wire _43969_;
  wire _43970_;
  wire _43971_;
  wire _43972_;
  wire _43973_;
  wire _43974_;
  wire _43975_;
  wire _43976_;
  wire _43977_;
  wire _43978_;
  wire _43979_;
  wire _43980_;
  wire _43981_;
  wire _43982_;
  wire _43983_;
  wire _43984_;
  wire _43985_;
  wire _43986_;
  wire _43987_;
  wire _43988_;
  wire _43989_;
  wire _43990_;
  wire _43991_;
  wire _43992_;
  wire _43993_;
  wire _43994_;
  wire _43995_;
  wire _43996_;
  wire _43997_;
  wire _43998_;
  wire _43999_;
  wire _44000_;
  wire _44001_;
  wire _44002_;
  wire _44003_;
  wire _44004_;
  wire _44005_;
  wire _44006_;
  wire [7:0] ACC_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] PCON_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [7:0] ie_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [6:0] \oc8051_golden_model_1.n0988 ;
  wire \oc8051_golden_model_1.n0989 ;
  wire \oc8051_golden_model_1.n0990 ;
  wire \oc8051_golden_model_1.n0991 ;
  wire \oc8051_golden_model_1.n0992 ;
  wire \oc8051_golden_model_1.n0993 ;
  wire \oc8051_golden_model_1.n0994 ;
  wire \oc8051_golden_model_1.n0995 ;
  wire \oc8051_golden_model_1.n0996 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire [7:0] \oc8051_golden_model_1.n1004 ;
  wire [7:0] \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire \oc8051_golden_model_1.n1018 ;
  wire \oc8051_golden_model_1.n1019 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire [7:0] \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1043 ;
  wire [7:0] \oc8051_golden_model_1.n1044 ;
  wire [3:0] \oc8051_golden_model_1.n1137 ;
  wire [3:0] \oc8051_golden_model_1.n1139 ;
  wire [3:0] \oc8051_golden_model_1.n1141 ;
  wire [3:0] \oc8051_golden_model_1.n1142 ;
  wire [3:0] \oc8051_golden_model_1.n1143 ;
  wire [3:0] \oc8051_golden_model_1.n1144 ;
  wire [3:0] \oc8051_golden_model_1.n1145 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1147 ;
  wire \oc8051_golden_model_1.n1194 ;
  wire \oc8051_golden_model_1.n1239 ;
  wire [8:0] \oc8051_golden_model_1.n1240 ;
  wire [8:0] \oc8051_golden_model_1.n1241 ;
  wire [7:0] \oc8051_golden_model_1.n1242 ;
  wire \oc8051_golden_model_1.n1243 ;
  wire [2:0] \oc8051_golden_model_1.n1244 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [1:0] \oc8051_golden_model_1.n1246 ;
  wire [7:0] \oc8051_golden_model_1.n1247 ;
  wire [6:0] \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1251 ;
  wire \oc8051_golden_model_1.n1252 ;
  wire \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1255 ;
  wire \oc8051_golden_model_1.n1256 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [7:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1280 ;
  wire [7:0] \oc8051_golden_model_1.n1281 ;
  wire [15:0] \oc8051_golden_model_1.n1323 ;
  wire [7:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire \oc8051_golden_model_1.n1328 ;
  wire \oc8051_golden_model_1.n1329 ;
  wire \oc8051_golden_model_1.n1330 ;
  wire \oc8051_golden_model_1.n1331 ;
  wire \oc8051_golden_model_1.n1332 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire \oc8051_golden_model_1.n1340 ;
  wire [7:0] \oc8051_golden_model_1.n1341 ;
  wire [8:0] \oc8051_golden_model_1.n1343 ;
  wire [8:0] \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire [3:0] \oc8051_golden_model_1.n1349 ;
  wire [4:0] \oc8051_golden_model_1.n1350 ;
  wire [4:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [8:0] \oc8051_golden_model_1.n1356 ;
  wire \oc8051_golden_model_1.n1364 ;
  wire [7:0] \oc8051_golden_model_1.n1365 ;
  wire [6:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1381 ;
  wire [7:0] \oc8051_golden_model_1.n1382 ;
  wire [8:0] \oc8051_golden_model_1.n1404 ;
  wire \oc8051_golden_model_1.n1405 ;
  wire [4:0] \oc8051_golden_model_1.n1410 ;
  wire \oc8051_golden_model_1.n1411 ;
  wire \oc8051_golden_model_1.n1419 ;
  wire [7:0] \oc8051_golden_model_1.n1420 ;
  wire [6:0] \oc8051_golden_model_1.n1421 ;
  wire \oc8051_golden_model_1.n1436 ;
  wire [7:0] \oc8051_golden_model_1.n1437 ;
  wire [8:0] \oc8051_golden_model_1.n1439 ;
  wire [8:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1442 ;
  wire [3:0] \oc8051_golden_model_1.n1443 ;
  wire [4:0] \oc8051_golden_model_1.n1444 ;
  wire [4:0] \oc8051_golden_model_1.n1446 ;
  wire \oc8051_golden_model_1.n1447 ;
  wire [8:0] \oc8051_golden_model_1.n1448 ;
  wire \oc8051_golden_model_1.n1455 ;
  wire [7:0] \oc8051_golden_model_1.n1456 ;
  wire [6:0] \oc8051_golden_model_1.n1457 ;
  wire \oc8051_golden_model_1.n1472 ;
  wire [7:0] \oc8051_golden_model_1.n1473 ;
  wire [8:0] \oc8051_golden_model_1.n1476 ;
  wire \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1484 ;
  wire [7:0] \oc8051_golden_model_1.n1485 ;
  wire [6:0] \oc8051_golden_model_1.n1486 ;
  wire [7:0] \oc8051_golden_model_1.n1487 ;
  wire [8:0] \oc8051_golden_model_1.n1489 ;
  wire [8:0] \oc8051_golden_model_1.n1491 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [4:0] \oc8051_golden_model_1.n1493 ;
  wire [4:0] \oc8051_golden_model_1.n1495 ;
  wire \oc8051_golden_model_1.n1496 ;
  wire [8:0] \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire [4:0] \oc8051_golden_model_1.n1524 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire [7:0] \oc8051_golden_model_1.n1526 ;
  wire [6:0] \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [8:0] \oc8051_golden_model_1.n1530 ;
  wire \oc8051_golden_model_1.n1531 ;
  wire \oc8051_golden_model_1.n1538 ;
  wire [7:0] \oc8051_golden_model_1.n1539 ;
  wire [6:0] \oc8051_golden_model_1.n1540 ;
  wire [7:0] \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [6:0] \oc8051_golden_model_1.n1543 ;
  wire [7:0] \oc8051_golden_model_1.n1544 ;
  wire [8:0] \oc8051_golden_model_1.n1547 ;
  wire [8:0] \oc8051_golden_model_1.n1548 ;
  wire [7:0] \oc8051_golden_model_1.n1549 ;
  wire [7:0] \oc8051_golden_model_1.n1550 ;
  wire [6:0] \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1552 ;
  wire \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire \oc8051_golden_model_1.n1555 ;
  wire \oc8051_golden_model_1.n1556 ;
  wire \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire \oc8051_golden_model_1.n1559 ;
  wire \oc8051_golden_model_1.n1566 ;
  wire [7:0] \oc8051_golden_model_1.n1567 ;
  wire [7:0] \oc8051_golden_model_1.n1568 ;
  wire [8:0] \oc8051_golden_model_1.n1571 ;
  wire [8:0] \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire [4:0] \oc8051_golden_model_1.n1575 ;
  wire [4:0] \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1585 ;
  wire [7:0] \oc8051_golden_model_1.n1586 ;
  wire [6:0] \oc8051_golden_model_1.n1587 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [7:0] \oc8051_golden_model_1.n1603 ;
  wire [8:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1608 ;
  wire [4:0] \oc8051_golden_model_1.n1610 ;
  wire \oc8051_golden_model_1.n1611 ;
  wire \oc8051_golden_model_1.n1618 ;
  wire [7:0] \oc8051_golden_model_1.n1619 ;
  wire [6:0] \oc8051_golden_model_1.n1620 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [7:0] \oc8051_golden_model_1.n1636 ;
  wire [8:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1641 ;
  wire [4:0] \oc8051_golden_model_1.n1643 ;
  wire \oc8051_golden_model_1.n1644 ;
  wire \oc8051_golden_model_1.n1651 ;
  wire [7:0] \oc8051_golden_model_1.n1652 ;
  wire [6:0] \oc8051_golden_model_1.n1653 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [7:0] \oc8051_golden_model_1.n1669 ;
  wire [8:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1674 ;
  wire [4:0] \oc8051_golden_model_1.n1676 ;
  wire \oc8051_golden_model_1.n1677 ;
  wire \oc8051_golden_model_1.n1684 ;
  wire [7:0] \oc8051_golden_model_1.n1685 ;
  wire [6:0] \oc8051_golden_model_1.n1686 ;
  wire \oc8051_golden_model_1.n1701 ;
  wire [7:0] \oc8051_golden_model_1.n1702 ;
  wire [7:0] \oc8051_golden_model_1.n1727 ;
  wire [6:0] \oc8051_golden_model_1.n1728 ;
  wire [7:0] \oc8051_golden_model_1.n1729 ;
  wire \oc8051_golden_model_1.n1784 ;
  wire [7:0] \oc8051_golden_model_1.n1785 ;
  wire \oc8051_golden_model_1.n1801 ;
  wire [7:0] \oc8051_golden_model_1.n1802 ;
  wire \oc8051_golden_model_1.n1818 ;
  wire [7:0] \oc8051_golden_model_1.n1819 ;
  wire \oc8051_golden_model_1.n1835 ;
  wire [7:0] \oc8051_golden_model_1.n1836 ;
  wire [7:0] \oc8051_golden_model_1.n1859 ;
  wire [6:0] \oc8051_golden_model_1.n1860 ;
  wire [7:0] \oc8051_golden_model_1.n1861 ;
  wire \oc8051_golden_model_1.n1916 ;
  wire [7:0] \oc8051_golden_model_1.n1917 ;
  wire \oc8051_golden_model_1.n1933 ;
  wire [7:0] \oc8051_golden_model_1.n1934 ;
  wire \oc8051_golden_model_1.n1950 ;
  wire [7:0] \oc8051_golden_model_1.n1951 ;
  wire \oc8051_golden_model_1.n1967 ;
  wire [7:0] \oc8051_golden_model_1.n1968 ;
  wire \oc8051_golden_model_1.n2065 ;
  wire [7:0] \oc8051_golden_model_1.n2066 ;
  wire \oc8051_golden_model_1.n2082 ;
  wire [7:0] \oc8051_golden_model_1.n2083 ;
  wire \oc8051_golden_model_1.n2099 ;
  wire [7:0] \oc8051_golden_model_1.n2100 ;
  wire \oc8051_golden_model_1.n2116 ;
  wire [7:0] \oc8051_golden_model_1.n2117 ;
  wire \oc8051_golden_model_1.n2121 ;
  wire [6:0] \oc8051_golden_model_1.n2122 ;
  wire [7:0] \oc8051_golden_model_1.n2123 ;
  wire [6:0] \oc8051_golden_model_1.n2124 ;
  wire [7:0] \oc8051_golden_model_1.n2125 ;
  wire \oc8051_golden_model_1.n2140 ;
  wire [7:0] \oc8051_golden_model_1.n2141 ;
  wire \oc8051_golden_model_1.n2180 ;
  wire [7:0] \oc8051_golden_model_1.n2181 ;
  wire [6:0] \oc8051_golden_model_1.n2182 ;
  wire [7:0] \oc8051_golden_model_1.n2183 ;
  wire [3:0] \oc8051_golden_model_1.n2190 ;
  wire \oc8051_golden_model_1.n2191 ;
  wire [7:0] \oc8051_golden_model_1.n2192 ;
  wire [6:0] \oc8051_golden_model_1.n2193 ;
  wire \oc8051_golden_model_1.n2208 ;
  wire [7:0] \oc8051_golden_model_1.n2209 ;
  wire [7:0] \oc8051_golden_model_1.n2421 ;
  wire \oc8051_golden_model_1.n2424 ;
  wire \oc8051_golden_model_1.n2426 ;
  wire \oc8051_golden_model_1.n2432 ;
  wire [7:0] \oc8051_golden_model_1.n2433 ;
  wire [6:0] \oc8051_golden_model_1.n2434 ;
  wire \oc8051_golden_model_1.n2449 ;
  wire [7:0] \oc8051_golden_model_1.n2450 ;
  wire \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2456 ;
  wire \oc8051_golden_model_1.n2462 ;
  wire [7:0] \oc8051_golden_model_1.n2463 ;
  wire [6:0] \oc8051_golden_model_1.n2464 ;
  wire \oc8051_golden_model_1.n2479 ;
  wire [7:0] \oc8051_golden_model_1.n2480 ;
  wire \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2486 ;
  wire \oc8051_golden_model_1.n2492 ;
  wire [7:0] \oc8051_golden_model_1.n2493 ;
  wire [6:0] \oc8051_golden_model_1.n2494 ;
  wire \oc8051_golden_model_1.n2509 ;
  wire [7:0] \oc8051_golden_model_1.n2510 ;
  wire \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2516 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire [7:0] \oc8051_golden_model_1.n2523 ;
  wire [6:0] \oc8051_golden_model_1.n2524 ;
  wire \oc8051_golden_model_1.n2539 ;
  wire [7:0] \oc8051_golden_model_1.n2540 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire [7:0] \oc8051_golden_model_1.n2545 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire [7:0] \oc8051_golden_model_1.n2548 ;
  wire [15:0] \oc8051_golden_model_1.n2552 ;
  wire \oc8051_golden_model_1.n2558 ;
  wire [7:0] \oc8051_golden_model_1.n2559 ;
  wire [6:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2575 ;
  wire [7:0] \oc8051_golden_model_1.n2576 ;
  wire \oc8051_golden_model_1.n2579 ;
  wire [7:0] \oc8051_golden_model_1.n2580 ;
  wire [6:0] \oc8051_golden_model_1.n2581 ;
  wire [7:0] \oc8051_golden_model_1.n2582 ;
  wire \oc8051_golden_model_1.n2614 ;
  wire [7:0] \oc8051_golden_model_1.n2615 ;
  wire [6:0] \oc8051_golden_model_1.n2616 ;
  wire [7:0] \oc8051_golden_model_1.n2617 ;
  wire \oc8051_golden_model_1.n2622 ;
  wire [7:0] \oc8051_golden_model_1.n2623 ;
  wire [6:0] \oc8051_golden_model_1.n2624 ;
  wire [7:0] \oc8051_golden_model_1.n2625 ;
  wire \oc8051_golden_model_1.n2630 ;
  wire [7:0] \oc8051_golden_model_1.n2631 ;
  wire [6:0] \oc8051_golden_model_1.n2632 ;
  wire [7:0] \oc8051_golden_model_1.n2633 ;
  wire \oc8051_golden_model_1.n2638 ;
  wire [7:0] \oc8051_golden_model_1.n2639 ;
  wire [6:0] \oc8051_golden_model_1.n2640 ;
  wire [7:0] \oc8051_golden_model_1.n2641 ;
  wire \oc8051_golden_model_1.n2646 ;
  wire [7:0] \oc8051_golden_model_1.n2647 ;
  wire [6:0] \oc8051_golden_model_1.n2648 ;
  wire [7:0] \oc8051_golden_model_1.n2649 ;
  wire [7:0] \oc8051_golden_model_1.n2674 ;
  wire [6:0] \oc8051_golden_model_1.n2675 ;
  wire [7:0] \oc8051_golden_model_1.n2676 ;
  wire [3:0] \oc8051_golden_model_1.n2677 ;
  wire [7:0] \oc8051_golden_model_1.n2678 ;
  wire \oc8051_golden_model_1.n2679 ;
  wire \oc8051_golden_model_1.n2680 ;
  wire \oc8051_golden_model_1.n2681 ;
  wire \oc8051_golden_model_1.n2682 ;
  wire \oc8051_golden_model_1.n2683 ;
  wire \oc8051_golden_model_1.n2684 ;
  wire \oc8051_golden_model_1.n2685 ;
  wire \oc8051_golden_model_1.n2686 ;
  wire \oc8051_golden_model_1.n2693 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [6:0] \oc8051_golden_model_1.n2715 ;
  wire [7:0] \oc8051_golden_model_1.n2731 ;
  wire \oc8051_golden_model_1.n2732 ;
  wire \oc8051_golden_model_1.n2733 ;
  wire \oc8051_golden_model_1.n2734 ;
  wire \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2736 ;
  wire \oc8051_golden_model_1.n2737 ;
  wire \oc8051_golden_model_1.n2738 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire \oc8051_golden_model_1.n2746 ;
  wire [7:0] \oc8051_golden_model_1.n2747 ;
  wire \oc8051_golden_model_1.n2748 ;
  wire \oc8051_golden_model_1.n2749 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2762 ;
  wire [7:0] \oc8051_golden_model_1.n2763 ;
  wire [7:0] \oc8051_golden_model_1.n2795 ;
  wire [6:0] \oc8051_golden_model_1.n2796 ;
  wire [7:0] \oc8051_golden_model_1.n2797 ;
  wire \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire [6:0] \oc8051_golden_model_1.n2818 ;
  wire \oc8051_golden_model_1.n2833 ;
  wire [7:0] \oc8051_golden_model_1.n2834 ;
  wire [7:0] \oc8051_golden_model_1.n2838 ;
  wire [3:0] \oc8051_golden_model_1.n2839 ;
  wire [7:0] \oc8051_golden_model_1.n2840 ;
  wire \oc8051_golden_model_1.n2841 ;
  wire \oc8051_golden_model_1.n2842 ;
  wire \oc8051_golden_model_1.n2843 ;
  wire \oc8051_golden_model_1.n2844 ;
  wire \oc8051_golden_model_1.n2845 ;
  wire \oc8051_golden_model_1.n2846 ;
  wire \oc8051_golden_model_1.n2847 ;
  wire \oc8051_golden_model_1.n2848 ;
  wire \oc8051_golden_model_1.n2855 ;
  wire [7:0] \oc8051_golden_model_1.n2856 ;
  wire \oc8051_golden_model_1.n2874 ;
  wire [7:0] \oc8051_golden_model_1.n2875 ;
  wire \oc8051_golden_model_1.n2891 ;
  wire [7:0] \oc8051_golden_model_1.n2892 ;
  wire [7:0] \oc8051_golden_model_1.n2893 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not _44007_ (_41755_, rst);
  not _44008_ (_15496_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _44009_ (_15507_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _44010_ (_15518_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15507_);
  and _44011_ (_15529_, _15518_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44012_ (_15540_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15507_);
  and _44013_ (_15551_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15507_);
  nor _44014_ (_15562_, _15551_, _15540_);
  and _44015_ (_15573_, _15562_, _15529_);
  nor _44016_ (_15584_, _15573_, _15496_);
  and _44017_ (_15595_, _15496_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44018_ (_15606_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _44019_ (_15617_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15606_);
  nor _44020_ (_15628_, _15617_, _15595_);
  not _44021_ (_15639_, _15628_);
  and _44022_ (_15650_, _15639_, _15573_);
  or _44023_ (_15661_, _15650_, _15584_);
  and _44024_ (_22440_, _15661_, _41755_);
  nor _44025_ (_15682_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _44026_ (_15693_, _15682_);
  and _44027_ (_15704_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _44028_ (_15715_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _44029_ (_15725_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _44030_ (_15736_, _15725_);
  not _44031_ (_15747_, _15617_);
  nor _44032_ (_15758_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _44033_ (_15769_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _44034_ (_15780_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15769_);
  nor _44035_ (_15791_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not _44036_ (_15802_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _44037_ (_15813_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15802_);
  nor _44038_ (_15824_, _15813_, _15791_);
  nor _44039_ (_15835_, _15824_, _15780_);
  not _44040_ (_15846_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _44041_ (_15857_, _15780_, _15846_);
  nor _44042_ (_15868_, _15857_, _15835_);
  and _44043_ (_15879_, _15868_, _15758_);
  not _44044_ (_15890_, _15879_);
  and _44045_ (_15901_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44046_ (_15912_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _44047_ (_15923_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _44048_ (_15934_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _15923_);
  and _44049_ (_15945_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _44050_ (_15956_, _15945_, _15912_);
  and _44051_ (_15967_, _15956_, _15890_);
  nor _44052_ (_15978_, _15967_, _15747_);
  not _44053_ (_15989_, _15595_);
  nor _44054_ (_16000_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _44055_ (_16011_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15802_);
  nor _44056_ (_16022_, _16011_, _16000_);
  nor _44057_ (_16033_, _16022_, _15780_);
  not _44058_ (_16044_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _44059_ (_16055_, _15780_, _16044_);
  nor _44060_ (_16065_, _16055_, _16033_);
  and _44061_ (_16076_, _16065_, _15758_);
  not _44062_ (_16087_, _16076_);
  and _44063_ (_16098_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _44064_ (_16109_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _44065_ (_16120_, _16109_, _16098_);
  and _44066_ (_16131_, _16120_, _16087_);
  nor _44067_ (_16142_, _16131_, _15989_);
  nor _44068_ (_16153_, _16142_, _15978_);
  nor _44069_ (_16164_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _44070_ (_16175_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15802_);
  nor _44071_ (_16186_, _16175_, _16164_);
  nor _44072_ (_16197_, _16186_, _15780_);
  not _44073_ (_16208_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _44074_ (_16219_, _15780_, _16208_);
  nor _44075_ (_16230_, _16219_, _16197_);
  and _44076_ (_16241_, _16230_, _15758_);
  not _44077_ (_16252_, _16241_);
  and _44078_ (_16263_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _44079_ (_16274_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44080_ (_16285_, _16274_, _16263_);
  and _44081_ (_16296_, _16285_, _16252_);
  nor _44082_ (_16307_, _16296_, _15639_);
  nor _44083_ (_16318_, _16307_, _15682_);
  and _44084_ (_16329_, _16318_, _16153_);
  nor _44085_ (_16340_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor _44086_ (_16351_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15802_);
  nor _44087_ (_16362_, _16351_, _16340_);
  nor _44088_ (_16373_, _16362_, _15780_);
  not _44089_ (_16384_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _44090_ (_16394_, _15780_, _16384_);
  nor _44091_ (_16405_, _16394_, _16373_);
  and _44092_ (_16416_, _16405_, _15758_);
  not _44093_ (_16427_, _16416_);
  and _44094_ (_16438_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _44095_ (_16449_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _44096_ (_16460_, _16449_, _16438_);
  and _44097_ (_16471_, _16460_, _16427_);
  and _44098_ (_16482_, _16471_, _15682_);
  nor _44099_ (_16493_, _16482_, _16329_);
  not _44100_ (_16504_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44101_ (_16515_, _16504_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44102_ (_16526_, _16515_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44103_ (_16537_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _44104_ (_16548_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44105_ (_16570_, _16548_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44106_ (_16571_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _44107_ (_16582_, _16571_, _16537_);
  not _44108_ (_16593_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44109_ (_16604_, _16515_, _16593_);
  and _44110_ (_16615_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _44111_ (_16626_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44112_ (_16637_, _16626_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _44113_ (_16648_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor _44114_ (_16659_, _16648_, _16615_);
  and _44115_ (_16670_, _16659_, _16582_);
  and _44116_ (_16681_, _16548_, _16593_);
  and _44117_ (_16692_, _16681_, _16405_);
  and _44118_ (_16703_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _44119_ (_16714_, _16703_, _16593_);
  and _44120_ (_16725_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _44121_ (_16736_, _16703_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _44122_ (_16746_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _44123_ (_16757_, _16746_, _16725_);
  not _44124_ (_16768_, _16757_);
  nor _44125_ (_16779_, _16768_, _16692_);
  and _44126_ (_16790_, _16779_, _16670_);
  not _44127_ (_16801_, _16790_);
  and _44128_ (_16812_, _16801_, _16493_);
  not _44129_ (_16823_, _16812_);
  nor _44130_ (_16834_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _44131_ (_16845_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15802_);
  nor _44132_ (_16856_, _16845_, _16834_);
  nor _44133_ (_16867_, _16856_, _15780_);
  not _44134_ (_16878_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _44135_ (_16889_, _15780_, _16878_);
  nor _44136_ (_16900_, _16889_, _16867_);
  and _44137_ (_16911_, _16900_, _15758_);
  not _44138_ (_16922_, _16911_);
  and _44139_ (_16933_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _44140_ (_16944_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _44141_ (_16955_, _16944_, _16933_);
  and _44142_ (_16966_, _16955_, _16922_);
  nor _44143_ (_16977_, _16966_, _15747_);
  nor _44144_ (_16988_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor _44145_ (_16999_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15802_);
  nor _44146_ (_17010_, _16999_, _16988_);
  nor _44147_ (_17021_, _17010_, _15780_);
  not _44148_ (_17032_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _44149_ (_17043_, _15780_, _17032_);
  nor _44150_ (_17054_, _17043_, _17021_);
  and _44151_ (_17065_, _17054_, _15758_);
  not _44152_ (_17075_, _17065_);
  and _44153_ (_17086_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _44154_ (_17097_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44155_ (_17108_, _17097_, _17086_);
  and _44156_ (_17119_, _17108_, _17075_);
  nor _44157_ (_17130_, _17119_, _15989_);
  nor _44158_ (_17141_, _17130_, _16977_);
  nor _44159_ (_17152_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _44160_ (_17162_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15802_);
  nor _44161_ (_17173_, _17162_, _17152_);
  nor _44162_ (_17184_, _17173_, _15780_);
  not _44163_ (_17195_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _44164_ (_17206_, _15780_, _17195_);
  nor _44165_ (_17217_, _17206_, _17184_);
  and _44166_ (_17228_, _17217_, _15758_);
  not _44167_ (_17239_, _17228_);
  and _44168_ (_17250_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _44169_ (_17260_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44170_ (_17271_, _17260_, _17250_);
  and _44171_ (_17292_, _17271_, _17239_);
  nor _44172_ (_17293_, _17292_, _15639_);
  nor _44173_ (_17314_, _17293_, _15682_);
  and _44174_ (_17315_, _17314_, _17141_);
  nor _44175_ (_17326_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor _44176_ (_17337_, _15802_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor _44177_ (_17347_, _17337_, _17326_);
  nor _44178_ (_17358_, _17347_, _15780_);
  not _44179_ (_17369_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _44180_ (_17380_, _15780_, _17369_);
  nor _44181_ (_17391_, _17380_, _17358_);
  and _44182_ (_17402_, _17391_, _15758_);
  not _44183_ (_17413_, _17402_);
  and _44184_ (_17424_, _15901_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _44185_ (_17434_, _15934_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _44186_ (_17445_, _17434_, _17424_);
  and _44187_ (_17456_, _17445_, _17413_);
  and _44188_ (_17467_, _17456_, _15682_);
  nor _44189_ (_17478_, _17467_, _17315_);
  and _44190_ (_17489_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _44191_ (_17500_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _44192_ (_17511_, _17500_, _17489_);
  and _44193_ (_17521_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _44194_ (_17532_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _44195_ (_17543_, _17532_, _17521_);
  and _44196_ (_17554_, _17543_, _17511_);
  and _44197_ (_17565_, _17391_, _16681_);
  and _44198_ (_17576_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _44199_ (_17587_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _44200_ (_17598_, _17587_, _17576_);
  not _44201_ (_17608_, _17598_);
  nor _44202_ (_17619_, _17608_, _17565_);
  and _44203_ (_17630_, _17619_, _17554_);
  not _44204_ (_17641_, _17630_);
  and _44205_ (_17652_, _17641_, _17478_);
  and _44206_ (_17663_, _17652_, _16823_);
  not _44207_ (_17674_, _17663_);
  and _44208_ (_17685_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _44209_ (_17696_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _44210_ (_17706_, _17696_, _17685_);
  and _44211_ (_17717_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _44212_ (_17728_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _44213_ (_17739_, _17728_, _17717_);
  and _44214_ (_17750_, _17739_, _17706_);
  and _44215_ (_17761_, _17054_, _16681_);
  and _44216_ (_17772_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _44217_ (_17783_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44218_ (_17794_, _17783_, _17772_);
  not _44219_ (_17804_, _17794_);
  nor _44220_ (_17815_, _17804_, _17761_);
  and _44221_ (_17826_, _17815_, _17750_);
  not _44222_ (_17837_, _17826_);
  and _44223_ (_17848_, _17837_, _17478_);
  and _44224_ (_17859_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _44225_ (_17870_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _44226_ (_17881_, _17870_, _17859_);
  and _44227_ (_17892_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _44228_ (_17903_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _44229_ (_17914_, _17903_, _17892_);
  and _44230_ (_17924_, _17914_, _17881_);
  and _44231_ (_17935_, _16681_, _16065_);
  and _44232_ (_17946_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _44233_ (_17957_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _44234_ (_17968_, _17957_, _17946_);
  not _44235_ (_17979_, _17968_);
  nor _44236_ (_17990_, _17979_, _17935_);
  and _44237_ (_18001_, _17990_, _17924_);
  not _44238_ (_18012_, _18001_);
  and _44239_ (_18023_, _18012_, _16493_);
  and _44240_ (_18034_, _17848_, _18023_);
  nor _44241_ (_18044_, _16812_, _18034_);
  and _44242_ (_18055_, _16801_, _18034_);
  nor _44243_ (_18066_, _18055_, _18044_);
  and _44244_ (_18077_, _18066_, _17848_);
  and _44245_ (_18088_, _17652_, _16812_);
  and _44246_ (_18099_, _16801_, _17478_);
  and _44247_ (_18110_, _17641_, _16493_);
  nor _44248_ (_18121_, _18110_, _18099_);
  nor _44249_ (_18132_, _18121_, _18088_);
  and _44250_ (_18143_, _18132_, _18077_);
  and _44251_ (_18153_, _18132_, _18055_);
  nor _44252_ (_18164_, _18153_, _18143_);
  nor _44253_ (_18175_, _18164_, _17674_);
  and _44254_ (_18186_, _17478_, _18012_);
  and _44255_ (_18197_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _44256_ (_18208_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _44257_ (_18219_, _18208_, _18197_);
  and _44258_ (_18230_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _44259_ (_18241_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _44260_ (_18252_, _18241_, _18230_);
  and _44261_ (_18263_, _18252_, _18219_);
  and _44262_ (_18273_, _16900_, _16681_);
  and _44263_ (_18284_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _44264_ (_18295_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _44265_ (_18306_, _18295_, _18284_);
  not _44266_ (_18317_, _18306_);
  nor _44267_ (_18328_, _18317_, _18273_);
  and _44268_ (_18339_, _18328_, _18263_);
  not _44269_ (_18350_, _18339_);
  and _44270_ (_18361_, _18350_, _16493_);
  and _44271_ (_18372_, _18361_, _18186_);
  and _44272_ (_18383_, _17837_, _16493_);
  nor _44273_ (_18393_, _18383_, _18186_);
  nor _44274_ (_18404_, _18393_, _18034_);
  and _44275_ (_18415_, _18404_, _18372_);
  nor _44276_ (_18426_, _16812_, _17848_);
  nor _44277_ (_18437_, _18426_, _18077_);
  and _44278_ (_18448_, _18437_, _18415_);
  nor _44279_ (_18459_, _18132_, _18077_);
  nor _44280_ (_18470_, _18459_, _18143_);
  nor _44281_ (_18481_, _18470_, _18055_);
  nor _44282_ (_18492_, _18481_, _18153_);
  and _44283_ (_18502_, _18492_, _18448_);
  nor _44284_ (_18513_, _18492_, _18448_);
  nor _44285_ (_18524_, _18513_, _18502_);
  not _44286_ (_18535_, _18524_);
  and _44287_ (_18546_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _44288_ (_18557_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _44289_ (_18568_, _18557_, _18546_);
  and _44290_ (_18579_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _44291_ (_18589_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _44292_ (_18600_, _18589_, _18579_);
  and _44293_ (_18611_, _18600_, _18568_);
  and _44294_ (_18622_, _17217_, _16681_);
  and _44295_ (_18633_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _44296_ (_18644_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44297_ (_18655_, _18644_, _18633_);
  not _44298_ (_18666_, _18655_);
  nor _44299_ (_18676_, _18666_, _18622_);
  and _44300_ (_18687_, _18676_, _18611_);
  not _44301_ (_18698_, _18687_);
  and _44302_ (_18709_, _18698_, _17478_);
  and _44303_ (_18720_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _44304_ (_18731_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _44305_ (_18742_, _18731_, _18720_);
  and _44306_ (_18753_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _44307_ (_18763_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _44308_ (_18774_, _18763_, _18753_);
  and _44309_ (_18785_, _18774_, _18742_);
  and _44310_ (_18796_, _16681_, _15868_);
  and _44311_ (_18807_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _44312_ (_18818_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor _44313_ (_18829_, _18818_, _18807_);
  not _44314_ (_18840_, _18829_);
  nor _44315_ (_18851_, _18840_, _18796_);
  and _44316_ (_18861_, _18851_, _18785_);
  not _44317_ (_18872_, _18861_);
  and _44318_ (_18883_, _18872_, _16493_);
  and _44319_ (_18894_, _18883_, _18709_);
  and _44320_ (_18905_, _18698_, _16493_);
  not _44321_ (_18916_, _18905_);
  and _44322_ (_18927_, _18872_, _17478_);
  and _44323_ (_18938_, _18927_, _18916_);
  and _44324_ (_18948_, _18938_, _18361_);
  nor _44325_ (_18959_, _18948_, _18894_);
  and _44326_ (_18970_, _18350_, _17478_);
  nor _44327_ (_18981_, _18970_, _18023_);
  nor _44328_ (_18992_, _18981_, _18372_);
  not _44329_ (_19003_, _18992_);
  nor _44330_ (_19014_, _19003_, _18959_);
  nor _44331_ (_19025_, _18404_, _18372_);
  nor _44332_ (_19035_, _19025_, _18415_);
  and _44333_ (_19046_, _19035_, _19014_);
  nor _44334_ (_19057_, _18437_, _18415_);
  nor _44335_ (_19068_, _19057_, _18448_);
  and _44336_ (_19079_, _19068_, _19046_);
  and _44337_ (_19090_, _16526_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _44338_ (_19101_, _16570_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _44339_ (_19112_, _19101_, _19090_);
  and _44340_ (_19122_, _16637_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _44341_ (_19133_, _16604_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _44342_ (_19144_, _19133_, _19122_);
  and _44343_ (_19155_, _19144_, _19112_);
  and _44344_ (_19166_, _16681_, _16230_);
  and _44345_ (_19177_, _16736_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _44346_ (_19188_, _16714_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44347_ (_19199_, _19188_, _19177_);
  not _44348_ (_19210_, _19199_);
  nor _44349_ (_19221_, _19210_, _19166_);
  and _44350_ (_19231_, _19221_, _19155_);
  not _44351_ (_19242_, _19231_);
  and _44352_ (_19253_, _19242_, _17478_);
  and _44353_ (_19264_, _19253_, _18905_);
  nor _44354_ (_19275_, _18883_, _18709_);
  nor _44355_ (_19286_, _19275_, _18894_);
  and _44356_ (_19297_, _19286_, _19264_);
  nor _44357_ (_19308_, _18938_, _18361_);
  nor _44358_ (_19319_, _19308_, _18948_);
  and _44359_ (_19330_, _19319_, _19297_);
  and _44360_ (_19340_, _19003_, _18959_);
  nor _44361_ (_19351_, _19340_, _19014_);
  and _44362_ (_19362_, _19351_, _19330_);
  nor _44363_ (_19373_, _19035_, _19014_);
  nor _44364_ (_19384_, _19373_, _19046_);
  and _44365_ (_19395_, _19384_, _19362_);
  nor _44366_ (_19406_, _19068_, _19046_);
  nor _44367_ (_19417_, _19406_, _19079_);
  and _44368_ (_19428_, _19417_, _19395_);
  nor _44369_ (_19439_, _19428_, _19079_);
  nor _44370_ (_19450_, _19439_, _18535_);
  nor _44371_ (_19460_, _19450_, _18502_);
  and _44372_ (_19471_, _18164_, _17674_);
  nor _44373_ (_19482_, _19471_, _18175_);
  not _44374_ (_19493_, _19482_);
  nor _44375_ (_19504_, _19493_, _19460_);
  or _44376_ (_19515_, _19504_, _18088_);
  nor _44377_ (_19526_, _19515_, _18175_);
  nor _44378_ (_19537_, _19526_, _15736_);
  and _44379_ (_19548_, _19526_, _15736_);
  nor _44380_ (_19559_, _19548_, _19537_);
  not _44381_ (_19569_, _19559_);
  and _44382_ (_19580_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _44383_ (_19591_, _19493_, _19460_);
  nor _44384_ (_19602_, _19591_, _19504_);
  and _44385_ (_19613_, _19602_, _19580_);
  and _44386_ (_19624_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and _44387_ (_19635_, _19439_, _18535_);
  nor _44388_ (_19646_, _19635_, _19450_);
  and _44389_ (_19657_, _19646_, _19624_);
  nor _44390_ (_19668_, _19646_, _19624_);
  nor _44391_ (_19679_, _19668_, _19657_);
  not _44392_ (_19689_, _19679_);
  and _44393_ (_19700_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor _44394_ (_19711_, _19417_, _19395_);
  nor _44395_ (_19722_, _19711_, _19428_);
  and _44396_ (_19733_, _19722_, _19700_);
  nor _44397_ (_19744_, _19722_, _19700_);
  nor _44398_ (_19755_, _19744_, _19733_);
  not _44399_ (_19766_, _19755_);
  and _44400_ (_19777_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor _44401_ (_19788_, _19384_, _19362_);
  nor _44402_ (_19799_, _19788_, _19395_);
  and _44403_ (_19809_, _19799_, _19777_);
  nor _44404_ (_19820_, _19799_, _19777_);
  nor _44405_ (_19831_, _19820_, _19809_);
  not _44406_ (_19842_, _19831_);
  and _44407_ (_19853_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor _44408_ (_19864_, _19351_, _19330_);
  nor _44409_ (_19875_, _19864_, _19362_);
  and _44410_ (_19886_, _19875_, _19853_);
  and _44411_ (_19897_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor _44412_ (_19908_, _19319_, _19297_);
  nor _44413_ (_19918_, _19908_, _19330_);
  and _44414_ (_19929_, _19918_, _19897_);
  and _44415_ (_19940_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _44416_ (_19951_, _19286_, _19264_);
  nor _44417_ (_19962_, _19951_, _19297_);
  and _44418_ (_19973_, _19962_, _19940_);
  nor _44419_ (_19984_, _19918_, _19897_);
  nor _44420_ (_19995_, _19984_, _19929_);
  and _44421_ (_20005_, _19995_, _19973_);
  nor _44422_ (_20016_, _20005_, _19929_);
  not _44423_ (_20027_, _20016_);
  nor _44424_ (_20038_, _19875_, _19853_);
  nor _44425_ (_20049_, _20038_, _19886_);
  and _44426_ (_20060_, _20049_, _20027_);
  nor _44427_ (_20071_, _20060_, _19886_);
  nor _44428_ (_20082_, _20071_, _19842_);
  nor _44429_ (_20092_, _20082_, _19809_);
  nor _44430_ (_20103_, _20092_, _19766_);
  nor _44431_ (_20114_, _20103_, _19733_);
  nor _44432_ (_20125_, _20114_, _19689_);
  nor _44433_ (_20136_, _20125_, _19657_);
  nor _44434_ (_20147_, _19602_, _19580_);
  nor _44435_ (_20158_, _20147_, _19613_);
  not _44436_ (_20169_, _20158_);
  nor _44437_ (_20179_, _20169_, _20136_);
  nor _44438_ (_20190_, _20179_, _19613_);
  nor _44439_ (_20201_, _20190_, _19569_);
  nor _44440_ (_20212_, _20201_, _19537_);
  not _44441_ (_20223_, _20212_);
  and _44442_ (_20234_, _20223_, _15715_);
  and _44443_ (_20245_, _20234_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _44444_ (_20256_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _44445_ (_20266_, _20256_, _20245_);
  and _44446_ (_20277_, _20266_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _44447_ (_20288_, _20277_, _15704_);
  and _44448_ (_20299_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _44449_ (_20310_, _20299_, _20288_);
  and _44450_ (_20321_, _20288_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _44451_ (_20332_, _20321_, _20310_);
  and _44452_ (_24614_, _20332_, _41755_);
  nor _44453_ (_20352_, _15573_, _15606_);
  and _44454_ (_20363_, _15573_, _15606_);
  or _44455_ (_20374_, _20363_, _20352_);
  and _44456_ (_02465_, _20374_, _41755_);
  and _44457_ (_20395_, _19242_, _16493_);
  and _44458_ (_02660_, _20395_, _41755_);
  nor _44459_ (_20416_, _19253_, _18905_);
  nor _44460_ (_20427_, _20416_, _19264_);
  and _44461_ (_02854_, _20427_, _41755_);
  nor _44462_ (_20447_, _19962_, _19940_);
  nor _44463_ (_20458_, _20447_, _19973_);
  and _44464_ (_03058_, _20458_, _41755_);
  nor _44465_ (_20479_, _19995_, _19973_);
  nor _44466_ (_20490_, _20479_, _20005_);
  and _44467_ (_03269_, _20490_, _41755_);
  nor _44468_ (_20511_, _20049_, _20027_);
  nor _44469_ (_20522_, _20511_, _20060_);
  and _44470_ (_03470_, _20522_, _41755_);
  and _44471_ (_20542_, _20071_, _19842_);
  nor _44472_ (_20553_, _20542_, _20082_);
  and _44473_ (_03671_, _20553_, _41755_);
  and _44474_ (_20574_, _20092_, _19766_);
  nor _44475_ (_20585_, _20574_, _20103_);
  and _44476_ (_03872_, _20585_, _41755_);
  and _44477_ (_20605_, _20114_, _19689_);
  nor _44478_ (_20616_, _20605_, _20125_);
  and _44479_ (_04073_, _20616_, _41755_);
  and _44480_ (_20637_, _20169_, _20136_);
  nor _44481_ (_20648_, _20637_, _20179_);
  and _44482_ (_04174_, _20648_, _41755_);
  and _44483_ (_20669_, _20190_, _19569_);
  nor _44484_ (_20680_, _20669_, _20201_);
  and _44485_ (_04275_, _20680_, _41755_);
  nor _44486_ (_20700_, _20223_, _15715_);
  nor _44487_ (_20711_, _20700_, _20234_);
  and _44488_ (_04376_, _20711_, _41755_);
  and _44489_ (_20732_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _44490_ (_20743_, _20732_, _20234_);
  nor _44491_ (_20754_, _20743_, _20245_);
  and _44492_ (_04477_, _20754_, _41755_);
  nor _44493_ (_20774_, _20256_, _20245_);
  nor _44494_ (_20785_, _20774_, _20266_);
  and _44495_ (_04578_, _20785_, _41755_);
  and _44496_ (_20806_, _15693_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _44497_ (_20817_, _20806_, _20266_);
  nor _44498_ (_20828_, _20817_, _20277_);
  and _44499_ (_04679_, _20828_, _41755_);
  nor _44500_ (_20849_, _20277_, _15704_);
  nor _44501_ (_20859_, _20849_, _20288_);
  and _44502_ (_04780_, _20859_, _41755_);
  and _44503_ (_20880_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15507_);
  nor _44504_ (_20891_, _20880_, _15518_);
  not _44505_ (_20902_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _44506_ (_20913_, _15540_, _20902_);
  and _44507_ (_20924_, _20913_, _20891_);
  and _44508_ (_20935_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _44509_ (_20946_, _20935_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44510_ (_20956_, _20935_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44511_ (_20967_, _20956_, _20946_);
  and _44512_ (_00863_, _20967_, _41755_);
  and _44513_ (_00894_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _41755_);
  not _44514_ (_20998_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _44515_ (_21009_, _17292_, _20998_);
  and _44516_ (_21020_, _16966_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44517_ (_21031_, _21020_, _21009_);
  nor _44518_ (_21041_, _21031_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44519_ (_21052_, _17119_, _20998_);
  and _44520_ (_21063_, _17456_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _44521_ (_21074_, _21063_, _21052_);
  and _44522_ (_21085_, _21074_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44523_ (_21096_, _21085_, _21041_);
  nor _44524_ (_21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44525_ (_21118_, _21107_, _17630_);
  nor _44526_ (_21128_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor _44527_ (_21139_, _21128_, _21118_);
  not _44528_ (_21150_, _21139_);
  and _44529_ (_21161_, _16296_, _20998_);
  and _44530_ (_21172_, _15967_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44531_ (_21183_, _21172_, _21161_);
  nor _44532_ (_21194_, _21183_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44533_ (_21204_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44534_ (_21215_, _16131_, _20998_);
  and _44535_ (_21226_, _16471_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44536_ (_21237_, _21226_, _21215_);
  nor _44537_ (_21248_, _21237_, _21204_);
  nor _44538_ (_21259_, _21248_, _21194_);
  nor _44539_ (_21270_, _21259_, _21150_);
  and _44540_ (_21281_, _21259_, _21150_);
  nor _44541_ (_21292_, _21281_, _21270_);
  and _44542_ (_21302_, _21107_, _16790_);
  nor _44543_ (_21313_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor _44544_ (_21324_, _21313_, _21302_);
  not _44545_ (_21335_, _21324_);
  nor _44546_ (_21346_, _17292_, _20998_);
  nor _44547_ (_21357_, _21346_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44548_ (_21368_, _16966_, _20998_);
  and _44549_ (_21379_, _17119_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44550_ (_21389_, _21379_, _21368_);
  nor _44551_ (_21400_, _21389_, _21204_);
  nor _44552_ (_21411_, _21400_, _21357_);
  nor _44553_ (_21422_, _21411_, _21335_);
  and _44554_ (_21433_, _21411_, _21335_);
  nor _44555_ (_21444_, _21433_, _21422_);
  not _44556_ (_21455_, _21444_);
  nor _44557_ (_21466_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and _44558_ (_21476_, _21107_, _17826_);
  nor _44559_ (_21498_, _21476_, _21466_);
  not _44560_ (_21510_, _21498_);
  nor _44561_ (_21522_, _16296_, _20998_);
  nor _44562_ (_21534_, _21522_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44563_ (_21546_, _15967_, _20998_);
  and _44564_ (_21558_, _16131_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44565_ (_21559_, _21558_, _21546_);
  nor _44566_ (_21569_, _21559_, _21204_);
  nor _44567_ (_21580_, _21569_, _21534_);
  nor _44568_ (_21591_, _21580_, _21510_);
  and _44569_ (_21602_, _21580_, _21510_);
  nor _44570_ (_21613_, _21602_, _21591_);
  not _44571_ (_21624_, _21613_);
  and _44572_ (_21635_, _21031_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44573_ (_21646_, _21635_);
  nor _44574_ (_21656_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and _44575_ (_21667_, _21107_, _18001_);
  nor _44576_ (_21678_, _21667_, _21656_);
  and _44577_ (_21689_, _21678_, _21646_);
  and _44578_ (_21700_, _21183_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44579_ (_21711_, _21700_);
  and _44580_ (_21722_, _21107_, _18339_);
  nor _44581_ (_21733_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor _44582_ (_21743_, _21733_, _21722_);
  and _44583_ (_21754_, _21743_, _21711_);
  nor _44584_ (_21765_, _21743_, _21711_);
  nor _44585_ (_21776_, _21765_, _21754_);
  not _44586_ (_21787_, _21776_);
  and _44587_ (_21798_, _21346_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44588_ (_21809_, _21798_);
  and _44589_ (_21820_, _21107_, _18861_);
  nor _44590_ (_21830_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _44591_ (_21841_, _21830_, _21820_);
  and _44592_ (_21852_, _21841_, _21809_);
  and _44593_ (_21863_, _21522_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44594_ (_21874_, _21863_);
  nor _44595_ (_21885_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and _44596_ (_21896_, _21107_, _18687_);
  nor _44597_ (_21907_, _21896_, _21885_);
  nor _44598_ (_21917_, _21907_, _21874_);
  not _44599_ (_21928_, _21917_);
  nor _44600_ (_21939_, _21841_, _21809_);
  nor _44601_ (_21950_, _21939_, _21852_);
  and _44602_ (_21961_, _21950_, _21928_);
  nor _44603_ (_21972_, _21961_, _21852_);
  nor _44604_ (_21983_, _21972_, _21787_);
  nor _44605_ (_21994_, _21983_, _21754_);
  nor _44606_ (_22004_, _21678_, _21646_);
  nor _44607_ (_22015_, _22004_, _21689_);
  not _44608_ (_22026_, _22015_);
  nor _44609_ (_22037_, _22026_, _21994_);
  nor _44610_ (_22048_, _22037_, _21689_);
  nor _44611_ (_22069_, _22048_, _21624_);
  nor _44612_ (_22070_, _22069_, _21591_);
  nor _44613_ (_22081_, _22070_, _21455_);
  nor _44614_ (_22091_, _22081_, _21422_);
  not _44615_ (_22102_, _22091_);
  and _44616_ (_22113_, _22102_, _21292_);
  or _44617_ (_22124_, _22113_, _21270_);
  and _44618_ (_22135_, _17456_, _16471_);
  or _44619_ (_22146_, _22135_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _44620_ (_22157_, _21237_);
  and _44621_ (_22168_, _21074_, _22157_);
  nor _44622_ (_22178_, _21559_, _21389_);
  and _44623_ (_22189_, _22178_, _22168_);
  or _44624_ (_22200_, _22189_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44625_ (_22211_, _22200_, _22146_);
  and _44626_ (_22222_, _22211_, _22124_);
  and _44627_ (_22233_, _22222_, _21096_);
  nor _44628_ (_22244_, _22102_, _21292_);
  or _44629_ (_22255_, _22244_, _22113_);
  and _44630_ (_22266_, _22255_, _22233_);
  nor _44631_ (_22276_, _22233_, _21139_);
  nor _44632_ (_22287_, _22276_, _22266_);
  not _44633_ (_22298_, _22287_);
  and _44634_ (_22309_, _22287_, _21096_);
  not _44635_ (_22331_, _21259_);
  and _44636_ (_22332_, _22070_, _21455_);
  or _44637_ (_22343_, _22332_, _22081_);
  and _44638_ (_22354_, _22343_, _22233_);
  nor _44639_ (_22364_, _22233_, _21324_);
  nor _44640_ (_22375_, _22364_, _22354_);
  and _44641_ (_22386_, _22375_, _22331_);
  nor _44642_ (_22397_, _22375_, _22331_);
  nor _44643_ (_22408_, _22397_, _22386_);
  not _44644_ (_22419_, _22408_);
  not _44645_ (_22430_, _21411_);
  nor _44646_ (_22441_, _22233_, _21510_);
  and _44647_ (_22452_, _22048_, _21624_);
  nor _44648_ (_22463_, _22452_, _22069_);
  and _44649_ (_22474_, _22463_, _22233_);
  or _44650_ (_22485_, _22474_, _22441_);
  and _44651_ (_22496_, _22485_, _22430_);
  nor _44652_ (_22507_, _22485_, _22430_);
  not _44653_ (_22518_, _21580_);
  and _44654_ (_22529_, _22026_, _21994_);
  or _44655_ (_22539_, _22529_, _22037_);
  and _44656_ (_22550_, _22539_, _22233_);
  nor _44657_ (_22561_, _22233_, _21678_);
  nor _44658_ (_22572_, _22561_, _22550_);
  and _44659_ (_22583_, _22572_, _22518_);
  and _44660_ (_22594_, _21972_, _21787_);
  nor _44661_ (_22605_, _22594_, _21983_);
  not _44662_ (_22616_, _22605_);
  and _44663_ (_22626_, _22616_, _22233_);
  nor _44664_ (_22637_, _22233_, _21743_);
  nor _44665_ (_22648_, _22637_, _22626_);
  and _44666_ (_22659_, _22648_, _21646_);
  nor _44667_ (_22670_, _22648_, _21646_);
  nor _44668_ (_22681_, _22670_, _22659_);
  not _44669_ (_22692_, _22681_);
  nor _44670_ (_22703_, _21950_, _21928_);
  nor _44671_ (_22713_, _22703_, _21961_);
  not _44672_ (_22724_, _22713_);
  and _44673_ (_22735_, _22724_, _22233_);
  nor _44674_ (_22746_, _22233_, _21841_);
  nor _44675_ (_22757_, _22746_, _22735_);
  and _44676_ (_22768_, _22757_, _21711_);
  and _44677_ (_22779_, _22233_, _21863_);
  nor _44678_ (_22790_, _22779_, _21907_);
  and _44679_ (_22800_, _22779_, _21907_);
  nor _44680_ (_22811_, _22800_, _22790_);
  and _44681_ (_22822_, _22811_, _21809_);
  nor _44682_ (_22833_, _22811_, _21809_);
  nor _44683_ (_22844_, _22833_, _22822_);
  nor _44684_ (_22855_, _21107_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and _44685_ (_22866_, _21107_, _19231_);
  nor _44686_ (_22877_, _22866_, _22855_);
  nor _44687_ (_22887_, _22877_, _21874_);
  not _44688_ (_22898_, _22887_);
  and _44689_ (_22909_, _22898_, _22844_);
  nor _44690_ (_22920_, _22909_, _22822_);
  nor _44691_ (_22931_, _22757_, _21711_);
  nor _44692_ (_22942_, _22931_, _22768_);
  not _44693_ (_22953_, _22942_);
  nor _44694_ (_22964_, _22953_, _22920_);
  nor _44695_ (_22974_, _22964_, _22768_);
  nor _44696_ (_22985_, _22974_, _22692_);
  nor _44697_ (_23006_, _22985_, _22659_);
  nor _44698_ (_23007_, _22572_, _22518_);
  nor _44699_ (_23018_, _23007_, _22583_);
  not _44700_ (_23039_, _23018_);
  nor _44701_ (_23040_, _23039_, _23006_);
  nor _44702_ (_23051_, _23040_, _22583_);
  nor _44703_ (_23072_, _23051_, _22507_);
  nor _44704_ (_23073_, _23072_, _22496_);
  nor _44705_ (_23083_, _23073_, _22419_);
  or _44706_ (_23104_, _23083_, _22386_);
  or _44707_ (_23105_, _23104_, _22309_);
  and _44708_ (_23116_, _23105_, _22211_);
  nor _44709_ (_23137_, _23116_, _22298_);
  and _44710_ (_23138_, _22309_, _22211_);
  and _44711_ (_23149_, _23138_, _23104_);
  or _44712_ (_23170_, _23149_, _23137_);
  and _44713_ (_00915_, _23170_, _41755_);
  or _44714_ (_23181_, _22287_, _21096_);
  and _44715_ (_23201_, _23181_, _23116_);
  and _44716_ (_03015_, _23201_, _41755_);
  and _44717_ (_03026_, _22233_, _41755_);
  and _44718_ (_03047_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _41755_);
  and _44719_ (_03069_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _41755_);
  and _44720_ (_03090_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _41755_);
  or _44721_ (_23252_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44722_ (_23263_, _20935_, rst);
  and _44723_ (_03101_, _23263_, _23252_);
  and _44724_ (_23284_, _23201_, _21863_);
  or _44725_ (_23295_, _23284_, _22877_);
  nand _44726_ (_23305_, _23284_, _22877_);
  and _44727_ (_23316_, _23305_, _23295_);
  and _44728_ (_03112_, _23316_, _41755_);
  nor _44729_ (_23337_, _22898_, _22844_);
  or _44730_ (_23348_, _23337_, _22909_);
  nand _44731_ (_23359_, _23348_, _23201_);
  or _44732_ (_23370_, _23201_, _22811_);
  and _44733_ (_23381_, _23370_, _23359_);
  and _44734_ (_03123_, _23381_, _41755_);
  and _44735_ (_23402_, _22953_, _22920_);
  or _44736_ (_23413_, _23402_, _22964_);
  nand _44737_ (_23423_, _23413_, _23201_);
  or _44738_ (_23434_, _23201_, _22757_);
  and _44739_ (_23445_, _23434_, _23423_);
  and _44740_ (_03134_, _23445_, _41755_);
  and _44741_ (_23466_, _22974_, _22692_);
  or _44742_ (_23477_, _23466_, _22985_);
  nand _44743_ (_23488_, _23477_, _23201_);
  or _44744_ (_23499_, _23201_, _22648_);
  and _44745_ (_23510_, _23499_, _23488_);
  and _44746_ (_03145_, _23510_, _41755_);
  and _44747_ (_23531_, _23039_, _23006_);
  or _44748_ (_23541_, _23531_, _23040_);
  nand _44749_ (_23552_, _23541_, _23201_);
  or _44750_ (_23563_, _23201_, _22572_);
  and _44751_ (_23574_, _23563_, _23552_);
  and _44752_ (_03156_, _23574_, _41755_);
  or _44753_ (_23595_, _22507_, _22496_);
  and _44754_ (_23606_, _23595_, _23051_);
  nor _44755_ (_23617_, _23595_, _23051_);
  or _44756_ (_23628_, _23617_, _23606_);
  nand _44757_ (_23639_, _23628_, _23201_);
  or _44758_ (_23649_, _23201_, _22485_);
  and _44759_ (_23660_, _23649_, _23639_);
  and _44760_ (_03167_, _23660_, _41755_);
  and _44761_ (_23681_, _23073_, _22419_);
  or _44762_ (_23692_, _23681_, _23083_);
  nand _44763_ (_23703_, _23692_, _23201_);
  or _44764_ (_23714_, _23201_, _22375_);
  and _44765_ (_23725_, _23714_, _23703_);
  and _44766_ (_03178_, _23725_, _41755_);
  not _44767_ (_23746_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _44768_ (_23757_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15507_);
  and _44769_ (_23767_, _23757_, _23746_);
  and _44770_ (_23778_, _23767_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44771_ (_23789_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  not _44772_ (_23800_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44773_ (_23811_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15507_);
  and _44774_ (_23822_, _23811_, _23800_);
  and _44775_ (_23833_, _23822_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _44776_ (_23844_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44777_ (_23855_, _23844_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44778_ (_23866_, _23844_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44779_ (_23876_, _23866_, _23855_);
  and _44780_ (_23887_, _23876_, _23833_);
  nor _44781_ (_23898_, _23887_, _23789_);
  nor _44782_ (_23909_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44783_ (_23920_, _23909_, _23811_);
  and _44784_ (_23931_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _44785_ (_23942_, _23909_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _44786_ (_23953_, _23942_, _23811_);
  and _44787_ (_23964_, _23953_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  and _44788_ (_23975_, _23767_, _23800_);
  and _44789_ (_23985_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or _44790_ (_23996_, _23985_, _23964_);
  nor _44791_ (_24007_, _23996_, _23931_);
  and _44792_ (_24018_, _24007_, _23898_);
  and _44793_ (_24029_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor _44794_ (_24040_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _44795_ (_24051_, _24040_, _23844_);
  and _44796_ (_24062_, _24051_, _23833_);
  nor _44797_ (_24073_, _24062_, _24029_);
  and _44798_ (_24084_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _44799_ (_24095_, _23953_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _44800_ (_24105_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _44801_ (_24116_, _24105_, _24095_);
  nor _44802_ (_24127_, _24116_, _24084_);
  and _44803_ (_24138_, _24127_, _24073_);
  and _44804_ (_24149_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and _44805_ (_24160_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _44806_ (_24182_, _24160_, _24149_);
  and _44807_ (_24194_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not _44808_ (_24206_, _24194_);
  not _44809_ (_24218_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44810_ (_24229_, _23833_, _24218_);
  and _44811_ (_24241_, _23953_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _44812_ (_24253_, _24241_, _24229_);
  and _44813_ (_24254_, _24253_, _24206_);
  and _44814_ (_24265_, _24254_, _24182_);
  and _44815_ (_24276_, _24265_, _24138_);
  and _44816_ (_24287_, _24276_, _24018_);
  and _44817_ (_24298_, _23855_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _44818_ (_24309_, _24298_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _44819_ (_24320_, _24309_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _44820_ (_24331_, _24320_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _44821_ (_24341_, _24331_);
  not _44822_ (_24352_, _23833_);
  nor _44823_ (_24363_, _24320_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _44824_ (_24374_, _24363_, _24352_);
  and _44825_ (_24385_, _24374_, _24341_);
  not _44826_ (_24396_, _24385_);
  and _44827_ (_24407_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44828_ (_24418_, _24407_, _23811_);
  and _44829_ (_24429_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _44830_ (_24440_, _24429_, _24418_);
  and _44831_ (_24451_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _44832_ (_24461_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _44833_ (_24472_, _24461_, _24451_);
  and _44834_ (_24483_, _24472_, _24440_);
  and _44835_ (_24494_, _24483_, _24396_);
  nor _44836_ (_24505_, _24309_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _44837_ (_24516_, _24505_);
  nor _44838_ (_24527_, _24320_, _24352_);
  and _44839_ (_24538_, _24527_, _24516_);
  not _44840_ (_24549_, _24538_);
  and _44841_ (_24560_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _44842_ (_24571_, _24560_, _24418_);
  and _44843_ (_24581_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _44844_ (_24592_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _44845_ (_24603_, _24592_, _24581_);
  and _44846_ (_24615_, _24603_, _24571_);
  and _44847_ (_24626_, _24615_, _24549_);
  nor _44848_ (_24637_, _24626_, _24494_);
  not _44849_ (_24648_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _44850_ (_24659_, _24331_, _24648_);
  and _44851_ (_24669_, _24331_, _24648_);
  nor _44852_ (_24680_, _24669_, _24659_);
  nor _44853_ (_24691_, _24680_, _24352_);
  not _44854_ (_24702_, _24691_);
  and _44855_ (_24713_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor _44856_ (_24724_, _24713_, _24418_);
  and _44857_ (_24735_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _44858_ (_24746_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _44859_ (_24756_, _24746_, _24735_);
  and _44860_ (_24767_, _24756_, _24724_);
  and _44861_ (_24778_, _24767_, _24702_);
  not _44862_ (_24789_, _24778_);
  not _44863_ (_24800_, _24298_);
  nor _44864_ (_24811_, _23855_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _44865_ (_24822_, _24811_, _24352_);
  and _44866_ (_24833_, _24822_, _24800_);
  not _44867_ (_24844_, _24833_);
  and _44868_ (_24854_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and _44869_ (_24865_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _44870_ (_24876_, _24865_, _24854_);
  and _44871_ (_24887_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _44872_ (_24898_, _23953_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor _44873_ (_24909_, _24898_, _24887_);
  and _44874_ (_24920_, _24909_, _24876_);
  and _44875_ (_24931_, _24920_, _24844_);
  not _44876_ (_24942_, _24931_);
  and _44877_ (_24952_, _23920_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _44878_ (_24963_, _24952_, _24418_);
  and _44879_ (_24974_, _23778_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not _44880_ (_24985_, _24974_);
  and _44881_ (_24996_, _24985_, _24963_);
  nor _44882_ (_25007_, _24298_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _44883_ (_25018_, _25007_);
  nor _44884_ (_25029_, _24309_, _24352_);
  and _44885_ (_25039_, _25029_, _25018_);
  and _44886_ (_25050_, _23975_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and _44887_ (_25061_, _23953_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _44888_ (_25072_, _25061_, _25050_);
  not _44889_ (_25083_, _25072_);
  nor _44890_ (_25104_, _25083_, _25039_);
  and _44891_ (_25105_, _25104_, _24996_);
  nor _44892_ (_25116_, _25105_, _24942_);
  and _44893_ (_25127_, _25116_, _24789_);
  and _44894_ (_25147_, _25127_, _24637_);
  nand _44895_ (_25148_, _25147_, _24287_);
  and _44896_ (_25159_, _23170_, _20924_);
  not _44897_ (_25180_, _25159_);
  and _44898_ (_25181_, _20332_, _15573_);
  nor _44899_ (_25192_, _16790_, _16471_);
  and _44900_ (_25203_, _16790_, _16471_);
  nor _44901_ (_25214_, _25203_, _25192_);
  not _44902_ (_25234_, _25214_);
  nor _44903_ (_25235_, _17826_, _17119_);
  and _44904_ (_25246_, _17826_, _17119_);
  nor _44905_ (_25257_, _25246_, _25235_);
  nor _44906_ (_25268_, _18001_, _16131_);
  and _44907_ (_25279_, _25268_, _25257_);
  nor _44908_ (_25290_, _25279_, _25235_);
  nor _44909_ (_25301_, _25290_, _25234_);
  and _44910_ (_25312_, _18001_, _16131_);
  nor _44911_ (_25322_, _25312_, _25268_);
  nor _44912_ (_25333_, _18339_, _16966_);
  and _44913_ (_25344_, _18339_, _16966_);
  nor _44914_ (_25365_, _25344_, _25333_);
  nor _44915_ (_25366_, _18861_, _15967_);
  and _44916_ (_25377_, _18861_, _15967_);
  nor _44917_ (_25388_, _25377_, _25366_);
  not _44918_ (_25399_, _25388_);
  nor _44919_ (_25410_, _18687_, _17292_);
  nor _44920_ (_25420_, _19231_, _16296_);
  and _44921_ (_25431_, _18687_, _17292_);
  nor _44922_ (_25442_, _25431_, _25410_);
  and _44923_ (_25453_, _25442_, _25420_);
  nor _44924_ (_25464_, _25453_, _25410_);
  nor _44925_ (_25475_, _25464_, _25399_);
  nor _44926_ (_25486_, _25475_, _25366_);
  nor _44927_ (_25497_, _25486_, _25365_);
  and _44928_ (_25507_, _25486_, _25365_);
  nor _44929_ (_25518_, _25507_, _25497_);
  not _44930_ (_25539_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _44931_ (_25540_, _15780_, _25539_);
  not _44932_ (_25551_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _44933_ (_25562_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44934_ (_25573_, _25562_, _17347_);
  nor _44935_ (_25584_, _25573_, _25551_);
  nor _44936_ (_25595_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44937_ (_25605_, _25595_, _16022_);
  not _44938_ (_25616_, _25605_);
  not _44939_ (_25627_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _44940_ (_25638_, _25627_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44941_ (_25649_, _25638_, _16362_);
  not _44942_ (_25660_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44943_ (_25671_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25660_);
  and _44944_ (_25682_, _25671_, _17010_);
  nor _44945_ (_25693_, _25682_, _25649_);
  and _44946_ (_25703_, _25693_, _25616_);
  and _44947_ (_25714_, _25703_, _25584_);
  and _44948_ (_25735_, _25562_, _16856_);
  nor _44949_ (_25736_, _25735_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _44950_ (_25747_, _25671_, _17173_);
  not _44951_ (_25758_, _25747_);
  and _44952_ (_25769_, _25638_, _15824_);
  and _44953_ (_25780_, _25595_, _16186_);
  nor _44954_ (_25790_, _25780_, _25769_);
  and _44955_ (_25801_, _25790_, _25758_);
  and _44956_ (_25812_, _25801_, _25736_);
  nor _44957_ (_25823_, _25812_, _25714_);
  nor _44958_ (_25834_, _25823_, _15780_);
  nor _44959_ (_25845_, _25834_, _25540_);
  and _44960_ (_25856_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _44961_ (_25867_, _25856_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _44962_ (_25878_, _25867_);
  and _44963_ (_25888_, _25878_, _25845_);
  and _44964_ (_25899_, _25878_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _44965_ (_25910_, _25899_, _25888_);
  and _44966_ (_25921_, _19231_, _16296_);
  nor _44967_ (_25932_, _25921_, _25420_);
  not _44968_ (_25943_, _25932_);
  nor _44969_ (_25954_, _25943_, _25910_);
  and _44970_ (_25965_, _25954_, _25442_);
  and _44971_ (_25976_, _25464_, _25399_);
  nor _44972_ (_25987_, _25976_, _25475_);
  and _44973_ (_25998_, _25987_, _25965_);
  not _44974_ (_26009_, _25998_);
  nor _44975_ (_26020_, _26009_, _25518_);
  nor _44976_ (_26031_, _25486_, _25344_);
  or _44977_ (_26042_, _26031_, _25333_);
  or _44978_ (_26053_, _26042_, _26020_);
  and _44979_ (_26064_, _26053_, _25322_);
  and _44980_ (_26085_, _26064_, _25257_);
  and _44981_ (_26086_, _25290_, _25234_);
  nor _44982_ (_26097_, _26086_, _25301_);
  and _44983_ (_26108_, _26097_, _26085_);
  or _44984_ (_26119_, _26108_, _25301_);
  nor _44985_ (_26130_, _26119_, _25192_);
  nor _44986_ (_26141_, _17630_, _17456_);
  and _44987_ (_26152_, _17630_, _17456_);
  nor _44988_ (_26162_, _26152_, _26141_);
  not _44989_ (_26173_, _26162_);
  and _44990_ (_26194_, _26173_, _26130_);
  nor _44991_ (_26195_, _26173_, _26130_);
  not _44992_ (_26206_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _44993_ (_26217_, _20880_, _26206_);
  and _44994_ (_26228_, _26217_, _15562_);
  not _44995_ (_26239_, _26228_);
  or _44996_ (_26250_, _26239_, _26195_);
  nor _44997_ (_26261_, _26250_, _26194_);
  not _44998_ (_26272_, _26261_);
  not _44999_ (_26283_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _45000_ (_26294_, _15518_, _26283_);
  and _45001_ (_26305_, _26294_, _15562_);
  not _45002_ (_26316_, _26305_);
  not _45003_ (_26327_, _16471_);
  nor _45004_ (_26338_, _16790_, _26327_);
  not _45005_ (_26349_, _17119_);
  nor _45006_ (_26360_, _17826_, _26349_);
  not _45007_ (_26371_, _16131_);
  and _45008_ (_26382_, _18001_, _26371_);
  nor _45009_ (_26393_, _26382_, _25257_);
  nor _45010_ (_26404_, _26393_, _26360_);
  nor _45011_ (_26415_, _26404_, _25214_);
  nor _45012_ (_26426_, _26415_, _26338_);
  and _45013_ (_26437_, _26404_, _25214_);
  nor _45014_ (_26448_, _26437_, _26415_);
  not _45015_ (_26459_, _26448_);
  and _45016_ (_26470_, _26382_, _25257_);
  nor _45017_ (_26481_, _26470_, _26393_);
  not _45018_ (_26492_, _26481_);
  not _45019_ (_26503_, _25322_);
  not _45020_ (_26514_, _16296_);
  and _45021_ (_26525_, _19231_, _26514_);
  nor _45022_ (_26536_, _26525_, _25442_);
  not _45023_ (_26546_, _17292_);
  nor _45024_ (_26557_, _18687_, _26546_);
  nor _45025_ (_26568_, _26557_, _26536_);
  nor _45026_ (_26579_, _26568_, _25388_);
  not _45027_ (_26590_, _15967_);
  nor _45028_ (_26601_, _18861_, _26590_);
  nor _45029_ (_26612_, _26601_, _26579_);
  nor _45030_ (_26623_, _26612_, _25365_);
  and _45031_ (_26644_, _26612_, _25365_);
  nor _45032_ (_26645_, _26644_, _26623_);
  not _45033_ (_26656_, _26645_);
  and _45034_ (_26667_, _26568_, _25388_);
  nor _45035_ (_26678_, _26667_, _26579_);
  not _45036_ (_26689_, _26678_);
  and _45037_ (_26700_, _26525_, _25442_);
  nor _45038_ (_26711_, _26700_, _26536_);
  not _45039_ (_26722_, _26711_);
  nor _45040_ (_26733_, _25932_, _25910_);
  and _45041_ (_26744_, _26733_, _26722_);
  and _45042_ (_26755_, _26744_, _26689_);
  and _45043_ (_26766_, _26755_, _26656_);
  not _45044_ (_26777_, _16966_);
  or _45045_ (_26788_, _18339_, _26777_);
  and _45046_ (_26799_, _18339_, _26777_);
  or _45047_ (_26810_, _26612_, _26799_);
  and _45048_ (_26821_, _26810_, _26788_);
  or _45049_ (_26832_, _26821_, _26766_);
  and _45050_ (_26843_, _26832_, _26503_);
  and _45051_ (_26854_, _26843_, _26492_);
  and _45052_ (_26865_, _26854_, _26459_);
  nor _45053_ (_26876_, _26865_, _26426_);
  nor _45054_ (_26887_, _26876_, _26162_);
  and _45055_ (_26898_, _26876_, _26162_);
  nor _45056_ (_26908_, _26898_, _26887_);
  nor _45057_ (_26919_, _26908_, _26316_);
  and _45058_ (_26940_, _15551_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45059_ (_26941_, _26940_, _26294_);
  nor _45060_ (_26952_, _19231_, _18687_);
  and _45061_ (_26963_, _26952_, _18872_);
  and _45062_ (_26974_, _26963_, _18350_);
  and _45063_ (_26985_, _26974_, _18012_);
  and _45064_ (_26996_, _26985_, _17837_);
  and _45065_ (_27007_, _26996_, _16801_);
  and _45066_ (_27018_, _27007_, _25910_);
  not _45067_ (_27029_, _25910_);
  and _45068_ (_27050_, _16790_, _17826_);
  and _45069_ (_27051_, _18861_, _18687_);
  and _45070_ (_27062_, _27051_, _19231_);
  and _45071_ (_27073_, _27062_, _18339_);
  and _45072_ (_27084_, _27073_, _18001_);
  and _45073_ (_27095_, _27084_, _27050_);
  and _45074_ (_27106_, _27095_, _27029_);
  nor _45075_ (_27117_, _27106_, _27018_);
  and _45076_ (_27128_, _27117_, _17630_);
  nor _45077_ (_27139_, _27117_, _17630_);
  nor _45078_ (_27150_, _27139_, _27128_);
  and _45079_ (_27161_, _27150_, _26941_);
  not _45080_ (_27172_, _17456_);
  nor _45081_ (_27183_, _25910_, _27172_);
  not _45082_ (_27194_, _27183_);
  and _45083_ (_27205_, _25910_, _17630_);
  and _45084_ (_27216_, _26940_, _15529_);
  not _45085_ (_27227_, _27216_);
  nor _45086_ (_27238_, _27227_, _27205_);
  and _45087_ (_27249_, _27238_, _27194_);
  nor _45088_ (_27269_, _27249_, _27161_);
  and _45089_ (_27270_, _26217_, _20913_);
  nor _45090_ (_27281_, _27051_, _18339_);
  and _45091_ (_27292_, _27281_, _27270_);
  and _45092_ (_27303_, _27292_, _18012_);
  nor _45093_ (_27314_, _27303_, _17837_);
  and _45094_ (_27325_, _27314_, _16790_);
  nor _45095_ (_27336_, _27050_, _17630_);
  nor _45096_ (_27347_, _27336_, _27292_);
  and _45097_ (_27358_, _27347_, _25910_);
  nor _45098_ (_27369_, _27358_, _27325_);
  nor _45099_ (_27380_, _27369_, _17641_);
  and _45100_ (_27391_, _27369_, _17641_);
  nor _45101_ (_27402_, _27391_, _27380_);
  and _45102_ (_27413_, _27402_, _27270_);
  not _45103_ (_27424_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _45104_ (_27435_, _15551_, _27424_);
  and _45105_ (_27446_, _27435_, _26217_);
  not _45106_ (_27457_, _27446_);
  nor _45107_ (_27468_, _27457_, _26152_);
  and _45108_ (_27479_, _27435_, _20891_);
  and _45109_ (_27490_, _27479_, _26162_);
  nor _45110_ (_27501_, _27490_, _27468_);
  and _45111_ (_27512_, _27435_, _15518_);
  not _45112_ (_27533_, _27512_);
  nor _45113_ (_27534_, _27533_, _16790_);
  and _45114_ (_27545_, _26940_, _20891_);
  and _45115_ (_27556_, _27545_, _19242_);
  nor _45116_ (_27567_, _27556_, _27534_);
  and _45117_ (_27578_, _27567_, _27501_);
  and _45118_ (_27589_, _26940_, _26217_);
  not _45119_ (_27600_, _27589_);
  nor _45120_ (_27610_, _27600_, _25910_);
  and _45121_ (_27621_, _20913_, _15529_);
  and _45122_ (_27632_, _27621_, _26141_);
  and _45123_ (_27643_, _26294_, _20913_);
  and _45124_ (_27654_, _27643_, _17630_);
  nor _45125_ (_27665_, _27654_, _27632_);
  and _45126_ (_27676_, _20891_, _15562_);
  not _45127_ (_27687_, _27676_);
  nor _45128_ (_27698_, _27687_, _17630_);
  not _45129_ (_27709_, _27698_);
  nand _45130_ (_27720_, _27709_, _27665_);
  nor _45131_ (_27731_, _27720_, _27610_);
  and _45132_ (_27742_, _27731_, _27578_);
  not _45133_ (_27753_, _27742_);
  nor _45134_ (_27764_, _27753_, _27413_);
  and _45135_ (_27775_, _27764_, _27269_);
  not _45136_ (_27786_, _27775_);
  nor _45137_ (_27797_, _27786_, _26919_);
  and _45138_ (_27818_, _27797_, _26272_);
  not _45139_ (_27819_, _27818_);
  nor _45140_ (_27830_, _27819_, _25181_);
  and _45141_ (_27841_, _27830_, _25180_);
  not _45142_ (_27852_, _27841_);
  or _45143_ (_27863_, _27852_, _25148_);
  and _45144_ (_27874_, \oc8051_top_1.oc8051_decoder1.wr , _15507_);
  not _45145_ (_27885_, _27874_);
  nor _45146_ (_27896_, _27885_, _23822_);
  not _45147_ (_27907_, _27896_);
  nor _45148_ (_27918_, _27907_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not _45149_ (_27929_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _45150_ (_27940_, _25148_, _27929_);
  and _45151_ (_27951_, _27940_, _27918_);
  and _45152_ (_27962_, _27951_, _27863_);
  nor _45153_ (_27972_, _27896_, _27929_);
  nor _45154_ (_27983_, _26195_, _26141_);
  nor _45155_ (_27994_, _27983_, _26239_);
  not _45156_ (_28005_, _27994_);
  and _45157_ (_28016_, _17630_, _27172_);
  nor _45158_ (_28027_, _28016_, _26887_);
  nor _45159_ (_28038_, _28027_, _26316_);
  and _45160_ (_28049_, _25910_, _16790_);
  and _45161_ (_28060_, _28049_, _27314_);
  nor _45162_ (_28071_, _28060_, _27205_);
  not _45163_ (_28082_, _27270_);
  nor _45164_ (_28093_, _25910_, _17630_);
  not _45165_ (_28104_, _28093_);
  nor _45166_ (_28115_, _28104_, _27325_);
  nor _45167_ (_28126_, _28115_, _28082_);
  and _45168_ (_28137_, _28126_, _28071_);
  or _45169_ (_28148_, _28137_, _27292_);
  nor _45170_ (_28159_, _27676_, _25910_);
  nor _45171_ (_28170_, _27643_, _27029_);
  nor _45172_ (_28181_, _28170_, _28159_);
  not _45173_ (_28192_, _28181_);
  nor _45174_ (_28203_, _25899_, _25845_);
  not _45175_ (_28214_, _27479_);
  nor _45176_ (_28225_, _28214_, _25888_);
  nor _45177_ (_28236_, _28225_, _27446_);
  nor _45178_ (_28257_, _28236_, _28203_);
  not _45179_ (_28258_, _28257_);
  nor _45180_ (_28269_, _27600_, _19231_);
  and _45181_ (_28280_, _27435_, _15529_);
  not _45182_ (_28291_, _28280_);
  nor _45183_ (_28302_, _28291_, _17630_);
  nor _45184_ (_28313_, _28302_, _28269_);
  not _45185_ (_28323_, _28313_);
  not _45186_ (_28334_, _25845_);
  and _45187_ (_28345_, _27435_, _26294_);
  nor _45188_ (_28356_, _28345_, _27621_);
  nor _45189_ (_28367_, _28356_, _25867_);
  nor _45190_ (_28378_, _28367_, _28334_);
  and _45191_ (_28389_, _27545_, _25899_);
  nor _45192_ (_28400_, _28389_, _28345_);
  and _45193_ (_28411_, _28400_, _28334_);
  nor _45194_ (_28422_, _28411_, _28378_);
  nor _45195_ (_28443_, _28422_, _28323_);
  and _45196_ (_28444_, _28443_, _28258_);
  and _45197_ (_28455_, _28444_, _28192_);
  not _45198_ (_28466_, _28455_);
  nor _45199_ (_28477_, _28466_, _28148_);
  not _45200_ (_28488_, _28477_);
  nor _45201_ (_28499_, _28488_, _28038_);
  and _45202_ (_28510_, _28499_, _28005_);
  not _45203_ (_28521_, _24018_);
  nor _45204_ (_28532_, _24265_, _24138_);
  and _45205_ (_28543_, _28532_, _28521_);
  and _45206_ (_28554_, _28543_, _25147_);
  nand _45207_ (_28565_, _28554_, _28510_);
  and _45208_ (_28576_, _27896_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or _45209_ (_28587_, _28554_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _45210_ (_28598_, _28587_, _28576_);
  and _45211_ (_28609_, _28598_, _28565_);
  or _45212_ (_28620_, _28609_, _27972_);
  or _45213_ (_28631_, _28620_, _27962_);
  and _45214_ (_06696_, _28631_, _41755_);
  and _45215_ (_28652_, _23316_, _20924_);
  not _45216_ (_28663_, _28652_);
  and _45217_ (_28673_, _20648_, _15573_);
  and _45218_ (_28684_, _25943_, _25910_);
  nor _45219_ (_28695_, _28684_, _25954_);
  not _45220_ (_28706_, _28695_);
  nor _45221_ (_28717_, _26305_, _26228_);
  nor _45222_ (_28728_, _28717_, _28706_);
  nor _45223_ (_28739_, _28291_, _25910_);
  not _45224_ (_28750_, _28739_);
  nor _45225_ (_28761_, _28214_, _25420_);
  nor _45226_ (_28772_, _28761_, _27446_);
  or _45227_ (_28783_, _28772_, _25921_);
  and _45228_ (_28794_, _28345_, _17641_);
  and _45229_ (_28805_, _26940_, _26206_);
  not _45230_ (_28816_, _28805_);
  nor _45231_ (_28827_, _28816_, _18687_);
  nor _45232_ (_28838_, _28827_, _28794_);
  and _45233_ (_28849_, _27621_, _25420_);
  and _45234_ (_28860_, _27643_, _19231_);
  nor _45235_ (_28871_, _28860_, _28849_);
  nor _45236_ (_28882_, _27227_, _16296_);
  and _45237_ (_28893_, _26941_, _19231_);
  nor _45238_ (_28904_, _28893_, _28882_);
  nor _45239_ (_28915_, _27676_, _27270_);
  nor _45240_ (_28926_, _28915_, _19231_);
  not _45241_ (_28937_, _28926_);
  and _45242_ (_28948_, _28937_, _28904_);
  and _45243_ (_28959_, _28948_, _28871_);
  and _45244_ (_28980_, _28959_, _28838_);
  and _45245_ (_28981_, _28980_, _28783_);
  and _45246_ (_28992_, _28981_, _28750_);
  not _45247_ (_29002_, _28992_);
  nor _45248_ (_29013_, _29002_, _28728_);
  not _45249_ (_29024_, _29013_);
  nor _45250_ (_29035_, _29024_, _28673_);
  and _45251_ (_29046_, _29035_, _28663_);
  not _45252_ (_29057_, _29046_);
  or _45253_ (_29068_, _29057_, _25148_);
  not _45254_ (_29079_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _45255_ (_29090_, _25148_, _29079_);
  and _45256_ (_29101_, _29090_, _27918_);
  and _45257_ (_29112_, _29101_, _29068_);
  nor _45258_ (_29123_, _27896_, _29079_);
  not _45259_ (_29134_, _28510_);
  or _45260_ (_29145_, _29134_, _25148_);
  and _45261_ (_29156_, _29090_, _28576_);
  and _45262_ (_29167_, _29156_, _29145_);
  or _45263_ (_29178_, _29167_, _29123_);
  or _45264_ (_29189_, _29178_, _29112_);
  and _45265_ (_08932_, _29189_, _41755_);
  and _45266_ (_29210_, _20680_, _15573_);
  not _45267_ (_29221_, _29210_);
  and _45268_ (_29232_, _23381_, _20924_);
  nor _45269_ (_29243_, _27227_, _17292_);
  and _45270_ (_29254_, _19231_, _18687_);
  nor _45271_ (_29265_, _29254_, _26952_);
  not _45272_ (_29276_, _29265_);
  nor _45273_ (_29287_, _29276_, _25910_);
  and _45274_ (_29298_, _29276_, _25910_);
  nor _45275_ (_29309_, _29298_, _29287_);
  and _45276_ (_29320_, _29309_, _26941_);
  nor _45277_ (_29331_, _29320_, _29243_);
  nor _45278_ (_29341_, _27281_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _45279_ (_29352_, _29341_, _18698_);
  nor _45280_ (_29363_, _29341_, _18698_);
  nor _45281_ (_29374_, _29363_, _29352_);
  nor _45282_ (_29385_, _29374_, _28082_);
  not _45283_ (_29396_, _29385_);
  nor _45284_ (_29407_, _27687_, _18687_);
  nor _45285_ (_29418_, _28816_, _18861_);
  nor _45286_ (_29429_, _27533_, _19231_);
  or _45287_ (_29440_, _29429_, _29418_);
  nor _45288_ (_29451_, _29440_, _29407_);
  and _45289_ (_29462_, _27479_, _25442_);
  and _45290_ (_29473_, _27621_, _25410_);
  nor _45291_ (_29484_, _27457_, _25431_);
  and _45292_ (_29495_, _27643_, _18687_);
  or _45293_ (_29506_, _29495_, _29484_);
  or _45294_ (_29527_, _29506_, _29473_);
  nor _45295_ (_29528_, _29527_, _29462_);
  and _45296_ (_29539_, _29528_, _29451_);
  and _45297_ (_29550_, _29539_, _29396_);
  and _45298_ (_29561_, _29550_, _29331_);
  nor _45299_ (_29572_, _25442_, _25420_);
  or _45300_ (_29583_, _29572_, _25453_);
  and _45301_ (_29594_, _29583_, _25954_);
  nor _45302_ (_29605_, _29583_, _25954_);
  or _45303_ (_29616_, _29605_, _29594_);
  and _45304_ (_29627_, _29616_, _26228_);
  nor _45305_ (_29638_, _26733_, _26722_);
  nor _45306_ (_29648_, _29638_, _26744_);
  nor _45307_ (_29659_, _29648_, _26316_);
  nor _45308_ (_29670_, _29659_, _29627_);
  and _45309_ (_29681_, _29670_, _29561_);
  not _45310_ (_29692_, _29681_);
  nor _45311_ (_29703_, _29692_, _29232_);
  and _45312_ (_29714_, _29703_, _29221_);
  not _45313_ (_29725_, _29714_);
  or _45314_ (_29736_, _29725_, _25148_);
  not _45315_ (_29747_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _45316_ (_29758_, _25148_, _29747_);
  and _45317_ (_29769_, _29758_, _27918_);
  and _45318_ (_29790_, _29769_, _29736_);
  nor _45319_ (_29791_, _27896_, _29747_);
  not _45320_ (_29802_, _24265_);
  and _45321_ (_29813_, _29802_, _24138_);
  and _45322_ (_29824_, _29813_, _24018_);
  and _45323_ (_29835_, _29824_, _25147_);
  or _45324_ (_29846_, _29835_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _45325_ (_29857_, _29846_, _28576_);
  nand _45326_ (_29868_, _29835_, _28510_);
  and _45327_ (_29879_, _29868_, _29857_);
  or _45328_ (_29890_, _29879_, _29791_);
  or _45329_ (_29901_, _29890_, _29790_);
  and _45330_ (_08943_, _29901_, _41755_);
  and _45331_ (_29922_, _23445_, _20924_);
  not _45332_ (_29933_, _29922_);
  and _45333_ (_29944_, _20711_, _15573_);
  nor _45334_ (_29954_, _27227_, _15967_);
  nor _45335_ (_29965_, _29254_, _25910_);
  nor _45336_ (_29976_, _26952_, _27029_);
  nor _45337_ (_29987_, _29976_, _29965_);
  and _45338_ (_29998_, _29987_, _18872_);
  nor _45339_ (_30009_, _29987_, _18872_);
  nor _45340_ (_30020_, _30009_, _29998_);
  and _45341_ (_30031_, _30020_, _26941_);
  nor _45342_ (_30042_, _30031_, _29954_);
  nor _45343_ (_30053_, _26744_, _26689_);
  nor _45344_ (_30064_, _30053_, _26755_);
  nor _45345_ (_30075_, _30064_, _26316_);
  and _45346_ (_30096_, _27479_, _25388_);
  nor _45347_ (_30097_, _27457_, _25377_);
  not _45348_ (_30108_, _30097_);
  and _45349_ (_30119_, _27621_, _25366_);
  and _45350_ (_30130_, _27643_, _18861_);
  nor _45351_ (_30141_, _30130_, _30119_);
  nand _45352_ (_30152_, _30141_, _30108_);
  nor _45353_ (_30163_, _30152_, _30096_);
  nor _45354_ (_30174_, _27533_, _18687_);
  not _45355_ (_30185_, _30174_);
  nor _45356_ (_30196_, _27687_, _18861_);
  nor _45357_ (_30207_, _28816_, _18339_);
  nor _45358_ (_30218_, _30207_, _30196_);
  and _45359_ (_30229_, _30218_, _30185_);
  and _45360_ (_30240_, _30229_, _30163_);
  not _45361_ (_30251_, _30240_);
  nor _45362_ (_30262_, _30251_, _30075_);
  nor _45363_ (_30272_, _25987_, _25965_);
  nor _45364_ (_30283_, _30272_, _26239_);
  and _45365_ (_30294_, _30283_, _26009_);
  nor _45366_ (_30305_, _29363_, _18861_);
  and _45367_ (_30316_, _27051_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45368_ (_30327_, _30316_, _30305_);
  nor _45369_ (_30338_, _30327_, _28082_);
  nor _45370_ (_30349_, _30338_, _30294_);
  and _45371_ (_30360_, _30349_, _30262_);
  and _45372_ (_30371_, _30360_, _30042_);
  not _45373_ (_30382_, _30371_);
  nor _45374_ (_30393_, _30382_, _29944_);
  and _45375_ (_30404_, _30393_, _29933_);
  not _45376_ (_30425_, _30404_);
  or _45377_ (_30426_, _30425_, _25148_);
  not _45378_ (_30437_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _45379_ (_30448_, _25148_, _30437_);
  and _45380_ (_30459_, _30448_, _27918_);
  and _45381_ (_30470_, _30459_, _30426_);
  nor _45382_ (_30481_, _27896_, _30437_);
  nand _45383_ (_30493_, _25147_, _24018_);
  or _45384_ (_30514_, _28532_, _30493_);
  and _45385_ (_30525_, _30514_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _45386_ (_30536_, _24138_);
  and _45387_ (_30547_, _24018_, _24265_);
  and _45388_ (_30558_, _30547_, _30536_);
  not _45389_ (_30569_, _30558_);
  nor _45390_ (_30580_, _30569_, _28510_);
  and _45391_ (_30590_, _24018_, _24138_);
  and _45392_ (_30601_, _30590_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _45393_ (_30612_, _30601_, _30580_);
  and _45394_ (_30623_, _30612_, _25147_);
  or _45395_ (_30634_, _30623_, _30525_);
  and _45396_ (_30645_, _30634_, _28576_);
  or _45397_ (_30656_, _30645_, _30481_);
  or _45398_ (_30667_, _30656_, _30470_);
  and _45399_ (_08954_, _30667_, _41755_);
  and _45400_ (_30688_, _20754_, _15573_);
  not _45401_ (_30699_, _30688_);
  and _45402_ (_30710_, _23510_, _20924_);
  nor _45403_ (_30721_, _26755_, _26656_);
  nor _45404_ (_30732_, _30721_, _26766_);
  nor _45405_ (_30743_, _30732_, _26316_);
  not _45406_ (_30754_, _30743_);
  and _45407_ (_30765_, _26009_, _25518_);
  or _45408_ (_30776_, _30765_, _26239_);
  nor _45409_ (_30787_, _30776_, _26020_);
  not _45410_ (_30798_, _30787_);
  nor _45411_ (_30809_, _27227_, _16966_);
  nor _45412_ (_30820_, _27062_, _25910_);
  nor _45413_ (_30831_, _26963_, _27029_);
  nor _45414_ (_30842_, _30831_, _30820_);
  and _45415_ (_30853_, _30842_, _18350_);
  not _45416_ (_30864_, _26941_);
  nor _45417_ (_30875_, _30842_, _18350_);
  or _45418_ (_30886_, _30875_, _30864_);
  nor _45419_ (_30896_, _30886_, _30853_);
  nor _45420_ (_30917_, _30896_, _30809_);
  and _45421_ (_30918_, _27479_, _25365_);
  and _45422_ (_30929_, _27621_, _25333_);
  nor _45423_ (_30940_, _27457_, _25344_);
  and _45424_ (_30951_, _27643_, _18339_);
  or _45425_ (_30962_, _30951_, _30940_);
  or _45426_ (_30973_, _30962_, _30929_);
  nor _45427_ (_30984_, _30973_, _30918_);
  not _45428_ (_30995_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45429_ (_31006_, _27051_, _30995_);
  nor _45430_ (_31016_, _31006_, _18350_);
  not _45431_ (_31027_, _31016_);
  nor _45432_ (_31038_, _27281_, _28082_);
  and _45433_ (_31049_, _31038_, _31027_);
  nor _45434_ (_31060_, _27687_, _18339_);
  not _45435_ (_31071_, _31060_);
  nor _45436_ (_31082_, _28816_, _18001_);
  nor _45437_ (_31093_, _27533_, _18861_);
  nor _45438_ (_31104_, _31093_, _31082_);
  and _45439_ (_31115_, _31104_, _31071_);
  not _45440_ (_31126_, _31115_);
  nor _45441_ (_31146_, _31126_, _31049_);
  and _45442_ (_31147_, _31146_, _30984_);
  and _45443_ (_31158_, _31147_, _30917_);
  and _45444_ (_31169_, _31158_, _30798_);
  and _45445_ (_31180_, _31169_, _30754_);
  not _45446_ (_31191_, _31180_);
  nor _45447_ (_31202_, _31191_, _30710_);
  and _45448_ (_31213_, _31202_, _30699_);
  not _45449_ (_31224_, _31213_);
  or _45450_ (_31235_, _31224_, _25148_);
  not _45451_ (_31246_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _45452_ (_31257_, _25148_, _31246_);
  and _45453_ (_31268_, _31257_, _27918_);
  and _45454_ (_31278_, _31268_, _31235_);
  nor _45455_ (_31289_, _27896_, _31246_);
  and _45456_ (_31300_, _30493_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _45457_ (_31311_, _28532_, _24018_);
  not _45458_ (_31322_, _31311_);
  nor _45459_ (_31333_, _31322_, _28510_);
  nor _45460_ (_31344_, _30590_, _30547_);
  nor _45461_ (_31355_, _31344_, _31246_);
  or _45462_ (_31366_, _31355_, _31333_);
  and _45463_ (_31377_, _31366_, _25147_);
  or _45464_ (_31388_, _31377_, _31300_);
  and _45465_ (_31398_, _31388_, _28576_);
  or _45466_ (_31409_, _31398_, _31289_);
  or _45467_ (_31420_, _31409_, _31278_);
  and _45468_ (_08965_, _31420_, _41755_);
  and _45469_ (_31441_, _23574_, _20924_);
  not _45470_ (_31452_, _31441_);
  and _45471_ (_31463_, _20785_, _15573_);
  nor _45472_ (_31474_, _26832_, _25322_);
  and _45473_ (_31485_, _26832_, _25322_);
  nor _45474_ (_31496_, _31485_, _31474_);
  and _45475_ (_31507_, _31496_, _26305_);
  not _45476_ (_31518_, _31507_);
  nor _45477_ (_31528_, _26053_, _25322_);
  nor _45478_ (_31539_, _31528_, _26064_);
  and _45479_ (_31550_, _31539_, _26228_);
  and _45480_ (_31561_, _25910_, _18012_);
  nor _45481_ (_31572_, _25910_, _16131_);
  or _45482_ (_31583_, _31572_, _31561_);
  and _45483_ (_31594_, _31583_, _27216_);
  and _45484_ (_31605_, _26974_, _25910_);
  and _45485_ (_31616_, _27073_, _27029_);
  nor _45486_ (_31627_, _31616_, _31605_);
  nor _45487_ (_31638_, _31627_, _18001_);
  not _45488_ (_31648_, _31638_);
  and _45489_ (_31659_, _31627_, _18001_);
  nor _45490_ (_31670_, _31659_, _30864_);
  and _45491_ (_31681_, _31670_, _31648_);
  nor _45492_ (_31692_, _31681_, _31594_);
  nor _45493_ (_31703_, _27292_, _18012_);
  not _45494_ (_31724_, _31703_);
  nor _45495_ (_31725_, _27303_, _28082_);
  and _45496_ (_31736_, _31725_, _31724_);
  not _45497_ (_31747_, _31736_);
  and _45498_ (_31758_, _27479_, _25322_);
  nor _45499_ (_31769_, _27457_, _25312_);
  not _45500_ (_31779_, _31769_);
  and _45501_ (_31790_, _27621_, _25268_);
  and _45502_ (_31801_, _27643_, _18001_);
  nor _45503_ (_31812_, _31801_, _31790_);
  nand _45504_ (_31823_, _31812_, _31779_);
  nor _45505_ (_31834_, _31823_, _31758_);
  nor _45506_ (_31845_, _28816_, _17826_);
  not _45507_ (_31856_, _31845_);
  nor _45508_ (_31867_, _27687_, _18001_);
  nor _45509_ (_31878_, _27533_, _18339_);
  nor _45510_ (_31888_, _31878_, _31867_);
  and _45511_ (_31899_, _31888_, _31856_);
  and _45512_ (_31910_, _31899_, _31834_);
  and _45513_ (_31921_, _31910_, _31747_);
  and _45514_ (_31932_, _31921_, _31692_);
  not _45515_ (_31943_, _31932_);
  nor _45516_ (_31954_, _31943_, _31550_);
  and _45517_ (_31965_, _31954_, _31518_);
  not _45518_ (_31976_, _31965_);
  nor _45519_ (_31987_, _31976_, _31463_);
  and _45520_ (_31997_, _31987_, _31452_);
  not _45521_ (_32008_, _31997_);
  or _45522_ (_32019_, _32008_, _25148_);
  not _45523_ (_32030_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _45524_ (_32041_, _25148_, _32030_);
  and _45525_ (_32052_, _32041_, _27918_);
  and _45526_ (_32063_, _32052_, _32019_);
  nor _45527_ (_32074_, _27896_, _32030_);
  not _45528_ (_32085_, _25147_);
  and _45529_ (_32096_, _24276_, _28521_);
  nor _45530_ (_32106_, _24276_, _28521_);
  nor _45531_ (_32117_, _32106_, _32096_);
  or _45532_ (_32128_, _32117_, _32085_);
  and _45533_ (_32139_, _32128_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _45534_ (_32150_, _32096_, _29134_);
  and _45535_ (_32161_, _32106_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _45536_ (_32172_, _32161_, _32150_);
  and _45537_ (_32183_, _32172_, _25147_);
  or _45538_ (_32194_, _32183_, _32139_);
  and _45539_ (_32205_, _32194_, _28576_);
  or _45540_ (_32215_, _32205_, _32074_);
  or _45541_ (_32226_, _32215_, _32063_);
  and _45542_ (_08976_, _32226_, _41755_);
  and _45543_ (_32247_, _23660_, _20924_);
  not _45544_ (_32258_, _32247_);
  and _45545_ (_32269_, _20828_, _15573_);
  nor _45546_ (_32280_, _26843_, _26492_);
  nor _45547_ (_32291_, _32280_, _26854_);
  nor _45548_ (_32302_, _32291_, _26316_);
  not _45549_ (_32313_, _32302_);
  nor _45550_ (_32324_, _25268_, _25257_);
  or _45551_ (_32334_, _32324_, _25279_);
  and _45552_ (_32355_, _32334_, _26064_);
  nor _45553_ (_32356_, _32334_, _26064_);
  or _45554_ (_32367_, _32356_, _32355_);
  and _45555_ (_32378_, _32367_, _26228_);
  nor _45556_ (_32389_, _25910_, _17119_);
  and _45557_ (_32400_, _25910_, _17837_);
  nor _45558_ (_32411_, _32400_, _32389_);
  nor _45559_ (_32422_, _32411_, _27227_);
  nor _45560_ (_32433_, _26985_, _27029_);
  nor _45561_ (_32443_, _27084_, _25910_);
  nor _45562_ (_32454_, _32443_, _32433_);
  and _45563_ (_32465_, _32454_, _17837_);
  nor _45564_ (_32476_, _32454_, _17837_);
  or _45565_ (_32487_, _32476_, _30864_);
  nor _45566_ (_32498_, _32487_, _32465_);
  nor _45567_ (_32509_, _32498_, _32422_);
  not _45568_ (_32520_, _27358_);
  and _45569_ (_32531_, _32520_, _27314_);
  nor _45570_ (_32542_, _27358_, _27303_);
  nor _45571_ (_32552_, _32542_, _17826_);
  nor _45572_ (_32563_, _32552_, _32531_);
  nor _45573_ (_32574_, _32563_, _28082_);
  and _45574_ (_32585_, _27479_, _25257_);
  and _45575_ (_32596_, _27621_, _25235_);
  nor _45576_ (_32607_, _27457_, _25246_);
  and _45577_ (_32618_, _27643_, _17826_);
  or _45578_ (_32629_, _32618_, _32607_);
  or _45579_ (_32640_, _32629_, _32596_);
  nor _45580_ (_32660_, _32640_, _32585_);
  nor _45581_ (_32661_, _28816_, _16790_);
  nor _45582_ (_32672_, _27533_, _18001_);
  nor _45583_ (_32683_, _27687_, _17826_);
  or _45584_ (_32694_, _32683_, _32672_);
  nor _45585_ (_32705_, _32694_, _32661_);
  and _45586_ (_32716_, _32705_, _32660_);
  not _45587_ (_32727_, _32716_);
  nor _45588_ (_32738_, _32727_, _32574_);
  and _45589_ (_32749_, _32738_, _32509_);
  not _45590_ (_32760_, _32749_);
  nor _45591_ (_32770_, _32760_, _32378_);
  and _45592_ (_32781_, _32770_, _32313_);
  not _45593_ (_32792_, _32781_);
  nor _45594_ (_32803_, _32792_, _32269_);
  and _45595_ (_32814_, _32803_, _32258_);
  not _45596_ (_32825_, _32814_);
  or _45597_ (_32836_, _32825_, _25148_);
  not _45598_ (_32847_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _45599_ (_32858_, _25148_, _32847_);
  and _45600_ (_32869_, _32858_, _27918_);
  and _45601_ (_32879_, _32869_, _32836_);
  nor _45602_ (_32890_, _27896_, _32847_);
  and _45603_ (_32901_, _29813_, _28521_);
  and _45604_ (_32912_, _32901_, _25147_);
  nand _45605_ (_32923_, _32912_, _28510_);
  or _45606_ (_32934_, _32912_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _45607_ (_32945_, _32934_, _28576_);
  and _45608_ (_32956_, _32945_, _32923_);
  or _45609_ (_32967_, _32956_, _32890_);
  or _45610_ (_32978_, _32967_, _32879_);
  and _45611_ (_08987_, _32978_, _41755_);
  and _45612_ (_33008_, _23725_, _20924_);
  not _45613_ (_33009_, _33008_);
  and _45614_ (_33020_, _20859_, _15573_);
  nor _45615_ (_33031_, _26854_, _26459_);
  nor _45616_ (_33042_, _33031_, _26865_);
  nor _45617_ (_33053_, _33042_, _26316_);
  not _45618_ (_33064_, _33053_);
  nor _45619_ (_33075_, _26097_, _26085_);
  not _45620_ (_33086_, _33075_);
  nor _45621_ (_33097_, _26239_, _26108_);
  and _45622_ (_33107_, _33097_, _33086_);
  nor _45623_ (_33118_, _25910_, _26327_);
  or _45624_ (_33129_, _33118_, _27227_);
  nor _45625_ (_33140_, _33129_, _28049_);
  nor _45626_ (_33151_, _25910_, _17837_);
  nand _45627_ (_33162_, _33151_, _27084_);
  nand _45628_ (_33173_, _26996_, _25910_);
  and _45629_ (_33184_, _33173_, _33162_);
  and _45630_ (_33195_, _33184_, _16790_);
  nor _45631_ (_33206_, _33184_, _16790_);
  or _45632_ (_33216_, _33206_, _30864_);
  nor _45633_ (_33227_, _33216_, _33195_);
  nor _45634_ (_33238_, _33227_, _33140_);
  nor _45635_ (_33249_, _32531_, _16790_);
  and _45636_ (_33260_, _32531_, _16790_);
  nor _45637_ (_33271_, _33260_, _33249_);
  nor _45638_ (_33282_, _33271_, _28082_);
  nor _45639_ (_33293_, _27457_, _25203_);
  and _45640_ (_33304_, _27479_, _25214_);
  nor _45641_ (_33315_, _33304_, _33293_);
  and _45642_ (_33325_, _27621_, _25192_);
  and _45643_ (_33336_, _27643_, _16790_);
  nor _45644_ (_33347_, _33336_, _33325_);
  nor _45645_ (_33358_, _27687_, _16790_);
  not _45646_ (_33379_, _33358_);
  nor _45647_ (_33380_, _28816_, _17630_);
  nor _45648_ (_33391_, _27533_, _17826_);
  nor _45649_ (_33402_, _33391_, _33380_);
  and _45650_ (_33413_, _33402_, _33379_);
  and _45651_ (_33424_, _33413_, _33347_);
  and _45652_ (_33434_, _33424_, _33315_);
  not _45653_ (_33445_, _33434_);
  nor _45654_ (_33456_, _33445_, _33282_);
  and _45655_ (_33467_, _33456_, _33238_);
  not _45656_ (_33478_, _33467_);
  nor _45657_ (_33489_, _33478_, _33107_);
  and _45658_ (_33500_, _33489_, _33064_);
  not _45659_ (_33511_, _33500_);
  nor _45660_ (_33522_, _33511_, _33020_);
  and _45661_ (_33533_, _33522_, _33009_);
  not _45662_ (_33543_, _33533_);
  or _45663_ (_33554_, _33543_, _25148_);
  not _45664_ (_33565_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _45665_ (_33576_, _25148_, _33565_);
  and _45666_ (_33587_, _33576_, _27918_);
  and _45667_ (_33598_, _33587_, _33554_);
  nor _45668_ (_33609_, _27896_, _33565_);
  nor _45669_ (_33620_, _24018_, _24138_);
  and _45670_ (_33631_, _33620_, _24265_);
  and _45671_ (_33642_, _33631_, _25147_);
  nand _45672_ (_33652_, _33642_, _28510_);
  or _45673_ (_33663_, _33642_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _45674_ (_33674_, _33663_, _28576_);
  and _45675_ (_33685_, _33674_, _33652_);
  or _45676_ (_33696_, _33685_, _33609_);
  or _45677_ (_33707_, _33696_, _33598_);
  and _45678_ (_08998_, _33707_, _41755_);
  and _45679_ (_33728_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45680_ (_33739_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor _45681_ (_33750_, _33739_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _45682_ (_33760_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _45683_ (_33771_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _45684_ (_33782_, _33771_, _33760_);
  and _45685_ (_33793_, _33739_, _15507_);
  and _45686_ (_33804_, _33793_, _33782_);
  not _45687_ (_33815_, _33804_);
  and _45688_ (_33826_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _45689_ (_33837_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45690_ (_33848_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _45691_ (_33859_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45692_ (_33870_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _45693_ (_33880_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not _45694_ (_33901_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45695_ (_33902_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _33901_);
  and _45696_ (_33913_, _33902_, _33880_);
  and _45697_ (_33924_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not _45698_ (_33935_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _45699_ (_33946_, _33935_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45700_ (_33957_, _33946_, _33880_);
  and _45701_ (_33968_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _45702_ (_33979_, _33968_, _33924_);
  nor _45703_ (_33989_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _45704_ (_34000_, _33989_, _33880_);
  and _45705_ (_34011_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _45706_ (_34022_, _33989_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45707_ (_34033_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _45708_ (_34044_, _34033_, _34011_);
  and _45709_ (_34055_, _33989_, _33880_);
  and _45710_ (_34066_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _45711_ (_34077_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45712_ (_34088_, _34077_, _33880_);
  and _45713_ (_34098_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _45714_ (_34109_, _34098_, _34066_);
  and _45715_ (_34120_, _34109_, _34044_);
  and _45716_ (_34131_, _34120_, _33979_);
  nor _45717_ (_34142_, _34131_, _33870_);
  and _45718_ (_34153_, _34142_, _33859_);
  or _45719_ (_34173_, _34153_, _33848_);
  and _45720_ (_34174_, _34173_, _33837_);
  nor _45721_ (_34185_, _34174_, _33826_);
  nor _45722_ (_34196_, _34185_, _33815_);
  and _45723_ (_34207_, _33782_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _45724_ (_34218_, _34207_, _33815_);
  nor _45725_ (_34229_, _34218_, _34196_);
  not _45726_ (_34240_, _34229_);
  not _45727_ (_34251_, _33870_);
  and _45728_ (_34262_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _45729_ (_34273_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _45730_ (_34284_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _45731_ (_34294_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _45732_ (_34305_, _34294_, _34284_);
  and _45733_ (_34316_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _45734_ (_34327_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _45735_ (_34338_, _34327_, _34316_);
  nand _45736_ (_34349_, _34338_, _34305_);
  or _45737_ (_34360_, _34349_, _34273_);
  nor _45738_ (_34371_, _34360_, _34262_);
  and _45739_ (_34382_, _34371_, _34251_);
  and _45740_ (_34393_, _34382_, _33859_);
  nor _45741_ (_34404_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _33859_);
  nor _45742_ (_34414_, _34404_, _34393_);
  nor _45743_ (_34425_, _34414_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45744_ (_34436_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _33837_);
  nor _45745_ (_34447_, _34436_, _34425_);
  and _45746_ (_34458_, _34447_, _33804_);
  and _45747_ (_34469_, _33782_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _45748_ (_34480_, _34469_, _33815_);
  nor _45749_ (_34491_, _34480_, _34458_);
  not _45750_ (_34502_, _34491_);
  and _45751_ (_34513_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45752_ (_34524_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or _45753_ (_34534_, _33870_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45754_ (_34545_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _45755_ (_34556_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _45756_ (_34567_, _34556_, _34545_);
  and _45757_ (_34578_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _45758_ (_34589_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _45759_ (_34600_, _34589_, _34578_);
  and _45760_ (_34611_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _45761_ (_34622_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _45762_ (_34633_, _34622_, _34611_);
  and _45763_ (_34644_, _34633_, _34600_);
  and _45764_ (_34654_, _34644_, _34567_);
  nor _45765_ (_34665_, _34654_, _34534_);
  nor _45766_ (_34676_, _34665_, _34524_);
  nor _45767_ (_34687_, _34676_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45768_ (_34698_, _34687_, _34513_);
  nor _45769_ (_34709_, _34698_, _33815_);
  and _45770_ (_34720_, _33782_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _45771_ (_34731_, _34720_, _33815_);
  nor _45772_ (_34742_, _34731_, _34709_);
  and _45773_ (_34753_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45774_ (_34764_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45775_ (_34775_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _45776_ (_34795_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _45777_ (_34796_, _34795_, _34775_);
  and _45778_ (_34807_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _45779_ (_34818_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _45780_ (_34829_, _34818_, _34807_);
  and _45781_ (_34840_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _45782_ (_34851_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _45783_ (_34862_, _34851_, _34840_);
  and _45784_ (_34873_, _34862_, _34829_);
  and _45785_ (_34884_, _34873_, _34796_);
  nor _45786_ (_34895_, _34884_, _33870_);
  and _45787_ (_34906_, _34895_, _33859_);
  or _45788_ (_34916_, _34906_, _34764_);
  and _45789_ (_34927_, _34916_, _33837_);
  nor _45790_ (_34938_, _34927_, _34753_);
  nor _45791_ (_34949_, _34938_, _33815_);
  and _45792_ (_34960_, _33782_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _45793_ (_34971_, _34960_, _33815_);
  nor _45794_ (_34982_, _34971_, _34949_);
  and _45795_ (_34993_, _34982_, _34742_);
  and _45796_ (_35004_, _34993_, _34502_);
  and _45797_ (_35015_, _35004_, _34240_);
  and _45798_ (_35026_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _45799_ (_35037_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _45800_ (_35048_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _45801_ (_35059_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _45802_ (_35070_, _35059_, _35048_);
  and _45803_ (_35081_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _45804_ (_35092_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _45805_ (_35103_, _35092_, _35081_);
  nand _45806_ (_35114_, _35103_, _35070_);
  or _45807_ (_35125_, _35114_, _35037_);
  nor _45808_ (_35136_, _35125_, _35026_);
  and _45809_ (_35147_, _35136_, _34251_);
  and _45810_ (_35158_, _35147_, _33859_);
  nor _45811_ (_35169_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _33859_);
  nor _45812_ (_35180_, _35169_, _35158_);
  nor _45813_ (_35191_, _35180_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45814_ (_35202_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _33837_);
  nor _45815_ (_35213_, _35202_, _35191_);
  and _45816_ (_35224_, _35213_, _33804_);
  and _45817_ (_35235_, _33782_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _45818_ (_35246_, _35235_, _33815_);
  nor _45819_ (_35257_, _35246_, _35224_);
  and _45820_ (_35268_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45821_ (_35279_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45822_ (_35290_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _45823_ (_35301_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _45824_ (_35312_, _35301_, _35290_);
  and _45825_ (_35323_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _45826_ (_35334_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _45827_ (_35345_, _35334_, _35323_);
  and _45828_ (_35356_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _45829_ (_35367_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _45830_ (_35378_, _35367_, _35356_);
  and _45831_ (_35389_, _35378_, _35345_);
  and _45832_ (_35400_, _35389_, _35312_);
  nor _45833_ (_35411_, _35400_, _33870_);
  and _45834_ (_35422_, _35411_, _33859_);
  or _45835_ (_35433_, _35422_, _35279_);
  and _45836_ (_35444_, _35433_, _33837_);
  nor _45837_ (_35455_, _35444_, _35268_);
  nor _45838_ (_35466_, _35455_, _33815_);
  and _45839_ (_35477_, _33782_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _45840_ (_35488_, _35477_, _33815_);
  nor _45841_ (_35510_, _35488_, _35466_);
  not _45842_ (_35511_, _35510_);
  and _45843_ (_35533_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45844_ (_35534_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45845_ (_35556_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _45846_ (_35557_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _45847_ (_35579_, _35557_, _35556_);
  and _45848_ (_35580_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _45849_ (_35591_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _45850_ (_35602_, _35591_, _35580_);
  and _45851_ (_35613_, _35602_, _35579_);
  and _45852_ (_35624_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _45853_ (_35635_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _45854_ (_35646_, _35635_, _35624_);
  and _45855_ (_35657_, _35646_, _35613_);
  nor _45856_ (_35668_, _35657_, _34534_);
  or _45857_ (_35679_, _35668_, _35534_);
  and _45858_ (_35690_, _35679_, _33837_);
  nor _45859_ (_35701_, _35690_, _35533_);
  nor _45860_ (_35712_, _35701_, _33815_);
  and _45861_ (_35723_, _33782_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _45862_ (_35734_, _35723_, _33815_);
  nor _45863_ (_35745_, _35734_, _35712_);
  and _45864_ (_35756_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and _45865_ (_35767_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _45866_ (_35778_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _45867_ (_35789_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _45868_ (_35800_, _35789_, _35778_);
  and _45869_ (_35811_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _45870_ (_35822_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _45871_ (_35833_, _35822_, _35811_);
  and _45872_ (_35844_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _45873_ (_35855_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _45874_ (_35866_, _35855_, _35844_);
  and _45875_ (_35877_, _35866_, _35833_);
  and _45876_ (_35888_, _35877_, _35800_);
  nor _45877_ (_35899_, _35888_, _34534_);
  nor _45878_ (_35910_, _35899_, _35767_);
  nor _45879_ (_35921_, _35910_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45880_ (_35932_, _35921_, _35756_);
  nor _45881_ (_35943_, _35932_, _33815_);
  and _45882_ (_35954_, _33782_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _45883_ (_35965_, _35954_, _33815_);
  nor _45884_ (_35976_, _35965_, _35943_);
  not _45885_ (_35987_, _35976_);
  and _45886_ (_35998_, _35987_, _35745_);
  and _45887_ (_36009_, _35998_, _35511_);
  and _45888_ (_36020_, _36009_, _35257_);
  and _45889_ (_36031_, _36020_, _35015_);
  not _45890_ (_36042_, _35257_);
  and _45891_ (_36053_, _35745_, _35510_);
  and _45892_ (_36064_, _36053_, _35987_);
  and _45893_ (_36075_, _36064_, _36042_);
  nor _45894_ (_36086_, _35745_, _35510_);
  and _45895_ (_36097_, _36086_, _35976_);
  and _45896_ (_36108_, _36097_, _36042_);
  or _45897_ (_36119_, _36108_, _36075_);
  nand _45898_ (_36130_, _36119_, _35015_);
  not _45899_ (_36141_, _36130_);
  nor _45900_ (_36152_, _36141_, _36031_);
  and _45901_ (_36163_, _34229_, _34491_);
  and _45902_ (_36174_, _36163_, _34993_);
  not _45903_ (_36185_, _35745_);
  and _45904_ (_36196_, _36185_, _35510_);
  and _45905_ (_36207_, _36196_, _35987_);
  and _45906_ (_36218_, _36207_, _36042_);
  and _45907_ (_36229_, _36218_, _36174_);
  nor _45908_ (_36240_, _34742_, _34491_);
  and _45909_ (_36251_, _36240_, _34982_);
  and _45910_ (_36262_, _35257_, _36251_);
  and _45911_ (_36273_, _36064_, _36262_);
  nor _45912_ (_36284_, _36273_, _36229_);
  and _45913_ (_36295_, _35976_, _36185_);
  and _45914_ (_36306_, _36295_, _35510_);
  and _45915_ (_36317_, _36306_, _36262_);
  and _45916_ (_36328_, _36086_, _35987_);
  and _45917_ (_36339_, _36328_, _36262_);
  nor _45918_ (_36350_, _36339_, _36317_);
  and _45919_ (_36361_, _35004_, _34229_);
  and _45920_ (_36372_, _35976_, _35745_);
  and _45921_ (_36383_, _36372_, _35511_);
  and _45922_ (_36394_, _36383_, _36361_);
  and _45923_ (_36405_, _36097_, _36262_);
  nor _45924_ (_36416_, _36405_, _36394_);
  and _45925_ (_36427_, _36416_, _36350_);
  and _45926_ (_36437_, _36427_, _36284_);
  and _45927_ (_36448_, _36207_, _36251_);
  not _45928_ (_36459_, _34982_);
  nor _45929_ (_36470_, _35257_, _36459_);
  and _45930_ (_36481_, _36470_, _36240_);
  and _45931_ (_36492_, _36064_, _36481_);
  nor _45932_ (_36503_, _36492_, _36448_);
  and _45933_ (_36514_, _36372_, _35510_);
  and _45934_ (_36525_, _36514_, _36251_);
  and _45935_ (_36536_, _36009_, _36481_);
  nor _45936_ (_36547_, _36536_, _36525_);
  not _45937_ (_36557_, _36547_);
  nor _45938_ (_36568_, _35257_, _35511_);
  and _45939_ (_36579_, _36568_, _36295_);
  and _45940_ (_36590_, _36579_, _36251_);
  and _45941_ (_36601_, _36383_, _36251_);
  or _45942_ (_36612_, _36601_, _36590_);
  nor _45943_ (_36623_, _36612_, _36557_);
  and _45944_ (_36634_, _36623_, _36503_);
  and _45945_ (_36645_, _36634_, _36437_);
  and _45946_ (_36656_, _36645_, _36152_);
  nor _45947_ (_36667_, _36656_, _33750_);
  not _45948_ (_36678_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _45949_ (_36689_, _15507_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45950_ (_36700_, _36689_, _36678_);
  and _45951_ (_36711_, _36700_, _36097_);
  and _45952_ (_36722_, _36711_, _36174_);
  and _45953_ (_36733_, _36394_, _36689_);
  and _45954_ (_36744_, _36733_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or _45955_ (_36755_, _36744_, _36722_);
  nor _45956_ (_36766_, _36755_, _36667_);
  nor _45957_ (_36777_, _36766_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45958_ (_36788_, _36777_, _33728_);
  and _45959_ (_36798_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _45960_ (_36809_, _36009_, _36262_);
  not _45961_ (_36820_, _36809_);
  not _45962_ (_36831_, _34742_);
  and _45963_ (_36842_, _34982_, _36831_);
  and _45964_ (_36853_, _34240_, _34491_);
  and _45965_ (_36864_, _36853_, _36842_);
  and _45966_ (_36875_, _36328_, _35257_);
  and _45967_ (_36886_, _36875_, _36864_);
  and _45968_ (_36897_, _35998_, _36042_);
  and _45969_ (_36907_, _36897_, _36864_);
  nor _45970_ (_36918_, _36907_, _36886_);
  and _45971_ (_36929_, _36918_, _36820_);
  and _45972_ (_36940_, _36174_, _36207_);
  and _45973_ (_36951_, _36097_, _35257_);
  and _45974_ (_36962_, _35004_, _36951_);
  nor _45975_ (_36973_, _36962_, _36940_);
  not _45976_ (_36984_, _36394_);
  and _45977_ (_36995_, _35257_, _36459_);
  and _45978_ (_37006_, _36995_, _36009_);
  and _45979_ (_37016_, _35257_, _36514_);
  and _45980_ (_37027_, _37016_, _36864_);
  nor _45981_ (_37038_, _37027_, _37006_);
  and _45982_ (_37049_, _37038_, _36984_);
  and _45983_ (_37060_, _37049_, _36973_);
  nor _45984_ (_37071_, _36579_, _36383_);
  not _45985_ (_37082_, _36864_);
  nor _45986_ (_37093_, _37082_, _37071_);
  and _45987_ (_37104_, _36174_, _36383_);
  and _45988_ (_37115_, _37104_, _35257_);
  and _45989_ (_37126_, _36383_, _36042_);
  and _45990_ (_37136_, _36568_, _36372_);
  or _45991_ (_37147_, _37136_, _37126_);
  and _45992_ (_37158_, _37147_, _36174_);
  nor _45993_ (_37169_, _37158_, _37115_);
  not _45994_ (_37180_, _37169_);
  nor _45995_ (_37191_, _37180_, _37093_);
  and _45996_ (_37202_, _37191_, _37060_);
  and _45997_ (_37213_, _37202_, _36929_);
  and _45998_ (_37224_, _36306_, _35257_);
  and _45999_ (_37235_, _37224_, _35004_);
  not _46000_ (_37246_, _37235_);
  and _46001_ (_37257_, _37136_, _36864_);
  and _46002_ (_37268_, _36009_, _36042_);
  and _46003_ (_37279_, _36174_, _37268_);
  nor _46004_ (_37290_, _37279_, _37257_);
  and _46005_ (_37301_, _37290_, _37246_);
  and _46006_ (_37310_, _36108_, _36361_);
  and _46007_ (_37318_, _36864_, _36218_);
  nor _46008_ (_37326_, _37318_, _37310_);
  and _46009_ (_37333_, _37326_, _37301_);
  and _46010_ (_37341_, _36020_, _36174_);
  and _46011_ (_37349_, _37224_, _36864_);
  nor _46012_ (_37356_, _37349_, _37341_);
  and _46013_ (_37364_, _36361_, _37268_);
  and _46014_ (_37372_, _36207_, _35257_);
  and _46015_ (_37373_, _37372_, _36361_);
  nor _46016_ (_37374_, _37373_, _37364_);
  and _46017_ (_37376_, _37374_, _37356_);
  and _46018_ (_37387_, _37376_, _37333_);
  and _46019_ (_37398_, _36864_, _36951_);
  and _46020_ (_37409_, _37372_, _36864_);
  nor _46021_ (_37420_, _37409_, _37398_);
  and _46022_ (_37431_, _36064_, _35257_);
  and _46023_ (_37442_, _37431_, _36361_);
  and _46024_ (_37453_, _36579_, _35004_);
  nor _46025_ (_37464_, _37453_, _37442_);
  and _46026_ (_37475_, _37464_, _37420_);
  and _46027_ (_37486_, _36020_, _36361_);
  and _46028_ (_37497_, _36218_, _36361_);
  nor _46029_ (_37508_, _37497_, _37486_);
  and _46030_ (_37519_, _36075_, _36361_);
  and _46031_ (_37530_, _36864_, _37431_);
  nor _46032_ (_37541_, _37530_, _37519_);
  and _46033_ (_37552_, _37541_, _37508_);
  and _46034_ (_37563_, _37552_, _37475_);
  and _46035_ (_37574_, _37563_, _37387_);
  and _46036_ (_37580_, _37574_, _37213_);
  nor _46037_ (_37591_, _37580_, _33750_);
  and _46038_ (_37602_, _36689_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _46039_ (_37613_, _37602_, _36394_);
  not _46040_ (_37624_, _37613_);
  and _46041_ (_37635_, _36174_, _36295_);
  and _46042_ (_37646_, _37635_, _36700_);
  not _46043_ (_37657_, _36700_);
  and _46044_ (_37668_, _36383_, _35257_);
  and _46045_ (_37679_, _37668_, _36174_);
  and _46046_ (_37690_, _37136_, _36174_);
  nor _46047_ (_37701_, _37690_, _37679_);
  nor _46048_ (_37712_, _37701_, _37657_);
  nor _46049_ (_37723_, _37712_, _37646_);
  and _46050_ (_37734_, _37723_, _37624_);
  not _46051_ (_37745_, _37734_);
  nor _46052_ (_37756_, _37745_, _37591_);
  nor _46053_ (_37767_, _37756_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46054_ (_37778_, _37767_, _36798_);
  nor _46055_ (_37789_, _37778_, _36788_);
  and _46056_ (_37800_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46057_ (_37811_, _36163_, _36842_);
  and _46058_ (_37822_, _37811_, _37431_);
  and _46059_ (_37833_, _37811_, _36020_);
  nor _46060_ (_37844_, _37833_, _37822_);
  and _46061_ (_37855_, _37844_, _36152_);
  nor _46062_ (_37866_, _37855_, _33750_);
  or _46063_ (_37877_, _37866_, _37646_);
  not _46064_ (_37888_, _33750_);
  nor _46065_ (_37899_, _37844_, _37888_);
  nor _46066_ (_37910_, _37899_, _37877_);
  nor _46067_ (_37921_, _37910_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _46068_ (_37932_, _37921_, _37800_);
  and _46069_ (_37943_, _37932_, _41755_);
  and _46070_ (_09542_, _37943_, _37789_);
  and _46071_ (_37964_, _27918_, _24931_);
  and _46072_ (_37975_, _24626_, _24494_);
  and _46073_ (_37986_, _37975_, _25105_);
  and _46074_ (_37997_, _37986_, _24789_);
  and _46075_ (_38008_, _37997_, _29824_);
  and _46076_ (_38019_, _38008_, _37964_);
  not _46077_ (_38030_, _38019_);
  and _46078_ (_38041_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _46079_ (_38052_, _37997_, _24931_);
  and _46080_ (_38063_, _38052_, _24018_);
  and _46081_ (_38074_, _38063_, _29813_);
  and _46082_ (_38085_, _38074_, _27918_);
  not _46083_ (_38096_, _38085_);
  or _46084_ (_38107_, _20924_, _15573_);
  and _46085_ (_38118_, _26217_, _20902_);
  or _46086_ (_38129_, _27676_, _27512_);
  or _46087_ (_38140_, _38129_, _38118_);
  or _46088_ (_38151_, _38140_, _38107_);
  nor _46089_ (_38162_, _38151_, _28805_);
  nor _46090_ (_38173_, _38162_, _16790_);
  not _46091_ (_38184_, _38173_);
  and _46092_ (_38195_, _38184_, _33347_);
  and _46093_ (_38206_, _38195_, _33315_);
  and _46094_ (_38217_, _38206_, _33238_);
  nor _46095_ (_38227_, _38217_, _38096_);
  nor _46096_ (_38238_, _38227_, _38041_);
  and _46097_ (_38249_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _46098_ (_38260_, _38162_, _17826_);
  not _46099_ (_38270_, _38260_);
  and _46100_ (_38281_, _38270_, _32660_);
  and _46101_ (_38292_, _38281_, _32509_);
  nor _46102_ (_38303_, _38292_, _38096_);
  nor _46103_ (_38314_, _38303_, _38249_);
  and _46104_ (_38325_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _46105_ (_38331_, _38162_, _18001_);
  not _46106_ (_38332_, _38331_);
  and _46107_ (_38333_, _38332_, _31834_);
  and _46108_ (_38334_, _38333_, _31692_);
  nor _46109_ (_38335_, _38334_, _38096_);
  nor _46110_ (_38336_, _38335_, _38325_);
  and _46111_ (_38337_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _46112_ (_38338_, _38162_, _18339_);
  not _46113_ (_38339_, _38338_);
  and _46114_ (_38340_, _38339_, _30984_);
  and _46115_ (_38341_, _38340_, _30917_);
  nor _46116_ (_38342_, _38341_, _38096_);
  nor _46117_ (_38343_, _38342_, _38337_);
  and _46118_ (_38344_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _46119_ (_38345_, _38162_, _18861_);
  not _46120_ (_38346_, _38345_);
  and _46121_ (_38347_, _38346_, _30163_);
  and _46122_ (_38348_, _38347_, _30042_);
  nor _46123_ (_38349_, _38348_, _38096_);
  nor _46124_ (_38350_, _38349_, _38344_);
  and _46125_ (_38351_, _38030_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _46126_ (_38352_, _38162_, _18687_);
  not _46127_ (_38353_, _38352_);
  and _46128_ (_38354_, _38353_, _29528_);
  and _46129_ (_38355_, _38354_, _29331_);
  not _46130_ (_38356_, _38355_);
  and _46131_ (_38357_, _38356_, _38085_);
  nor _46132_ (_38358_, _38357_, _38351_);
  nor _46133_ (_38359_, _38019_, _24218_);
  nor _46134_ (_38360_, _38162_, _19231_);
  not _46135_ (_38361_, _38360_);
  and _46136_ (_38362_, _38361_, _28904_);
  and _46137_ (_38363_, _38362_, _28871_);
  and _46138_ (_38364_, _38363_, _28783_);
  not _46139_ (_38365_, _38364_);
  and _46140_ (_38366_, _38365_, _38085_);
  nor _46141_ (_38367_, _38366_, _38359_);
  and _46142_ (_38368_, _38367_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46143_ (_38369_, _38368_, _38358_);
  and _46144_ (_38370_, _38369_, _38350_);
  and _46145_ (_38371_, _38370_, _38343_);
  and _46146_ (_38372_, _38371_, _38336_);
  and _46147_ (_38373_, _38372_, _38314_);
  and _46148_ (_38374_, _38373_, _38238_);
  nor _46149_ (_38375_, _38019_, _24648_);
  nand _46150_ (_38376_, _38375_, _38374_);
  or _46151_ (_38377_, _38375_, _38374_);
  and _46152_ (_38378_, _38377_, _24352_);
  and _46153_ (_38379_, _38378_, _38376_);
  or _46154_ (_38380_, _38019_, _24691_);
  or _46155_ (_38381_, _38380_, _38379_);
  nor _46156_ (_38382_, _38162_, _17630_);
  not _46157_ (_38383_, _38382_);
  and _46158_ (_38384_, _38383_, _27665_);
  and _46159_ (_38385_, _38384_, _27501_);
  and _46160_ (_38386_, _38385_, _27269_);
  nand _46161_ (_38387_, _38386_, _38019_);
  and _46162_ (_38388_, _38387_, _38381_);
  and _46163_ (_09563_, _38388_, _41755_);
  not _46164_ (_38389_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _46165_ (_38390_, _38367_, _38389_);
  nor _46166_ (_38391_, _38367_, _38389_);
  nor _46167_ (_38392_, _38391_, _38390_);
  and _46168_ (_38393_, _38392_, _24352_);
  nor _46169_ (_38394_, _38393_, _24229_);
  nor _46170_ (_38395_, _38394_, _38085_);
  nor _46171_ (_38396_, _38395_, _38366_);
  nand _46172_ (_10690_, _38396_, _41755_);
  nor _46173_ (_38397_, _38368_, _38358_);
  nor _46174_ (_38398_, _38397_, _38369_);
  nor _46175_ (_38399_, _38398_, _23833_);
  nor _46176_ (_38400_, _38399_, _24062_);
  nor _46177_ (_38401_, _38400_, _38085_);
  nor _46178_ (_38402_, _38401_, _38357_);
  nand _46179_ (_10701_, _38402_, _41755_);
  nor _46180_ (_38403_, _38369_, _38350_);
  nor _46181_ (_38404_, _38403_, _38370_);
  nor _46182_ (_38405_, _38404_, _23833_);
  nor _46183_ (_38406_, _38405_, _23887_);
  nor _46184_ (_38407_, _38406_, _38085_);
  nor _46185_ (_38408_, _38407_, _38349_);
  nand _46186_ (_10712_, _38408_, _41755_);
  nor _46187_ (_38409_, _38370_, _38343_);
  nor _46188_ (_38410_, _38409_, _38371_);
  nor _46189_ (_38411_, _38410_, _23833_);
  nor _46190_ (_38412_, _38411_, _24833_);
  nor _46191_ (_38413_, _38412_, _38085_);
  nor _46192_ (_38414_, _38413_, _38342_);
  nor _46193_ (_10723_, _38414_, rst);
  nor _46194_ (_38415_, _38371_, _38336_);
  nor _46195_ (_38416_, _38415_, _38372_);
  nor _46196_ (_38417_, _38416_, _23833_);
  nor _46197_ (_38418_, _38417_, _25039_);
  nor _46198_ (_38419_, _38418_, _38085_);
  nor _46199_ (_38420_, _38419_, _38335_);
  nor _46200_ (_10734_, _38420_, rst);
  nor _46201_ (_38421_, _38372_, _38314_);
  nor _46202_ (_38422_, _38421_, _38373_);
  nor _46203_ (_38423_, _38422_, _23833_);
  nor _46204_ (_38424_, _38423_, _24538_);
  nor _46205_ (_38425_, _38424_, _38085_);
  nor _46206_ (_38426_, _38425_, _38303_);
  nor _46207_ (_10745_, _38426_, rst);
  nor _46208_ (_38427_, _38373_, _38238_);
  nor _46209_ (_38428_, _38427_, _38374_);
  nor _46210_ (_38429_, _38428_, _23833_);
  nor _46211_ (_38430_, _38429_, _24385_);
  nor _46212_ (_38431_, _38430_, _38085_);
  nor _46213_ (_38432_, _38431_, _38227_);
  nor _46214_ (_10756_, _38432_, rst);
  and _46215_ (_38433_, _37964_, _31311_);
  nand _46216_ (_38434_, _38433_, _37997_);
  nor _46217_ (_38435_, _38434_, _27841_);
  and _46218_ (_38436_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15507_);
  and _46219_ (_38437_, _38436_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46220_ (_38438_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _46221_ (_38439_, _38438_, _38437_);
  or _46222_ (_38440_, _38439_, _38435_);
  nor _46223_ (_38441_, _27687_, _17456_);
  nor _46224_ (_38442_, _28291_, _18339_);
  and _46225_ (_38443_, _25910_, _17119_);
  not _46226_ (_38444_, _38443_);
  nor _46227_ (_38445_, _17630_, _16296_);
  and _46228_ (_38446_, _38445_, _27007_);
  and _46229_ (_38447_, _38446_, _26546_);
  and _46230_ (_38448_, _38447_, _26590_);
  and _46231_ (_38449_, _38448_, _26777_);
  nor _46232_ (_38450_, _38449_, _27029_);
  and _46233_ (_38451_, _25910_, _16131_);
  nor _46234_ (_38452_, _38451_, _38450_);
  and _46235_ (_38453_, _38452_, _38444_);
  and _46236_ (_38454_, _27095_, _17630_);
  and _46237_ (_38455_, _16966_, _15967_);
  and _46238_ (_38456_, _17292_, _16296_);
  and _46239_ (_38457_, _38456_, _38455_);
  and _46240_ (_38458_, _38457_, _38454_);
  and _46241_ (_38459_, _17119_, _16131_);
  and _46242_ (_38460_, _38459_, _38458_);
  nor _46243_ (_38461_, _38460_, _25910_);
  not _46244_ (_38462_, _38461_);
  and _46245_ (_38463_, _38462_, _38453_);
  nor _46246_ (_38464_, _25910_, _16471_);
  and _46247_ (_38465_, _25910_, _16471_);
  nor _46248_ (_38466_, _38465_, _38464_);
  and _46249_ (_38467_, _38466_, _38463_);
  and _46250_ (_38468_, _38467_, _27172_);
  nor _46251_ (_38469_, _38467_, _27172_);
  nor _46252_ (_38470_, _38469_, _38468_);
  and _46253_ (_38471_, _38470_, _26941_);
  and _46254_ (_38472_, _25910_, _27172_);
  nor _46255_ (_38473_, _38472_, _28093_);
  nor _46256_ (_38474_, _38473_, _27227_);
  or _46257_ (_38475_, _38474_, _38471_);
  or _46258_ (_38476_, _38475_, _38442_);
  and _46259_ (_38477_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _46260_ (_38478_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _46261_ (_38479_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46262_ (_38480_, _38479_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46263_ (_38481_, _38480_, _38478_);
  nor _46264_ (_38482_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _46265_ (_38483_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46266_ (_38484_, _38483_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46267_ (_38485_, _38484_, _38482_);
  nor _46268_ (_38486_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _46269_ (_38487_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46270_ (_38488_, _38487_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46271_ (_38489_, _38488_, _38486_);
  not _46272_ (_38490_, _38489_);
  nor _46273_ (_38491_, _38490_, _27983_);
  nor _46274_ (_38492_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _46275_ (_38493_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _46276_ (_38494_, _38493_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46277_ (_38495_, _38494_, _38492_);
  and _46278_ (_38496_, _38495_, _38491_);
  nor _46279_ (_38497_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _46280_ (_38498_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _46281_ (_38499_, _38498_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46282_ (_38500_, _38499_, _38497_);
  and _46283_ (_38501_, _38500_, _38496_);
  and _46284_ (_38502_, _38501_, _38485_);
  nor _46285_ (_38503_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _46286_ (_38504_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _46287_ (_38505_, _38504_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46288_ (_38506_, _38505_, _38503_);
  and _46289_ (_38507_, _38506_, _38502_);
  and _46290_ (_38508_, _38507_, _38481_);
  nor _46291_ (_38509_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _46292_ (_38510_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _46293_ (_38511_, _38510_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46294_ (_38512_, _38511_, _38509_);
  and _46295_ (_38513_, _38512_, _38508_);
  nor _46296_ (_38514_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _46297_ (_38515_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _46298_ (_38516_, _38515_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46299_ (_38517_, _38516_, _38514_);
  nor _46300_ (_38518_, _38517_, _38513_);
  and _46301_ (_38519_, _38517_, _38513_);
  or _46302_ (_38520_, _38519_, _38518_);
  nor _46303_ (_38521_, _38520_, _26239_);
  and _46304_ (_38522_, _20616_, _15573_);
  or _46305_ (_38523_, _38522_, _38521_);
  or _46306_ (_38524_, _38523_, _38477_);
  or _46307_ (_38525_, _38524_, _38476_);
  nor _46308_ (_38526_, _38525_, _38441_);
  nand _46309_ (_38527_, _38526_, _38437_);
  and _46310_ (_38528_, _38527_, _41755_);
  and _46311_ (_12702_, _38528_, _38440_);
  and _46312_ (_38529_, _37964_, _30558_);
  and _46313_ (_38530_, _38529_, _37997_);
  nor _46314_ (_38531_, _38530_, _38437_);
  not _46315_ (_38532_, _38531_);
  nand _46316_ (_38533_, _38532_, _27841_);
  or _46317_ (_38534_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _46318_ (_38535_, _38534_, _41755_);
  and _46319_ (_12723_, _38535_, _38533_);
  nor _46320_ (_38536_, _38434_, _29046_);
  and _46321_ (_38537_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _46322_ (_38538_, _38537_, _38437_);
  or _46323_ (_38539_, _38538_, _38536_);
  nor _46324_ (_38540_, _27687_, _16296_);
  nor _46325_ (_38541_, _28291_, _18001_);
  nor _46326_ (_38542_, _27227_, _19231_);
  nor _46327_ (_38543_, _28093_, _27205_);
  not _46328_ (_38544_, _38543_);
  nor _46329_ (_38545_, _38544_, _27117_);
  nor _46330_ (_38546_, _38545_, _26514_);
  and _46331_ (_38547_, _38545_, _26514_);
  nor _46332_ (_38548_, _38547_, _38546_);
  and _46333_ (_38549_, _38548_, _26941_);
  or _46334_ (_38550_, _38549_, _38542_);
  or _46335_ (_38551_, _38550_, _38541_);
  and _46336_ (_38552_, _23201_, _20924_);
  and _46337_ (_38553_, _38490_, _27983_);
  nor _46338_ (_38554_, _38553_, _38491_);
  and _46339_ (_38555_, _38554_, _26228_);
  and _46340_ (_38556_, _20395_, _15573_);
  or _46341_ (_38557_, _38556_, _38555_);
  or _46342_ (_38558_, _38557_, _38552_);
  or _46343_ (_38559_, _38558_, _38551_);
  nor _46344_ (_38560_, _38559_, _38540_);
  nand _46345_ (_38561_, _38560_, _38437_);
  and _46346_ (_38562_, _38561_, _41755_);
  and _46347_ (_13599_, _38562_, _38539_);
  nor _46348_ (_38563_, _38434_, _29714_);
  and _46349_ (_38564_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _46350_ (_38565_, _38564_, _38437_);
  or _46351_ (_38566_, _38565_, _38563_);
  nor _46352_ (_38567_, _27687_, _17292_);
  nor _46353_ (_38568_, _28291_, _17826_);
  and _46354_ (_38569_, _38446_, _25910_);
  and _46355_ (_38570_, _38454_, _16296_);
  and _46356_ (_38571_, _38570_, _27029_);
  nor _46357_ (_38572_, _38571_, _38569_);
  and _46358_ (_38573_, _38572_, _17292_);
  nor _46359_ (_38574_, _38572_, _17292_);
  or _46360_ (_38575_, _38574_, _30864_);
  nor _46361_ (_38576_, _38575_, _38573_);
  nor _46362_ (_38577_, _27227_, _18687_);
  or _46363_ (_38578_, _38577_, _38576_);
  or _46364_ (_38579_, _38578_, _38568_);
  and _46365_ (_38580_, _22233_, _20924_);
  nor _46366_ (_38581_, _38495_, _38491_);
  not _46367_ (_38582_, _38581_);
  nor _46368_ (_38583_, _38496_, _26239_);
  and _46369_ (_38584_, _38583_, _38582_);
  and _46370_ (_38585_, _20427_, _15573_);
  or _46371_ (_38586_, _38585_, _38584_);
  or _46372_ (_38587_, _38586_, _38580_);
  or _46373_ (_38588_, _38587_, _38579_);
  nor _46374_ (_38589_, _38588_, _38567_);
  nand _46375_ (_38590_, _38589_, _38437_);
  and _46376_ (_38591_, _38590_, _41755_);
  and _46377_ (_13608_, _38591_, _38566_);
  nor _46378_ (_38592_, _38434_, _30404_);
  and _46379_ (_38593_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _46380_ (_38594_, _38593_, _38437_);
  or _46381_ (_38595_, _38594_, _38592_);
  nor _46382_ (_38596_, _27687_, _15967_);
  nor _46383_ (_38597_, _28291_, _16790_);
  and _46384_ (_38598_, _38570_, _17292_);
  and _46385_ (_38599_, _38598_, _27029_);
  and _46386_ (_38600_, _38447_, _25910_);
  nor _46387_ (_38601_, _38600_, _38599_);
  and _46388_ (_38602_, _38601_, _15967_);
  nor _46389_ (_38603_, _38601_, _15967_);
  nor _46390_ (_38604_, _38603_, _38602_);
  and _46391_ (_38605_, _38604_, _26941_);
  nor _46392_ (_38606_, _27227_, _18861_);
  or _46393_ (_38607_, _38606_, _38605_);
  or _46394_ (_38608_, _38607_, _38597_);
  and _46395_ (_38609_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _46396_ (_38610_, _38500_, _38496_);
  nor _46397_ (_38611_, _38610_, _38501_);
  and _46398_ (_38612_, _38611_, _26228_);
  and _46399_ (_38613_, _20458_, _15573_);
  or _46400_ (_38614_, _38613_, _38612_);
  or _46401_ (_38615_, _38614_, _38609_);
  or _46402_ (_38616_, _38615_, _38608_);
  nor _46403_ (_38617_, _38616_, _38596_);
  nand _46404_ (_38618_, _38617_, _38437_);
  and _46405_ (_38619_, _38618_, _41755_);
  and _46406_ (_13617_, _38619_, _38595_);
  nor _46407_ (_38620_, _38434_, _31213_);
  and _46408_ (_38621_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _46409_ (_38622_, _38621_, _38437_);
  or _46410_ (_38623_, _38622_, _38620_);
  nor _46411_ (_38624_, _27687_, _16966_);
  nor _46412_ (_38625_, _38448_, _26777_);
  not _46413_ (_38626_, _38625_);
  and _46414_ (_38627_, _38626_, _38450_);
  and _46415_ (_38628_, _38598_, _15967_);
  nor _46416_ (_38629_, _38628_, _16966_);
  nor _46417_ (_38630_, _38629_, _38458_);
  nor _46418_ (_38631_, _38630_, _25910_);
  nor _46419_ (_38632_, _38631_, _38627_);
  nor _46420_ (_38633_, _38632_, _30864_);
  nor _46421_ (_38634_, _27227_, _18339_);
  or _46422_ (_38635_, _38634_, _38633_);
  or _46423_ (_38636_, _38635_, _28302_);
  and _46424_ (_38637_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _46425_ (_38638_, _38501_, _38485_);
  not _46426_ (_38639_, _38638_);
  nor _46427_ (_38640_, _38502_, _26239_);
  and _46428_ (_38641_, _38640_, _38639_);
  and _46429_ (_38642_, _20490_, _15573_);
  or _46430_ (_38643_, _38642_, _38641_);
  or _46431_ (_38644_, _38643_, _38637_);
  or _46432_ (_38645_, _38644_, _38636_);
  nor _46433_ (_38646_, _38645_, _38624_);
  nand _46434_ (_38647_, _38646_, _38437_);
  and _46435_ (_38648_, _38647_, _41755_);
  and _46436_ (_13627_, _38648_, _38623_);
  nor _46437_ (_38649_, _38434_, _31997_);
  and _46438_ (_38650_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _46439_ (_38651_, _38650_, _38437_);
  or _46440_ (_38652_, _38651_, _38649_);
  nor _46441_ (_38653_, _27687_, _16131_);
  nor _46442_ (_38654_, _28291_, _19231_);
  nor _46443_ (_38655_, _38458_, _25910_);
  nor _46444_ (_38656_, _38655_, _38450_);
  nor _46445_ (_38657_, _38656_, _26371_);
  and _46446_ (_38658_, _38656_, _26371_);
  nor _46447_ (_38659_, _38658_, _38657_);
  and _46448_ (_38660_, _38659_, _26941_);
  nor _46449_ (_38661_, _25910_, _18012_);
  or _46450_ (_38662_, _38661_, _27227_);
  nor _46451_ (_38663_, _38662_, _38451_);
  or _46452_ (_38664_, _38663_, _38660_);
  or _46453_ (_38665_, _38664_, _38654_);
  and _46454_ (_38666_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _46455_ (_38667_, _38506_, _38502_);
  not _46456_ (_38668_, _38667_);
  nor _46457_ (_38669_, _38507_, _26239_);
  and _46458_ (_38670_, _38669_, _38668_);
  and _46459_ (_38671_, _20522_, _15573_);
  or _46460_ (_38672_, _38671_, _38670_);
  or _46461_ (_38673_, _38672_, _38666_);
  or _46462_ (_38674_, _38673_, _38665_);
  nor _46463_ (_38675_, _38674_, _38653_);
  nand _46464_ (_38676_, _38675_, _38437_);
  and _46465_ (_38677_, _38676_, _41755_);
  and _46466_ (_13636_, _38677_, _38652_);
  nor _46467_ (_38678_, _38434_, _32814_);
  and _46468_ (_38679_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _46469_ (_38680_, _38679_, _38437_);
  or _46470_ (_38681_, _38680_, _38678_);
  nor _46471_ (_38682_, _27687_, _17119_);
  nor _46472_ (_38683_, _28291_, _18687_);
  and _46473_ (_38684_, _38458_, _16131_);
  nor _46474_ (_38685_, _38684_, _25910_);
  not _46475_ (_38686_, _38685_);
  and _46476_ (_38687_, _38686_, _38452_);
  and _46477_ (_38688_, _38687_, _17119_);
  nor _46478_ (_38689_, _38687_, _17119_);
  or _46479_ (_38690_, _38689_, _38688_);
  and _46480_ (_38691_, _38690_, _26941_);
  nor _46481_ (_38692_, _33151_, _27227_);
  and _46482_ (_38693_, _38692_, _38444_);
  or _46483_ (_38694_, _38693_, _38691_);
  or _46484_ (_38695_, _38694_, _38683_);
  and _46485_ (_38696_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _46486_ (_38697_, _38507_, _38481_);
  not _46487_ (_38698_, _38697_);
  nor _46488_ (_38699_, _38508_, _26239_);
  and _46489_ (_38700_, _38699_, _38698_);
  and _46490_ (_38701_, _20553_, _15573_);
  or _46491_ (_38702_, _38701_, _38700_);
  or _46492_ (_38703_, _38702_, _38696_);
  or _46493_ (_38704_, _38703_, _38695_);
  nor _46494_ (_38705_, _38704_, _38682_);
  nand _46495_ (_38706_, _38705_, _38437_);
  and _46496_ (_38707_, _38706_, _41755_);
  and _46497_ (_13646_, _38707_, _38681_);
  nor _46498_ (_38708_, _38434_, _33533_);
  and _46499_ (_38709_, _38434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _46500_ (_38710_, _38709_, _38437_);
  or _46501_ (_38711_, _38710_, _38708_);
  nor _46502_ (_38712_, _27687_, _16471_);
  nor _46503_ (_38713_, _28291_, _18861_);
  nor _46504_ (_38714_, _38463_, _26327_);
  not _46505_ (_38715_, _38714_);
  and _46506_ (_38716_, _38463_, _26327_);
  nor _46507_ (_38717_, _38716_, _30864_);
  and _46508_ (_38718_, _38717_, _38715_);
  nor _46509_ (_38719_, _25910_, _16801_);
  or _46510_ (_38720_, _38719_, _27227_);
  nor _46511_ (_38721_, _38720_, _38465_);
  or _46512_ (_38722_, _38721_, _38718_);
  or _46513_ (_38723_, _38722_, _38713_);
  and _46514_ (_38724_, _20924_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _46515_ (_38725_, _38512_, _38508_);
  nor _46516_ (_38726_, _38725_, _38513_);
  and _46517_ (_38727_, _38726_, _26228_);
  and _46518_ (_38728_, _20585_, _15573_);
  or _46519_ (_38729_, _38728_, _38727_);
  or _46520_ (_38730_, _38729_, _38724_);
  or _46521_ (_38731_, _38730_, _38723_);
  nor _46522_ (_38732_, _38731_, _38712_);
  nand _46523_ (_38733_, _38732_, _38437_);
  and _46524_ (_38734_, _38733_, _41755_);
  and _46525_ (_13656_, _38734_, _38711_);
  nand _46526_ (_38735_, _38532_, _29046_);
  or _46527_ (_38736_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _46528_ (_38737_, _38736_, _41755_);
  and _46529_ (_13665_, _38737_, _38735_);
  nand _46530_ (_38738_, _38532_, _29714_);
  or _46531_ (_38739_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _46532_ (_38740_, _38739_, _41755_);
  and _46533_ (_13675_, _38740_, _38738_);
  nand _46534_ (_38741_, _38532_, _30404_);
  or _46535_ (_38742_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _46536_ (_38743_, _38742_, _41755_);
  and _46537_ (_13684_, _38743_, _38741_);
  nand _46538_ (_38744_, _38532_, _31213_);
  or _46539_ (_38745_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _46540_ (_38746_, _38745_, _41755_);
  and _46541_ (_13694_, _38746_, _38744_);
  nand _46542_ (_38747_, _38532_, _31997_);
  or _46543_ (_38748_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _46544_ (_38749_, _38748_, _41755_);
  and _46545_ (_13704_, _38749_, _38747_);
  nand _46546_ (_38750_, _38532_, _32814_);
  or _46547_ (_38751_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _46548_ (_38752_, _38751_, _41755_);
  and _46549_ (_13713_, _38752_, _38750_);
  nand _46550_ (_38753_, _38532_, _33533_);
  or _46551_ (_38754_, _38532_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _46552_ (_38755_, _38754_, _41755_);
  and _46553_ (_13722_, _38755_, _38753_);
  not _46554_ (_38756_, _24494_);
  and _46555_ (_38757_, _25116_, _24626_);
  and _46556_ (_38758_, _38757_, _38756_);
  and _46557_ (_38760_, _28576_, _24789_);
  and _46558_ (_38763_, _38760_, _38758_);
  not _46559_ (_38764_, _28543_);
  nor _46560_ (_38765_, _38764_, _28510_);
  not _46561_ (_38766_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _46562_ (_38767_, _28543_, _38766_);
  or _46563_ (_38768_, _38767_, _38765_);
  and _46564_ (_38769_, _38768_, _38763_);
  and _46565_ (_38770_, _27918_, _24287_);
  nor _46566_ (_38771_, _24494_, _24778_);
  and _46567_ (_38772_, _38757_, _38771_);
  and _46568_ (_38773_, _38772_, _38770_);
  nor _46569_ (_38782_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _46570_ (_38788_, _38782_);
  nand _46571_ (_38794_, _38788_, _28510_);
  and _46572_ (_38798_, _38772_, _28576_);
  and _46573_ (_38799_, _38782_, _38766_);
  nor _46574_ (_38800_, _38799_, _38798_);
  and _46575_ (_38801_, _38800_, _38794_);
  or _46576_ (_38802_, _38801_, _38773_);
  or _46577_ (_38803_, _38802_, _38769_);
  nand _46578_ (_38804_, _38773_, _38386_);
  and _46579_ (_38805_, _38804_, _38803_);
  and _46580_ (_16559_, _38805_, _41755_);
  not _46581_ (_38806_, _38773_);
  nor _46582_ (_38807_, _38806_, _38355_);
  and _46583_ (_38808_, _38763_, _29824_);
  or _46584_ (_38809_, _38808_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _46585_ (_38810_, _38809_, _38806_);
  nand _46586_ (_38811_, _38808_, _28510_);
  and _46587_ (_38812_, _38811_, _38810_);
  or _46588_ (_38813_, _38812_, _38807_);
  and _46589_ (_21487_, _38813_, _41755_);
  nor _46590_ (_38814_, _38806_, _38348_);
  and _46591_ (_38815_, _30569_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _46592_ (_38816_, _38815_, _30580_);
  and _46593_ (_38817_, _38816_, _38798_);
  and _46594_ (_38818_, _28016_, _26876_);
  not _46595_ (_38819_, _26876_);
  and _46596_ (_38820_, _28027_, _38819_);
  or _46597_ (_38822_, _38820_, _38818_);
  and _46598_ (_38824_, _38822_, _26305_);
  not _46599_ (_38825_, _26141_);
  nand _46600_ (_38826_, _26130_, _38825_);
  or _46601_ (_38827_, _26152_, _26130_);
  and _46602_ (_38828_, _26228_, _38827_);
  and _46603_ (_38829_, _38828_, _38826_);
  and _46604_ (_38830_, _38459_, _22135_);
  and _46605_ (_38831_, _38457_, _20924_);
  nand _46606_ (_38832_, _38831_, _38830_);
  nand _46607_ (_38833_, _38832_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46608_ (_38834_, _38833_, _38829_);
  or _46609_ (_38835_, _38834_, _38824_);
  or _46610_ (_38836_, _38835_, _33020_);
  or _46611_ (_38837_, _20680_, _20648_);
  or _46612_ (_38838_, _38837_, _20711_);
  or _46613_ (_38839_, _38838_, _20754_);
  or _46614_ (_38840_, _38839_, _20785_);
  or _46615_ (_38841_, _38840_, _20828_);
  and _46616_ (_38842_, _38841_, _15573_);
  or _46617_ (_38843_, _38842_, _38836_);
  or _46618_ (_38844_, _38843_, _25181_);
  nor _46619_ (_38845_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _46620_ (_38846_, _38845_, _38798_);
  and _46621_ (_38847_, _38846_, _38844_);
  or _46622_ (_38848_, _38847_, _38817_);
  and _46623_ (_38849_, _38848_, _38806_);
  or _46624_ (_38850_, _38849_, _38814_);
  and _46625_ (_21499_, _38850_, _41755_);
  not _46626_ (_38851_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand _46627_ (_38852_, _38798_, _31311_);
  nand _46628_ (_38853_, _38852_, _38851_);
  and _46629_ (_38854_, _38853_, _38806_);
  or _46630_ (_38855_, _38852_, _29134_);
  and _46631_ (_38856_, _38855_, _38854_);
  nor _46632_ (_38857_, _38806_, _38341_);
  or _46633_ (_38858_, _38857_, _38856_);
  and _46634_ (_21511_, _38858_, _41755_);
  not _46635_ (_38860_, _38798_);
  or _46636_ (_38863_, _38860_, _32117_);
  and _46637_ (_38869_, _38863_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _46638_ (_38874_, _32106_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _46639_ (_38881_, _38874_, _32150_);
  and _46640_ (_38888_, _38881_, _38798_);
  or _46641_ (_38898_, _38888_, _38869_);
  and _46642_ (_38899_, _38898_, _38806_);
  nor _46643_ (_38900_, _38806_, _38334_);
  or _46644_ (_38901_, _38900_, _38899_);
  and _46645_ (_21523_, _38901_, _41755_);
  nor _46646_ (_38902_, _38806_, _38292_);
  and _46647_ (_38903_, _38763_, _32901_);
  or _46648_ (_38904_, _38903_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _46649_ (_38905_, _38904_, _38806_);
  nand _46650_ (_38906_, _38903_, _28510_);
  and _46651_ (_38907_, _38906_, _38905_);
  or _46652_ (_38908_, _38907_, _38902_);
  and _46653_ (_21535_, _38908_, _41755_);
  nor _46654_ (_38909_, _38806_, _38217_);
  not _46655_ (_38910_, _33631_);
  nor _46656_ (_38911_, _38910_, _28510_);
  or _46657_ (_38912_, _33631_, _30995_);
  nand _46658_ (_38913_, _38912_, _38798_);
  or _46659_ (_38914_, _38913_, _38911_);
  and _46660_ (_38915_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _46661_ (_38916_, _26228_, _26053_);
  and _46662_ (_38917_, _26832_, _26305_);
  or _46663_ (_38918_, _38917_, _38916_);
  and _46664_ (_38919_, _38918_, _38915_);
  nand _46665_ (_38920_, _38915_, _27687_);
  and _46666_ (_38921_, _38920_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _46667_ (_38922_, _38921_, _38798_);
  or _46668_ (_38923_, _38922_, _38919_);
  and _46669_ (_38924_, _38923_, _38806_);
  and _46670_ (_38925_, _38924_, _38914_);
  or _46671_ (_38926_, _38925_, _38909_);
  and _46672_ (_21547_, _38926_, _41755_);
  not _46673_ (_38927_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46674_ (_38928_, _38436_, _38927_);
  and _46675_ (_38929_, _38928_, _38526_);
  nor _46676_ (_38930_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46677_ (_38931_, _38930_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46678_ (_38932_, _24287_, _24931_);
  not _46679_ (_38936_, _24626_);
  and _46680_ (_38947_, _25105_, _38936_);
  and _46681_ (_38950_, _38947_, _27918_);
  and _46682_ (_38951_, _38950_, _38932_);
  and _46683_ (_38952_, _38951_, _38771_);
  nor _46684_ (_38961_, _38952_, _38931_);
  nor _46685_ (_38969_, _38961_, _27841_);
  and _46686_ (_38970_, _25105_, _24931_);
  and _46687_ (_38971_, _38970_, _24637_);
  and _46688_ (_38972_, _38971_, _38760_);
  and _46689_ (_38973_, _38972_, _28543_);
  and _46690_ (_38974_, _38973_, _28510_);
  nor _46691_ (_38975_, _38973_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _46692_ (_38976_, _38928_);
  and _46693_ (_38977_, _38961_, _38976_);
  not _46694_ (_38978_, _38977_);
  nor _46695_ (_38979_, _38978_, _38975_);
  not _46696_ (_38980_, _38979_);
  nor _46697_ (_38981_, _38980_, _38974_);
  nor _46698_ (_38982_, _38981_, _38928_);
  not _46699_ (_38983_, _38982_);
  nor _46700_ (_38984_, _38983_, _38969_);
  nor _46701_ (_38985_, _38984_, _38929_);
  and _46702_ (_22320_, _38985_, _41755_);
  nor _46703_ (_38986_, _38961_, _29046_);
  and _46704_ (_38987_, _38972_, _24287_);
  and _46705_ (_38988_, _38987_, _28510_);
  nor _46706_ (_38989_, _38987_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _46707_ (_38990_, _38989_, _38978_);
  not _46708_ (_38991_, _38990_);
  nor _46709_ (_38992_, _38991_, _38988_);
  or _46710_ (_38993_, _38992_, _38986_);
  and _46711_ (_38994_, _38993_, _38976_);
  nor _46712_ (_38995_, _38976_, _38560_);
  or _46713_ (_38996_, _38995_, _38994_);
  and _46714_ (_24171_, _38996_, _41755_);
  and _46715_ (_38997_, _38928_, _38589_);
  nor _46716_ (_38998_, _38961_, _29714_);
  and _46717_ (_38999_, _38972_, _29824_);
  and _46718_ (_39000_, _38999_, _28510_);
  nor _46719_ (_39001_, _38999_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _46720_ (_39002_, _39001_, _38978_);
  not _46721_ (_39003_, _39002_);
  nor _46722_ (_39004_, _39003_, _39000_);
  nor _46723_ (_39005_, _39004_, _38928_);
  not _46724_ (_39006_, _39005_);
  nor _46725_ (_39007_, _39006_, _38998_);
  nor _46726_ (_39008_, _39007_, _38997_);
  and _46727_ (_24183_, _39008_, _41755_);
  nor _46728_ (_39009_, _38961_, _30404_);
  and _46729_ (_39010_, _38972_, _30558_);
  and _46730_ (_39011_, _39010_, _28510_);
  nor _46731_ (_39012_, _39010_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _46732_ (_39013_, _39012_, _38978_);
  not _46733_ (_39014_, _39013_);
  nor _46734_ (_39015_, _39014_, _39011_);
  or _46735_ (_39016_, _39015_, _39009_);
  and _46736_ (_39017_, _39016_, _38976_);
  nor _46737_ (_39018_, _38976_, _38617_);
  or _46738_ (_39019_, _39018_, _39017_);
  and _46739_ (_24195_, _39019_, _41755_);
  nor _46740_ (_39020_, _38961_, _31213_);
  not _46741_ (_39021_, _38972_);
  and _46742_ (_39022_, _38977_, _39021_);
  and _46743_ (_39023_, _39022_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _46744_ (_39024_, _31322_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _46745_ (_39025_, _39024_, _31333_);
  and _46746_ (_39026_, _38972_, _38976_);
  not _46747_ (_39027_, _39026_);
  nor _46748_ (_39028_, _39027_, _39025_);
  and _46749_ (_39029_, _39028_, _38977_);
  nor _46750_ (_39030_, _39029_, _39023_);
  and _46751_ (_39031_, _39030_, _38976_);
  not _46752_ (_39032_, _39031_);
  nor _46753_ (_39033_, _39032_, _39020_);
  and _46754_ (_39034_, _38928_, _38646_);
  or _46755_ (_39035_, _39034_, _39033_);
  nor _46756_ (_24207_, _39035_, rst);
  nor _46757_ (_39036_, _38961_, _31997_);
  and _46758_ (_39037_, _38972_, _32096_);
  and _46759_ (_39038_, _39037_, _28510_);
  nor _46760_ (_39039_, _39037_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _46761_ (_39040_, _39039_, _38978_);
  not _46762_ (_39041_, _39040_);
  nor _46763_ (_39042_, _39041_, _39038_);
  or _46764_ (_39043_, _39042_, _39036_);
  and _46765_ (_39044_, _39043_, _38976_);
  nor _46766_ (_39045_, _38976_, _38675_);
  or _46767_ (_39046_, _39045_, _39044_);
  and _46768_ (_24219_, _39046_, _41755_);
  nor _46769_ (_39047_, _38961_, _32814_);
  and _46770_ (_39048_, _38972_, _32901_);
  and _46771_ (_39049_, _39048_, _28510_);
  nor _46772_ (_39050_, _39048_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _46773_ (_39051_, _39050_, _38978_);
  not _46774_ (_39052_, _39051_);
  nor _46775_ (_39053_, _39052_, _39049_);
  or _46776_ (_39054_, _39053_, _39047_);
  and _46777_ (_39055_, _39054_, _38976_);
  nor _46778_ (_39056_, _38976_, _38705_);
  or _46779_ (_39057_, _39056_, _39055_);
  and _46780_ (_24230_, _39057_, _41755_);
  nor _46781_ (_39058_, _38961_, _33533_);
  and _46782_ (_39059_, _38972_, _33631_);
  and _46783_ (_39060_, _39059_, _28510_);
  nor _46784_ (_39061_, _39059_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _46785_ (_39062_, _39061_, _38978_);
  not _46786_ (_39063_, _39062_);
  nor _46787_ (_39064_, _39063_, _39060_);
  or _46788_ (_39065_, _39064_, _39058_);
  and _46789_ (_39066_, _39065_, _38976_);
  nor _46790_ (_39067_, _38976_, _38732_);
  or _46791_ (_39068_, _39067_, _39066_);
  and _46792_ (_24242_, _39068_, _41755_);
  and _46793_ (_39069_, _38052_, _28543_);
  nand _46794_ (_39070_, _39069_, _28510_);
  or _46795_ (_39071_, _39069_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46796_ (_39072_, _39071_, _28576_);
  and _46797_ (_39073_, _39072_, _39070_);
  and _46798_ (_39074_, _37997_, _38932_);
  nand _46799_ (_39075_, _39074_, _38386_);
  or _46800_ (_39076_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46801_ (_39077_, _39076_, _27918_);
  and _46802_ (_39078_, _39077_, _39075_);
  and _46803_ (_39079_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _46804_ (_39080_, _39079_, rst);
  or _46805_ (_39081_, _39080_, _39078_);
  or _46806_ (_35499_, _39081_, _39073_);
  nor _46807_ (_39082_, _38756_, _24778_);
  and _46808_ (_39083_, _38757_, _39082_);
  and _46809_ (_39084_, _39083_, _28543_);
  nand _46810_ (_39085_, _39084_, _28510_);
  or _46811_ (_39086_, _39084_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46812_ (_39087_, _39086_, _28576_);
  and _46813_ (_39088_, _39087_, _39085_);
  and _46814_ (_39089_, _39083_, _24287_);
  not _46815_ (_39090_, _39089_);
  nor _46816_ (_39091_, _39090_, _38386_);
  and _46817_ (_39092_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _46818_ (_39093_, _39092_, _39091_);
  and _46819_ (_39094_, _39093_, _27918_);
  and _46820_ (_39095_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _46821_ (_39096_, _39095_, rst);
  or _46822_ (_39097_, _39096_, _39094_);
  or _46823_ (_35522_, _39097_, _39088_);
  and _46824_ (_39098_, _38936_, _24494_);
  and _46825_ (_39099_, _39098_, _38970_);
  and _46826_ (_39100_, _39099_, _24789_);
  and _46827_ (_39101_, _39100_, _28543_);
  nand _46828_ (_39102_, _39101_, _28510_);
  or _46829_ (_39103_, _39101_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _46830_ (_39104_, _39103_, _28576_);
  and _46831_ (_39105_, _39104_, _39102_);
  and _46832_ (_39106_, _38947_, _39082_);
  and _46833_ (_39107_, _39106_, _38932_);
  not _46834_ (_39108_, _39107_);
  nor _46835_ (_39109_, _39108_, _38386_);
  and _46836_ (_39110_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46837_ (_39111_, _39110_, _39109_);
  and _46838_ (_39112_, _39111_, _27918_);
  and _46839_ (_39113_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46840_ (_39114_, _39113_, rst);
  or _46841_ (_39115_, _39114_, _39112_);
  or _46842_ (_35545_, _39115_, _39105_);
  and _46843_ (_39116_, _39098_, _25127_);
  and _46844_ (_39117_, _39116_, _28543_);
  nand _46845_ (_39118_, _39117_, _28510_);
  or _46846_ (_39119_, _39117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _46847_ (_39120_, _39119_, _28576_);
  and _46848_ (_39121_, _39120_, _39118_);
  nor _46849_ (_39122_, _25105_, _24626_);
  and _46850_ (_39123_, _39082_, _39122_);
  and _46851_ (_39124_, _39123_, _38932_);
  not _46852_ (_39125_, _39124_);
  nor _46853_ (_39126_, _39125_, _38386_);
  and _46854_ (_39127_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46855_ (_39128_, _39127_, _39126_);
  and _46856_ (_39129_, _39128_, _27918_);
  and _46857_ (_39130_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46858_ (_39131_, _39130_, rst);
  or _46859_ (_39132_, _39131_, _39129_);
  or _46860_ (_35568_, _39132_, _39121_);
  not _46861_ (_39133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _46862_ (_39134_, _39074_, _39133_);
  nand _46863_ (_39135_, _38052_, _24287_);
  nor _46864_ (_39136_, _39135_, _28510_);
  or _46865_ (_39137_, _39136_, _39134_);
  and _46866_ (_39138_, _39137_, _28576_);
  and _46867_ (_39139_, _39074_, _38365_);
  or _46868_ (_39140_, _39139_, _39134_);
  and _46869_ (_39141_, _39140_, _27918_);
  nor _46870_ (_39142_, _27896_, _39133_);
  or _46871_ (_39143_, _39142_, rst);
  or _46872_ (_39144_, _39143_, _39141_);
  or _46873_ (_41155_, _39144_, _39138_);
  or _46874_ (_39161_, _38074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46875_ (_39172_, _39161_, _28576_);
  nand _46876_ (_39182_, _38074_, _28510_);
  and _46877_ (_39188_, _39182_, _39172_);
  nand _46878_ (_39198_, _39074_, _38355_);
  or _46879_ (_39209_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46880_ (_39220_, _39209_, _27918_);
  and _46881_ (_39231_, _39220_, _39198_);
  and _46882_ (_39242_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _46883_ (_39253_, _39242_, rst);
  or _46884_ (_39264_, _39253_, _39231_);
  or _46885_ (_41157_, _39264_, _39188_);
  not _46886_ (_39285_, _31344_);
  nand _46887_ (_39296_, _38052_, _39285_);
  and _46888_ (_39307_, _39296_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46889_ (_39318_, _30590_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46890_ (_39329_, _39318_, _30580_);
  and _46891_ (_39340_, _39329_, _38052_);
  or _46892_ (_39351_, _39340_, _39307_);
  and _46893_ (_39357_, _39351_, _28576_);
  nand _46894_ (_39358_, _39074_, _38348_);
  or _46895_ (_39359_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46896_ (_39360_, _39359_, _27918_);
  and _46897_ (_39361_, _39360_, _39358_);
  and _46898_ (_39362_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46899_ (_39363_, _39362_, rst);
  or _46900_ (_39364_, _39363_, _39361_);
  or _46901_ (_41158_, _39364_, _39357_);
  not _46902_ (_39365_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor _46903_ (_39366_, _38063_, _39365_);
  nor _46904_ (_39367_, _31344_, _39365_);
  or _46905_ (_39368_, _39367_, _31333_);
  and _46906_ (_39369_, _39368_, _38052_);
  or _46907_ (_39370_, _39369_, _39366_);
  and _46908_ (_39371_, _39370_, _28576_);
  nand _46909_ (_39372_, _39074_, _38341_);
  or _46910_ (_39373_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46911_ (_39374_, _39373_, _27918_);
  and _46912_ (_39375_, _39374_, _39372_);
  nor _46913_ (_39376_, _27896_, _39365_);
  or _46914_ (_39377_, _39376_, rst);
  or _46915_ (_39378_, _39377_, _39375_);
  or _46916_ (_41160_, _39378_, _39371_);
  not _46917_ (_39379_, _38052_);
  or _46918_ (_39380_, _39379_, _32117_);
  and _46919_ (_39381_, _39380_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46920_ (_39382_, _32106_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46921_ (_39383_, _39382_, _32150_);
  and _46922_ (_39384_, _39383_, _38052_);
  or _46923_ (_39385_, _39384_, _39381_);
  and _46924_ (_39386_, _39385_, _28576_);
  nand _46925_ (_39387_, _39074_, _38334_);
  or _46926_ (_39388_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46927_ (_39389_, _39388_, _27918_);
  and _46928_ (_39390_, _39389_, _39387_);
  and _46929_ (_39391_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46930_ (_39392_, _39391_, rst);
  or _46931_ (_39393_, _39392_, _39390_);
  or _46932_ (_41162_, _39393_, _39386_);
  and _46933_ (_39394_, _38052_, _32901_);
  nand _46934_ (_39395_, _39394_, _28510_);
  or _46935_ (_39396_, _39394_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46936_ (_39397_, _39396_, _28576_);
  and _46937_ (_39398_, _39397_, _39395_);
  nand _46938_ (_39399_, _39074_, _38292_);
  or _46939_ (_39400_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46940_ (_39401_, _39400_, _27918_);
  and _46941_ (_39402_, _39401_, _39399_);
  and _46942_ (_39403_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _46943_ (_39404_, _39403_, rst);
  or _46944_ (_39405_, _39404_, _39402_);
  or _46945_ (_41164_, _39405_, _39398_);
  and _46946_ (_39406_, _38052_, _33631_);
  nand _46947_ (_39407_, _39406_, _28510_);
  or _46948_ (_39408_, _39406_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _46949_ (_39409_, _39408_, _28576_);
  and _46950_ (_39410_, _39409_, _39407_);
  nand _46951_ (_39411_, _39074_, _38217_);
  or _46952_ (_39412_, _39074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _46953_ (_39413_, _39412_, _27918_);
  and _46954_ (_39414_, _39413_, _39411_);
  and _46955_ (_39415_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _46956_ (_39416_, _39415_, rst);
  or _46957_ (_39417_, _39416_, _39414_);
  or _46958_ (_41165_, _39417_, _39410_);
  nand _46959_ (_39418_, _39089_, _28510_);
  or _46960_ (_39419_, _39089_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _46961_ (_39420_, _39419_, _28576_);
  and _46962_ (_39421_, _39420_, _39418_);
  and _46963_ (_39422_, _39089_, _38365_);
  and _46964_ (_39423_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _46965_ (_39424_, _39423_, _39422_);
  and _46966_ (_39425_, _39424_, _27918_);
  and _46967_ (_39426_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _46968_ (_39427_, _39426_, rst);
  or _46969_ (_39428_, _39427_, _39425_);
  or _46970_ (_41167_, _39428_, _39421_);
  and _46971_ (_39429_, _39083_, _29824_);
  nand _46972_ (_39430_, _39429_, _28510_);
  or _46973_ (_39431_, _39429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _46974_ (_39432_, _39431_, _28576_);
  and _46975_ (_39433_, _39432_, _39430_);
  nor _46976_ (_39434_, _39090_, _38355_);
  and _46977_ (_39435_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _46978_ (_39436_, _39435_, _39434_);
  and _46979_ (_39437_, _39436_, _27918_);
  and _46980_ (_39438_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _46981_ (_39439_, _39438_, rst);
  or _46982_ (_39440_, _39439_, _39437_);
  or _46983_ (_41169_, _39440_, _39433_);
  and _46984_ (_39441_, _39083_, _30558_);
  nand _46985_ (_39442_, _39441_, _28510_);
  or _46986_ (_39443_, _39441_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _46987_ (_39444_, _39443_, _28576_);
  and _46988_ (_39445_, _39444_, _39442_);
  nor _46989_ (_39446_, _39090_, _38348_);
  and _46990_ (_39447_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _46991_ (_39448_, _39447_, _39446_);
  and _46992_ (_39449_, _39448_, _27918_);
  and _46993_ (_39450_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _46994_ (_39451_, _39450_, rst);
  or _46995_ (_39452_, _39451_, _39449_);
  or _46996_ (_41171_, _39452_, _39445_);
  and _46997_ (_39453_, _39083_, _31311_);
  nand _46998_ (_39454_, _39453_, _28510_);
  or _46999_ (_39455_, _39453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _47000_ (_39456_, _39455_, _28576_);
  and _47001_ (_39457_, _39456_, _39454_);
  nor _47002_ (_39458_, _39090_, _38341_);
  and _47003_ (_39459_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _47004_ (_39460_, _39459_, _39458_);
  and _47005_ (_39461_, _39460_, _27918_);
  and _47006_ (_39462_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _47007_ (_39463_, _39462_, rst);
  or _47008_ (_39464_, _39463_, _39461_);
  or _47009_ (_41172_, _39464_, _39457_);
  and _47010_ (_39465_, _39083_, _32096_);
  nand _47011_ (_39466_, _39465_, _28510_);
  or _47012_ (_39467_, _39465_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _47013_ (_39468_, _39467_, _28576_);
  and _47014_ (_39469_, _39468_, _39466_);
  nor _47015_ (_39470_, _39090_, _38334_);
  and _47016_ (_39471_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _47017_ (_39472_, _39471_, _39470_);
  and _47018_ (_39473_, _39472_, _27918_);
  and _47019_ (_39474_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _47020_ (_39475_, _39474_, rst);
  or _47021_ (_39476_, _39475_, _39473_);
  or _47022_ (_41174_, _39476_, _39469_);
  and _47023_ (_39477_, _39083_, _32901_);
  nand _47024_ (_39478_, _39477_, _28510_);
  or _47025_ (_39479_, _39477_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _47026_ (_39480_, _39479_, _28576_);
  and _47027_ (_39481_, _39480_, _39478_);
  nor _47028_ (_39482_, _39090_, _38292_);
  and _47029_ (_39483_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _47030_ (_39484_, _39483_, _39482_);
  and _47031_ (_39485_, _39484_, _27918_);
  and _47032_ (_39486_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _47033_ (_39487_, _39486_, rst);
  or _47034_ (_39488_, _39487_, _39485_);
  or _47035_ (_41176_, _39488_, _39481_);
  and _47036_ (_39489_, _39083_, _33631_);
  nand _47037_ (_39490_, _39489_, _28510_);
  or _47038_ (_39491_, _39489_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _47039_ (_39492_, _39491_, _28576_);
  and _47040_ (_39493_, _39492_, _39490_);
  nor _47041_ (_39494_, _39090_, _38217_);
  and _47042_ (_39495_, _39090_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _47043_ (_39496_, _39495_, _39494_);
  and _47044_ (_39497_, _39496_, _27918_);
  and _47045_ (_39498_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _47046_ (_39499_, _39498_, rst);
  or _47047_ (_39500_, _39499_, _39497_);
  or _47048_ (_41178_, _39500_, _39493_);
  nand _47049_ (_39501_, _39107_, _28510_);
  or _47050_ (_39502_, _39107_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _47051_ (_39503_, _39502_, _28576_);
  and _47052_ (_39504_, _39503_, _39501_);
  and _47053_ (_39505_, _39107_, _38365_);
  and _47054_ (_39506_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _47055_ (_39507_, _39506_, _39505_);
  and _47056_ (_39508_, _39507_, _27918_);
  and _47057_ (_39509_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _47058_ (_39510_, _39509_, rst);
  or _47059_ (_39511_, _39510_, _39508_);
  or _47060_ (_41179_, _39511_, _39504_);
  and _47061_ (_39512_, _39100_, _29824_);
  nand _47062_ (_39513_, _39512_, _28510_);
  or _47063_ (_39514_, _39512_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _47064_ (_39515_, _39514_, _28576_);
  and _47065_ (_39516_, _39515_, _39513_);
  nor _47066_ (_39517_, _39108_, _38355_);
  and _47067_ (_39518_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _47068_ (_39519_, _39518_, _39517_);
  and _47069_ (_39520_, _39519_, _27918_);
  and _47070_ (_39521_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _47071_ (_39522_, _39521_, rst);
  or _47072_ (_39523_, _39522_, _39520_);
  or _47073_ (_41181_, _39523_, _39516_);
  and _47074_ (_39524_, _39100_, _30558_);
  nand _47075_ (_39525_, _39524_, _28510_);
  or _47076_ (_39526_, _39524_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _47077_ (_39527_, _39526_, _28576_);
  and _47078_ (_39528_, _39527_, _39525_);
  nor _47079_ (_39529_, _39108_, _38348_);
  and _47080_ (_39530_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _47081_ (_39531_, _39530_, _39529_);
  and _47082_ (_39532_, _39531_, _27918_);
  and _47083_ (_39533_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _47084_ (_39534_, _39533_, rst);
  or _47085_ (_39535_, _39534_, _39532_);
  or _47086_ (_41183_, _39535_, _39528_);
  and _47087_ (_39536_, _39100_, _31311_);
  nand _47088_ (_39537_, _39536_, _28510_);
  or _47089_ (_39538_, _39536_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _47090_ (_39539_, _39538_, _28576_);
  and _47091_ (_39540_, _39539_, _39537_);
  nor _47092_ (_39541_, _39108_, _38341_);
  and _47093_ (_39542_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _47094_ (_39543_, _39542_, _39541_);
  and _47095_ (_39544_, _39543_, _27918_);
  and _47096_ (_39545_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _47097_ (_39546_, _39545_, rst);
  or _47098_ (_39547_, _39546_, _39544_);
  or _47099_ (_41185_, _39547_, _39540_);
  and _47100_ (_39548_, _39100_, _32096_);
  nand _47101_ (_39549_, _39548_, _28510_);
  or _47102_ (_39550_, _39548_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _47103_ (_39551_, _39550_, _28576_);
  and _47104_ (_39552_, _39551_, _39549_);
  nor _47105_ (_39553_, _39108_, _38334_);
  and _47106_ (_39554_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _47107_ (_39555_, _39554_, _39553_);
  and _47108_ (_39556_, _39555_, _27918_);
  and _47109_ (_39557_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _47110_ (_39558_, _39557_, rst);
  or _47111_ (_39559_, _39558_, _39556_);
  or _47112_ (_41186_, _39559_, _39552_);
  and _47113_ (_39560_, _39100_, _32901_);
  nand _47114_ (_39561_, _39560_, _28510_);
  or _47115_ (_39562_, _39560_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _47116_ (_39564_, _39562_, _28576_);
  and _47117_ (_39565_, _39564_, _39561_);
  nor _47118_ (_39566_, _39108_, _38292_);
  and _47119_ (_39567_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _47120_ (_39568_, _39567_, _39566_);
  and _47121_ (_39569_, _39568_, _27918_);
  and _47122_ (_39570_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _47123_ (_39571_, _39570_, rst);
  or _47124_ (_39572_, _39571_, _39569_);
  or _47125_ (_41188_, _39572_, _39565_);
  and _47126_ (_39573_, _39100_, _33631_);
  nand _47127_ (_39574_, _39573_, _28510_);
  or _47128_ (_39575_, _39573_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _47129_ (_39576_, _39575_, _28576_);
  and _47130_ (_39577_, _39576_, _39574_);
  nor _47131_ (_39578_, _39108_, _38217_);
  and _47132_ (_39579_, _39108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _47133_ (_39580_, _39579_, _39578_);
  and _47134_ (_39581_, _39580_, _27918_);
  and _47135_ (_39582_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _47136_ (_39583_, _39582_, rst);
  or _47137_ (_39584_, _39583_, _39581_);
  or _47138_ (_41190_, _39584_, _39577_);
  and _47139_ (_39585_, _39116_, _24287_);
  nand _47140_ (_39586_, _39585_, _28510_);
  or _47141_ (_39587_, _39585_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _47142_ (_39588_, _39587_, _28576_);
  and _47143_ (_39589_, _39588_, _39586_);
  and _47144_ (_39590_, _39124_, _38365_);
  and _47145_ (_39591_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _47146_ (_39592_, _39591_, _39590_);
  and _47147_ (_39593_, _39592_, _27918_);
  and _47148_ (_39598_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _47149_ (_39599_, _39598_, rst);
  or _47150_ (_39600_, _39599_, _39593_);
  or _47151_ (_41192_, _39600_, _39589_);
  and _47152_ (_39601_, _39116_, _29824_);
  nand _47153_ (_39602_, _39601_, _28510_);
  or _47154_ (_39603_, _39601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _47155_ (_39604_, _39603_, _28576_);
  and _47156_ (_39605_, _39604_, _39602_);
  nor _47157_ (_39606_, _39125_, _38355_);
  and _47158_ (_39607_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47159_ (_39608_, _39607_, _39606_);
  and _47160_ (_39609_, _39608_, _27918_);
  and _47161_ (_39610_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47162_ (_39611_, _39610_, rst);
  or _47163_ (_39612_, _39611_, _39609_);
  or _47164_ (_41193_, _39612_, _39605_);
  and _47165_ (_39613_, _39116_, _30558_);
  nand _47166_ (_39614_, _39613_, _28510_);
  or _47167_ (_39615_, _39613_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _47168_ (_39616_, _39615_, _28576_);
  and _47169_ (_39617_, _39616_, _39614_);
  nor _47170_ (_39618_, _39125_, _38348_);
  and _47171_ (_39619_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47172_ (_39620_, _39619_, _39618_);
  and _47173_ (_39621_, _39620_, _27918_);
  and _47174_ (_39622_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47175_ (_39623_, _39622_, rst);
  or _47176_ (_39624_, _39623_, _39621_);
  or _47177_ (_41195_, _39624_, _39617_);
  and _47178_ (_39625_, _39116_, _31311_);
  nand _47179_ (_39626_, _39625_, _28510_);
  or _47180_ (_39627_, _39625_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _47181_ (_39628_, _39627_, _28576_);
  and _47182_ (_39629_, _39628_, _39626_);
  nor _47183_ (_39630_, _39125_, _38341_);
  and _47184_ (_39631_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47185_ (_39632_, _39631_, _39630_);
  and _47186_ (_39633_, _39632_, _27918_);
  and _47187_ (_39634_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47188_ (_39635_, _39634_, rst);
  or _47189_ (_39636_, _39635_, _39633_);
  or _47190_ (_41197_, _39636_, _39629_);
  and _47191_ (_39637_, _39116_, _32096_);
  nand _47192_ (_39638_, _39637_, _28510_);
  or _47193_ (_39639_, _39637_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47194_ (_39640_, _39639_, _28576_);
  and _47195_ (_39641_, _39640_, _39638_);
  nor _47196_ (_39642_, _39125_, _38334_);
  and _47197_ (_39643_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47198_ (_39644_, _39643_, _39642_);
  and _47199_ (_39645_, _39644_, _27918_);
  and _47200_ (_39646_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47201_ (_39647_, _39646_, rst);
  or _47202_ (_39648_, _39647_, _39645_);
  or _47203_ (_41198_, _39648_, _39641_);
  and _47204_ (_39649_, _39116_, _32901_);
  nand _47205_ (_39650_, _39649_, _28510_);
  or _47206_ (_39651_, _39649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _47207_ (_39652_, _39651_, _28576_);
  and _47208_ (_39653_, _39652_, _39650_);
  nor _47209_ (_39654_, _39125_, _38292_);
  and _47210_ (_39655_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47211_ (_39656_, _39655_, _39654_);
  and _47212_ (_39657_, _39656_, _27918_);
  and _47213_ (_39658_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47214_ (_39666_, _39658_, rst);
  or _47215_ (_39667_, _39666_, _39657_);
  or _47216_ (_41200_, _39667_, _39653_);
  and _47217_ (_39668_, _39116_, _33631_);
  nand _47218_ (_39669_, _39668_, _28510_);
  or _47219_ (_39670_, _39668_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _47220_ (_39671_, _39670_, _28576_);
  and _47221_ (_39672_, _39671_, _39669_);
  nor _47222_ (_39673_, _39125_, _38217_);
  and _47223_ (_39674_, _39125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47224_ (_39675_, _39674_, _39673_);
  and _47225_ (_39676_, _39675_, _27918_);
  and _47226_ (_39677_, _27907_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47227_ (_39678_, _39677_, rst);
  or _47228_ (_39679_, _39678_, _39676_);
  or _47229_ (_41202_, _39679_, _39672_);
  nor _47230_ (_39680_, _25105_, _24931_);
  and _47231_ (_39681_, _39680_, _39098_);
  and _47232_ (_39682_, _39681_, _38760_);
  and _47233_ (_39683_, _39682_, _28543_);
  nand _47234_ (_39684_, _39683_, _28510_);
  and _47235_ (_39685_, _38770_, _24942_);
  and _47236_ (_39686_, _39685_, _39123_);
  not _47237_ (_39687_, _39686_);
  or _47238_ (_39688_, _39683_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _47239_ (_39689_, _39688_, _39687_);
  and _47240_ (_39690_, _39689_, _39684_);
  nor _47241_ (_39691_, _39687_, _38386_);
  or _47242_ (_39692_, _39691_, _39690_);
  and _47243_ (_41698_, _39692_, _41755_);
  and _47244_ (_39693_, _25105_, _24942_);
  and _47245_ (_39694_, _39693_, _38760_);
  and _47246_ (_39695_, _39694_, _39098_);
  and _47247_ (_39696_, _39695_, _28543_);
  nand _47248_ (_39697_, _39696_, _28510_);
  and _47249_ (_39698_, _39685_, _39106_);
  not _47250_ (_39699_, _39698_);
  or _47251_ (_39700_, _39696_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47252_ (_39701_, _39700_, _39699_);
  and _47253_ (_39702_, _39701_, _39697_);
  nor _47254_ (_39703_, _39699_, _38386_);
  or _47255_ (_39704_, _39703_, _39702_);
  and _47256_ (_41701_, _39704_, _41755_);
  or _47257_ (_39705_, _24276_, _30547_);
  and _47258_ (_39706_, _39705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47259_ (_39707_, _39706_, _38911_);
  and _47260_ (_39708_, _39694_, _37975_);
  and _47261_ (_39713_, _39708_, _39707_);
  and _47262_ (_39714_, _39685_, _37997_);
  nand _47263_ (_39715_, _39708_, _24265_);
  and _47264_ (_39716_, _39715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47265_ (_39717_, _39716_, _39714_);
  or _47266_ (_39718_, _39717_, _39713_);
  nand _47267_ (_39719_, _39714_, _38217_);
  and _47268_ (_39720_, _39719_, _41755_);
  and _47269_ (_41702_, _39720_, _39718_);
  not _47270_ (_39721_, _39714_);
  not _47271_ (_39722_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _47272_ (_39723_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _47273_ (_39724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47274_ (_39725_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39724_);
  and _47275_ (_39726_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47276_ (_39727_, _39726_, _39725_);
  nor _47277_ (_39737_, _39727_, _39723_);
  or _47278_ (_39738_, _39737_, _39722_);
  and _47279_ (_39739_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _47280_ (_39740_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _47281_ (_39741_, _39740_, _39739_);
  nor _47282_ (_39742_, _39741_, _39723_);
  and _47283_ (_39743_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39724_);
  and _47284_ (_39744_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47285_ (_39745_, _39744_, _39743_);
  nand _47286_ (_39746_, _39745_, _39742_);
  or _47287_ (_39747_, _39746_, _39738_);
  and _47288_ (_39748_, _39747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor _47289_ (_39749_, _24018_, _24931_);
  and _47290_ (_39750_, _28576_, _28532_);
  and _47291_ (_39751_, _39750_, _37997_);
  and _47292_ (_39752_, _39751_, _39749_);
  or _47293_ (_39753_, _39752_, _39748_);
  and _47294_ (_39754_, _39753_, _39721_);
  nand _47295_ (_39755_, _39752_, _28510_);
  and _47296_ (_39756_, _39755_, _39754_);
  nor _47297_ (_39757_, _39721_, _38386_);
  or _47298_ (_39758_, _39757_, _39756_);
  and _47299_ (_41705_, _39758_, _41755_);
  nor _47300_ (_39759_, _39745_, _39723_);
  nand _47301_ (_39760_, _39759_, _39741_);
  or _47302_ (_39761_, _39760_, _39738_);
  and _47303_ (_39762_, _39761_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _47304_ (_39763_, _28576_, _29813_);
  and _47305_ (_39764_, _39763_, _37997_);
  and _47306_ (_39765_, _39764_, _39749_);
  or _47307_ (_39766_, _39765_, _39762_);
  and _47308_ (_39767_, _39766_, _39721_);
  nand _47309_ (_39768_, _39765_, _28510_);
  and _47310_ (_39769_, _39768_, _39767_);
  nor _47311_ (_39770_, _39721_, _38292_);
  or _47312_ (_39771_, _39770_, _39769_);
  and _47313_ (_41707_, _39771_, _41755_);
  not _47314_ (_39772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _47315_ (_39773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _39772_);
  nand _47316_ (_39774_, _39737_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _47317_ (_39775_, _39759_, _39742_);
  or _47318_ (_39776_, _39775_, _39774_);
  and _47319_ (_39777_, _39776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _47320_ (_39778_, _39777_, _39773_);
  nor _47321_ (_39779_, _28521_, _24931_);
  and _47322_ (_39780_, _39764_, _39779_);
  or _47323_ (_39781_, _39780_, _39778_);
  and _47324_ (_39782_, _39781_, _39721_);
  nand _47325_ (_39783_, _39780_, _28510_);
  and _47326_ (_39784_, _39783_, _39782_);
  nor _47327_ (_39785_, _39721_, _38355_);
  or _47328_ (_39786_, _39785_, _39784_);
  and _47329_ (_41709_, _39786_, _41755_);
  and _47330_ (_39787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _47331_ (_39788_, _39774_, _39760_);
  and _47332_ (_39789_, _39788_, _39787_);
  and _47333_ (_39790_, _39751_, _39779_);
  or _47334_ (_39791_, _39790_, _39789_);
  and _47335_ (_39792_, _39791_, _39721_);
  nand _47336_ (_39793_, _39790_, _28510_);
  and _47337_ (_39794_, _39793_, _39792_);
  nor _47338_ (_39795_, _39721_, _38341_);
  or _47339_ (_39796_, _39795_, _39794_);
  and _47340_ (_41711_, _39796_, _41755_);
  and _47341_ (_39797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47342_ (_39798_, _39797_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _47343_ (_39799_, _39798_);
  and _47344_ (_39800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47345_ (_39801_, _39800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47346_ (_39802_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47347_ (_39803_, _39802_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _47348_ (_39804_, _39803_, _39801_);
  and _47349_ (_39805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _47350_ (_39806_, _39805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  not _47351_ (_39807_, _39806_);
  and _47352_ (_39808_, _39807_, _39804_);
  and _47353_ (_39809_, _39808_, _39799_);
  not _47354_ (_39810_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47355_ (_39811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47356_ (_39812_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39724_);
  or _47357_ (_39813_, _39812_, _39811_);
  nor _47358_ (_39814_, _39813_, _39810_);
  nor _47359_ (_39815_, _39814_, _39723_);
  nor _47360_ (_39816_, _39815_, _39809_);
  and _47361_ (_39817_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _47362_ (_39818_, _39817_, _39724_);
  and _47363_ (_39819_, _39818_, _39816_);
  and _47364_ (_39820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39723_);
  not _47365_ (_39821_, _39820_);
  not _47366_ (_39822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47367_ (_39823_, _39800_, _39822_);
  not _47368_ (_39824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47369_ (_39825_, _39802_, _39824_);
  nor _47370_ (_39826_, _39825_, _39823_);
  not _47371_ (_39827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _47372_ (_39828_, _39805_, _39827_);
  not _47373_ (_39829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _47374_ (_39830_, _39797_, _39829_);
  nor _47375_ (_39831_, _39830_, _39828_);
  and _47376_ (_39832_, _39831_, _39826_);
  nor _47377_ (_39833_, _39832_, _39821_);
  nand _47378_ (_39834_, _39833_, _39818_);
  and _47379_ (_39835_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41755_);
  nand _47380_ (_39836_, _39835_, _39834_);
  nor _47381_ (_41743_, _39836_, _39819_);
  nor _47382_ (_39837_, _39817_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _47383_ (_39838_, _39837_);
  nor _47384_ (_39839_, _39833_, _39816_);
  nor _47385_ (_39840_, _39839_, _39838_);
  nand _47386_ (_39841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41755_);
  nor _47387_ (_41744_, _39841_, _39840_);
  and _47388_ (_39842_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _47389_ (_39843_, _39804_);
  or _47390_ (_39844_, _39843_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _47391_ (_39845_, _39844_, _39842_);
  or _47392_ (_39846_, _39808_, _39739_);
  and _47393_ (_39847_, _39846_, _39845_);
  and _47394_ (_39848_, _39847_, _39816_);
  or _47395_ (_39849_, _39848_, _39817_);
  and _47396_ (_39850_, _39839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _47397_ (_39851_, _39816_);
  and _47398_ (_39852_, _39833_, _39851_);
  and _47399_ (_39853_, _39830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47400_ (_39854_, _39853_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _47401_ (_39855_, _39826_);
  and _47402_ (_39856_, _39828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47403_ (_39857_, _39856_, _39855_);
  and _47404_ (_39858_, _39857_, _39854_);
  and _47405_ (_39859_, _39855_, _39739_);
  or _47406_ (_39860_, _39859_, _39858_);
  and _47407_ (_39861_, _39860_, _39852_);
  or _47408_ (_39862_, _39861_, _39850_);
  or _47409_ (_39863_, _39862_, _39849_);
  not _47410_ (_39864_, _39817_);
  or _47411_ (_39865_, _39864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _47412_ (_39866_, _39865_, _41755_);
  and _47413_ (_41746_, _39866_, _39863_);
  and _47414_ (_39867_, _39798_, _39724_);
  or _47415_ (_39868_, _39843_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _47416_ (_39869_, _39868_, _39867_);
  or _47417_ (_39870_, _39808_, _39740_);
  and _47418_ (_39871_, _39870_, _39869_);
  and _47419_ (_39872_, _39871_, _39816_);
  or _47420_ (_39873_, _39872_, _39817_);
  and _47421_ (_39874_, _39839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47422_ (_39875_, _39830_, _39724_);
  or _47423_ (_39876_, _39875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47424_ (_39877_, _39828_, _39724_);
  nor _47425_ (_39878_, _39877_, _39855_);
  and _47426_ (_39879_, _39878_, _39876_);
  and _47427_ (_39880_, _39855_, _39740_);
  or _47428_ (_39881_, _39880_, _39879_);
  and _47429_ (_39882_, _39881_, _39852_);
  or _47430_ (_39883_, _39882_, _39874_);
  or _47431_ (_39884_, _39883_, _39873_);
  or _47432_ (_39885_, _39864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47433_ (_39886_, _39885_, _41755_);
  and _47434_ (_41748_, _39886_, _39884_);
  nand _47435_ (_39887_, _39839_, _39723_);
  nor _47436_ (_39888_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _47437_ (_39889_, _39888_, _39817_);
  and _47438_ (_39890_, _39889_, _41755_);
  and _47439_ (_41750_, _39890_, _39887_);
  and _47440_ (_39891_, _39839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _47441_ (_39892_, _39724_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _47442_ (_39893_, _39892_, _39888_);
  nor _47443_ (_39894_, _39893_, _39851_);
  or _47444_ (_39895_, _39894_, _39817_);
  or _47445_ (_39896_, _39895_, _39891_);
  or _47446_ (_39897_, _39893_, _39864_);
  and _47447_ (_39898_, _39897_, _41755_);
  and _47448_ (_41752_, _39898_, _39896_);
  and _47449_ (_39899_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41755_);
  and _47450_ (_41754_, _39899_, _39817_);
  nor _47451_ (_39900_, _39839_, _39817_);
  and _47452_ (_39901_, _39817_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _47453_ (_39902_, _39901_, _39900_);
  and _47454_ (_42678_, _39902_, _41755_);
  and _47455_ (_39903_, _39817_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _47456_ (_39904_, _39903_, _39900_);
  and _47457_ (_42680_, _39904_, _41755_);
  and _47458_ (_39905_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _41755_);
  and _47459_ (_42682_, _39905_, _39817_);
  not _47460_ (_39906_, _39823_);
  nor _47461_ (_39907_, _39830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _47462_ (_39908_, _39907_, _39828_);
  or _47463_ (_39909_, _39908_, _39825_);
  and _47464_ (_39910_, _39909_, _39906_);
  and _47465_ (_39911_, _39910_, _39852_);
  not _47466_ (_39912_, _39801_);
  or _47467_ (_39913_, _39798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _47468_ (_39914_, _39913_, _39807_);
  or _47469_ (_39915_, _39914_, _39803_);
  and _47470_ (_39916_, _39915_, _39912_);
  and _47471_ (_39917_, _39916_, _39816_);
  or _47472_ (_39918_, _39917_, _39817_);
  or _47473_ (_39919_, _39918_, _39911_);
  or _47474_ (_39920_, _39864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _47475_ (_39921_, _39920_, _41755_);
  and _47476_ (_42684_, _39921_, _39919_);
  nand _47477_ (_39922_, _39826_, _39820_);
  nor _47478_ (_39923_, _39922_, _39831_);
  or _47479_ (_39924_, _39923_, _39816_);
  nand _47480_ (_39925_, _39816_, _39843_);
  and _47481_ (_39926_, _39925_, _39924_);
  or _47482_ (_39927_, _39926_, _39817_);
  or _47483_ (_39928_, _39864_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _47484_ (_39929_, _39928_, _41755_);
  and _47485_ (_42686_, _39929_, _39927_);
  and _47486_ (_39930_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _41755_);
  and _47487_ (_42688_, _39930_, _39817_);
  and _47488_ (_39931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _41755_);
  and _47489_ (_42690_, _39931_, _39817_);
  nand _47490_ (_39932_, _39839_, _39837_);
  nor _47491_ (_39933_, _39817_, _39816_);
  or _47492_ (_39934_, _39933_, _39724_);
  and _47493_ (_39935_, _39934_, _41755_);
  and _47494_ (_42692_, _39935_, _39932_);
  not _47495_ (_39936_, _39900_);
  and _47496_ (_39937_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _47497_ (_39938_, _39867_);
  and _47498_ (_39939_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _47499_ (_39940_, _39806_, _39724_);
  or _47500_ (_39941_, _39940_, _39803_);
  or _47501_ (_39942_, _39941_, _39939_);
  not _47502_ (_39943_, _39803_);
  or _47503_ (_39944_, _39943_, _39726_);
  and _47504_ (_39945_, _39944_, _39942_);
  or _47505_ (_39946_, _39945_, _39801_);
  or _47506_ (_39947_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39724_);
  or _47507_ (_39948_, _39947_, _39912_);
  and _47508_ (_39949_, _39948_, _39816_);
  and _47509_ (_39950_, _39949_, _39946_);
  not _47510_ (_39951_, _39875_);
  and _47511_ (_39952_, _39951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _47512_ (_39953_, _39877_, _39825_);
  or _47513_ (_39954_, _39953_, _39952_);
  not _47514_ (_39955_, _39825_);
  or _47515_ (_39956_, _39955_, _39726_);
  and _47516_ (_39957_, _39956_, _39906_);
  and _47517_ (_39958_, _39957_, _39954_);
  and _47518_ (_39959_, _39947_, _39823_);
  or _47519_ (_39960_, _39959_, _39958_);
  and _47520_ (_39961_, _39960_, _39852_);
  or _47521_ (_39962_, _39961_, _39950_);
  and _47522_ (_39963_, _39962_, _39864_);
  or _47523_ (_39964_, _39963_, _39937_);
  and _47524_ (_42694_, _39964_, _41755_);
  and _47525_ (_39965_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _47526_ (_39966_, _39938_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _47527_ (_39967_, _39966_, _39941_);
  or _47528_ (_39968_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39724_);
  or _47529_ (_39969_, _39968_, _39943_);
  and _47530_ (_39970_, _39969_, _39912_);
  and _47531_ (_39971_, _39970_, _39967_);
  and _47532_ (_39972_, _39801_, _39744_);
  or _47533_ (_39973_, _39972_, _39971_);
  and _47534_ (_39974_, _39973_, _39816_);
  and _47535_ (_39975_, _39951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _47536_ (_39976_, _39975_, _39953_);
  or _47537_ (_39977_, _39968_, _39955_);
  and _47538_ (_39978_, _39977_, _39906_);
  and _47539_ (_39979_, _39978_, _39976_);
  and _47540_ (_39980_, _39823_, _39744_);
  or _47541_ (_39981_, _39980_, _39979_);
  and _47542_ (_39982_, _39981_, _39852_);
  or _47543_ (_39983_, _39982_, _39974_);
  and _47544_ (_39984_, _39983_, _39864_);
  or _47545_ (_39985_, _39984_, _39965_);
  and _47546_ (_42696_, _39985_, _41755_);
  and _47547_ (_39986_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not _47548_ (_39987_, _39842_);
  and _47549_ (_39988_, _39987_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _47550_ (_39989_, _39806_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47551_ (_39990_, _39989_, _39803_);
  or _47552_ (_39991_, _39990_, _39988_);
  or _47553_ (_39992_, _39943_, _39725_);
  and _47554_ (_39993_, _39992_, _39991_);
  or _47555_ (_39994_, _39993_, _39801_);
  or _47556_ (_39995_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47557_ (_39996_, _39995_, _39912_);
  and _47558_ (_39997_, _39996_, _39816_);
  and _47559_ (_39998_, _39997_, _39994_);
  not _47560_ (_39999_, _39853_);
  and _47561_ (_40000_, _39999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _47562_ (_40001_, _39856_, _39825_);
  or _47563_ (_40002_, _40001_, _40000_);
  or _47564_ (_40003_, _39955_, _39725_);
  and _47565_ (_40004_, _40003_, _39906_);
  and _47566_ (_40005_, _40004_, _40002_);
  and _47567_ (_40006_, _39995_, _39823_);
  or _47568_ (_40007_, _40006_, _40005_);
  and _47569_ (_40008_, _40007_, _39852_);
  or _47570_ (_40009_, _40008_, _39998_);
  and _47571_ (_40010_, _40009_, _39864_);
  or _47572_ (_40011_, _40010_, _39986_);
  and _47573_ (_42698_, _40011_, _41755_);
  and _47574_ (_40012_, _39936_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _47575_ (_40013_, _39987_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _47576_ (_40014_, _40013_, _39990_);
  or _47577_ (_40015_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _47578_ (_40016_, _40015_, _39943_);
  and _47579_ (_40017_, _40016_, _39912_);
  and _47580_ (_40018_, _40017_, _40014_);
  and _47581_ (_40019_, _39801_, _39743_);
  or _47582_ (_40020_, _40019_, _40018_);
  and _47583_ (_40021_, _40020_, _39816_);
  and _47584_ (_40022_, _39999_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _47585_ (_40023_, _40022_, _40001_);
  or _47586_ (_40024_, _40015_, _39955_);
  and _47587_ (_40025_, _40024_, _39906_);
  and _47588_ (_40026_, _40025_, _40023_);
  and _47589_ (_40027_, _39823_, _39743_);
  or _47590_ (_40028_, _40027_, _40026_);
  and _47591_ (_40029_, _40028_, _39852_);
  or _47592_ (_40030_, _40029_, _40021_);
  and _47593_ (_40031_, _40030_, _39864_);
  or _47594_ (_40032_, _40031_, _40012_);
  and _47595_ (_42700_, _40032_, _41755_);
  and _47596_ (_40033_, _39837_, _39816_);
  nand _47597_ (_40034_, _39837_, _39833_);
  and _47598_ (_40035_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _47599_ (_40036_, _40035_, _40033_);
  and _47600_ (_42702_, _40036_, _41755_);
  and _47601_ (_40037_, _39834_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _47602_ (_40038_, _40037_, _39819_);
  and _47603_ (_42704_, _40038_, _41755_);
  and _47604_ (_40039_, _39708_, _24287_);
  or _47605_ (_40040_, _40039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _47606_ (_40041_, _40040_, _39721_);
  nand _47607_ (_40042_, _40039_, _28510_);
  and _47608_ (_40043_, _40042_, _40041_);
  and _47609_ (_40044_, _39714_, _38365_);
  or _47610_ (_40045_, _40044_, _40043_);
  and _47611_ (_42706_, _40045_, _41755_);
  and _47612_ (_40046_, _39708_, _30558_);
  nand _47613_ (_40047_, _40046_, _28510_);
  or _47614_ (_40048_, _40046_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _47615_ (_40049_, _40048_, _39721_);
  and _47616_ (_40050_, _40049_, _40047_);
  nor _47617_ (_40051_, _39721_, _38348_);
  or _47618_ (_40052_, _40051_, _40050_);
  and _47619_ (_42708_, _40052_, _41755_);
  and _47620_ (_40053_, _39708_, _32096_);
  nand _47621_ (_40054_, _40053_, _28510_);
  or _47622_ (_40055_, _40053_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _47623_ (_40056_, _40055_, _39721_);
  and _47624_ (_40057_, _40056_, _40054_);
  nor _47625_ (_40058_, _39721_, _38334_);
  or _47626_ (_40059_, _40058_, _40057_);
  and _47627_ (_42709_, _40059_, _41755_);
  and _47628_ (_40060_, _39695_, _24287_);
  nand _47629_ (_40061_, _40060_, _28510_);
  or _47630_ (_40062_, _40060_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47631_ (_40063_, _40062_, _39699_);
  and _47632_ (_40064_, _40063_, _40061_);
  and _47633_ (_40065_, _39698_, _38365_);
  or _47634_ (_40066_, _40065_, _40064_);
  and _47635_ (_42711_, _40066_, _41755_);
  and _47636_ (_40067_, _39695_, _29824_);
  nand _47637_ (_40068_, _40067_, _28510_);
  or _47638_ (_40069_, _40067_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47639_ (_40070_, _40069_, _39699_);
  and _47640_ (_40071_, _40070_, _40068_);
  nor _47641_ (_40072_, _39699_, _38355_);
  or _47642_ (_40073_, _40072_, _40071_);
  and _47643_ (_42713_, _40073_, _41755_);
  and _47644_ (_40074_, _30590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _47645_ (_40075_, _40074_, _30580_);
  and _47646_ (_40076_, _40075_, _39695_);
  nand _47647_ (_40077_, _39695_, _39285_);
  and _47648_ (_40078_, _40077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _47649_ (_40079_, _40078_, _39698_);
  or _47650_ (_40080_, _40079_, _40076_);
  nand _47651_ (_40081_, _39698_, _38348_);
  and _47652_ (_40082_, _40081_, _41755_);
  and _47653_ (_42715_, _40082_, _40080_);
  and _47654_ (_40083_, _39695_, _31311_);
  nand _47655_ (_40084_, _40083_, _28510_);
  or _47656_ (_40085_, _40083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47657_ (_40086_, _40085_, _39699_);
  and _47658_ (_40087_, _40086_, _40084_);
  nor _47659_ (_40088_, _39699_, _38341_);
  or _47660_ (_40089_, _40088_, _40087_);
  and _47661_ (_42717_, _40089_, _41755_);
  and _47662_ (_40090_, _39695_, _32096_);
  nand _47663_ (_40091_, _40090_, _28510_);
  or _47664_ (_40092_, _40090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _47665_ (_40093_, _40092_, _39699_);
  and _47666_ (_40094_, _40093_, _40091_);
  nor _47667_ (_40095_, _39699_, _38334_);
  or _47668_ (_40096_, _40095_, _40094_);
  and _47669_ (_42719_, _40096_, _41755_);
  and _47670_ (_40097_, _39695_, _32901_);
  nand _47671_ (_40098_, _40097_, _28510_);
  or _47672_ (_40099_, _40097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _47673_ (_40100_, _40099_, _39699_);
  and _47674_ (_40101_, _40100_, _40098_);
  nor _47675_ (_40102_, _39699_, _38292_);
  or _47676_ (_40103_, _40102_, _40101_);
  and _47677_ (_42721_, _40103_, _41755_);
  and _47678_ (_40104_, _39695_, _33631_);
  nand _47679_ (_40105_, _40104_, _28510_);
  or _47680_ (_40106_, _40104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _47681_ (_40107_, _40106_, _39699_);
  and _47682_ (_40108_, _40107_, _40105_);
  nor _47683_ (_40109_, _39699_, _38217_);
  or _47684_ (_40110_, _40109_, _40108_);
  and _47685_ (_42723_, _40110_, _41755_);
  and _47686_ (_40111_, _39682_, _24287_);
  nand _47687_ (_40112_, _40111_, _28510_);
  or _47688_ (_40113_, _40111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47689_ (_40114_, _40113_, _39687_);
  and _47690_ (_40115_, _40114_, _40112_);
  and _47691_ (_40116_, _39686_, _38365_);
  or _47692_ (_40117_, _40116_, _40115_);
  and _47693_ (_42725_, _40117_, _41755_);
  and _47694_ (_40118_, _39682_, _29824_);
  nand _47695_ (_40119_, _40118_, _28510_);
  or _47696_ (_40120_, _40118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47697_ (_40121_, _40120_, _39687_);
  and _47698_ (_40122_, _40121_, _40119_);
  nor _47699_ (_40123_, _39687_, _38355_);
  or _47700_ (_40124_, _40123_, _40122_);
  and _47701_ (_42727_, _40124_, _41755_);
  and _47702_ (_40125_, _30590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _47703_ (_40126_, _40125_, _30580_);
  and _47704_ (_40127_, _40126_, _39682_);
  nand _47705_ (_40128_, _39682_, _39285_);
  and _47706_ (_40129_, _40128_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _47707_ (_40130_, _40129_, _39686_);
  or _47708_ (_40131_, _40130_, _40127_);
  nand _47709_ (_40132_, _39686_, _38348_);
  and _47710_ (_40133_, _40132_, _41755_);
  and _47711_ (_42729_, _40133_, _40131_);
  and _47712_ (_40134_, _39682_, _31311_);
  nand _47713_ (_40135_, _40134_, _28510_);
  or _47714_ (_40136_, _40134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _47715_ (_40137_, _40136_, _39687_);
  and _47716_ (_40138_, _40137_, _40135_);
  nor _47717_ (_40139_, _39687_, _38341_);
  or _47718_ (_40140_, _40139_, _40138_);
  and _47719_ (_42731_, _40140_, _41755_);
  and _47720_ (_40141_, _39682_, _32096_);
  nand _47721_ (_40142_, _40141_, _28510_);
  or _47722_ (_40143_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _47723_ (_40144_, _40143_, _39687_);
  and _47724_ (_40145_, _40144_, _40142_);
  nor _47725_ (_40146_, _39687_, _38334_);
  or _47726_ (_40147_, _40146_, _40145_);
  and _47727_ (_42733_, _40147_, _41755_);
  and _47728_ (_40148_, _39682_, _32901_);
  nand _47729_ (_40149_, _40148_, _28510_);
  or _47730_ (_40150_, _40148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _47731_ (_40151_, _40150_, _39687_);
  and _47732_ (_40152_, _40151_, _40149_);
  nor _47733_ (_40153_, _39687_, _38292_);
  or _47734_ (_40154_, _40153_, _40152_);
  and _47735_ (_42735_, _40154_, _41755_);
  and _47736_ (_40155_, _39682_, _33631_);
  nand _47737_ (_40156_, _40155_, _28510_);
  or _47738_ (_40157_, _40155_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _47739_ (_40158_, _40157_, _39687_);
  and _47740_ (_40159_, _40158_, _40156_);
  nor _47741_ (_40160_, _39687_, _38217_);
  or _47742_ (_40161_, _40160_, _40159_);
  and _47743_ (_42737_, _40161_, _41755_);
  and _47744_ (_40162_, _38388_, _37789_);
  not _47745_ (_40163_, _40162_);
  not _47746_ (_40164_, _36788_);
  and _47747_ (_40165_, _37778_, _40164_);
  nor _47748_ (_40166_, _38773_, _38851_);
  nor _47749_ (_40167_, _40166_, _38857_);
  nor _47750_ (_40168_, _40167_, _34229_);
  and _47751_ (_40169_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  not _47752_ (_40170_, _40169_);
  and _47753_ (_40171_, _40167_, _34240_);
  and _47754_ (_40172_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _47755_ (_40173_, _40167_, _34240_);
  and _47756_ (_40174_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor _47757_ (_40175_, _40174_, _40172_);
  and _47758_ (_40176_, _40175_, _40170_);
  nand _47759_ (_40177_, _34229_, _29802_);
  or _47760_ (_40178_, _34229_, _29802_);
  nor _47761_ (_40179_, _24778_, _23822_);
  nor _47762_ (_40180_, _40179_, _27885_);
  not _47763_ (_40181_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _47764_ (_40182_, _30590_, _40181_);
  and _47765_ (_40183_, _40182_, _40180_);
  and _47766_ (_40184_, _40183_, _40178_);
  and _47767_ (_40185_, _40184_, _40177_);
  and _47768_ (_40186_, _40167_, _24942_);
  nor _47769_ (_40187_, _40167_, _24942_);
  nor _47770_ (_40188_, _40187_, _40186_);
  and _47771_ (_40189_, _40188_, _40185_);
  and _47772_ (_40190_, _40167_, _34229_);
  and _47773_ (_40191_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _47774_ (_40192_, _40191_, _40189_);
  and _47775_ (_40193_, _40192_, _40176_);
  and _47776_ (_40194_, _40189_, _38386_);
  or _47777_ (_40195_, _40194_, _40193_);
  not _47778_ (_40196_, _40195_);
  and _47779_ (_40197_, _40196_, _40165_);
  nor _47780_ (_40198_, _37778_, _40164_);
  not _47781_ (_40199_, _33793_);
  and _47782_ (_40200_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _47783_ (_40201_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _47784_ (_40202_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _47785_ (_40203_, _40202_, _40201_);
  and _47786_ (_40204_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _47787_ (_40205_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _47788_ (_40206_, _40205_, _40204_);
  and _47789_ (_40207_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _47790_ (_40208_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _47791_ (_40209_, _40208_, _40207_);
  and _47792_ (_40210_, _40209_, _40206_);
  and _47793_ (_40211_, _40210_, _40203_);
  and _47794_ (_40212_, _34251_, _33793_);
  not _47795_ (_40213_, _40212_);
  nor _47796_ (_40214_, _40213_, _40211_);
  nor _47797_ (_40215_, _40214_, _40200_);
  not _47798_ (_40216_, _40215_);
  and _47799_ (_40217_, _40216_, _40198_);
  nor _47800_ (_40218_, _40217_, _40197_);
  and _47801_ (_40219_, _40218_, _37932_);
  and _47802_ (_40220_, _40219_, _40163_);
  nor _47803_ (_40221_, _37519_, _37180_);
  nor _47804_ (_40222_, _37341_, _37310_);
  nor _47805_ (_40223_, _37442_, _37279_);
  and _47806_ (_40224_, _40223_, _40222_);
  and _47807_ (_40225_, _37508_, _37374_);
  and _47808_ (_40226_, _40225_, _40224_);
  and _47809_ (_40227_, _40226_, _40221_);
  nor _47810_ (_40228_, _40227_, _33750_);
  and _47811_ (_40229_, _37126_, _36174_);
  nor _47812_ (_40230_, _37690_, _40229_);
  nor _47813_ (_40231_, _40230_, _37657_);
  nor _47814_ (_40232_, _40231_, _40228_);
  not _47815_ (_40233_, _40232_);
  and _47816_ (_40234_, _40233_, _40220_);
  and _47817_ (_40235_, _40165_, _37932_);
  not _47818_ (_40236_, _38292_);
  and _47819_ (_40237_, _40189_, _40236_);
  and _47820_ (_40238_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _47821_ (_40239_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _47822_ (_40240_, _40239_, _40238_);
  and _47823_ (_40241_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and _47824_ (_40242_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _47825_ (_40243_, _40242_, _40241_);
  and _47826_ (_40244_, _40243_, _40240_);
  nor _47827_ (_40245_, _40244_, _40189_);
  nor _47828_ (_40246_, _40245_, _40237_);
  not _47829_ (_40247_, _40246_);
  and _47830_ (_40248_, _40247_, _40235_);
  not _47831_ (_40249_, _40198_);
  nor _47832_ (_40250_, _40165_, _37932_);
  and _47833_ (_40251_, _40250_, _40249_);
  nor _47834_ (_40252_, _40251_, _40248_);
  and _47835_ (_40253_, _37932_, _37789_);
  not _47836_ (_40254_, _38426_);
  and _47837_ (_40255_, _40254_, _40253_);
  and _47838_ (_40256_, _40198_, _37932_);
  and _47839_ (_40257_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _47840_ (_40258_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _47841_ (_40259_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _47842_ (_40260_, _40259_, _40258_);
  and _47843_ (_40261_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _47844_ (_40262_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _47845_ (_40263_, _40262_, _40261_);
  and _47846_ (_40264_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _47847_ (_40265_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _47848_ (_40266_, _40265_, _40264_);
  and _47849_ (_40267_, _40266_, _40263_);
  and _47850_ (_40268_, _40267_, _40260_);
  nor _47851_ (_40269_, _40268_, _40213_);
  nor _47852_ (_40270_, _40269_, _40257_);
  not _47853_ (_40271_, _40270_);
  and _47854_ (_40272_, _40271_, _40256_);
  nor _47855_ (_40273_, _40272_, _40255_);
  and _47856_ (_40274_, _40273_, _40252_);
  not _47857_ (_40275_, _40274_);
  and _47858_ (_40276_, _40275_, _40234_);
  and _47859_ (_40277_, _37778_, _36788_);
  and _47860_ (_40278_, _40277_, _37932_);
  and _47861_ (_40279_, _40278_, _36831_);
  and _47862_ (_40280_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _47863_ (_40281_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _47864_ (_40282_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _47865_ (_40283_, _40282_, _40281_);
  and _47866_ (_40284_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _47867_ (_40285_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _47868_ (_40286_, _40285_, _40284_);
  and _47869_ (_40287_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _47870_ (_40288_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _47871_ (_40289_, _40288_, _40287_);
  and _47872_ (_40290_, _40289_, _40286_);
  and _47873_ (_40291_, _40290_, _40283_);
  nor _47874_ (_40292_, _40291_, _40213_);
  nor _47875_ (_40293_, _40292_, _40280_);
  not _47876_ (_40294_, _40293_);
  and _47877_ (_40295_, _40294_, _40256_);
  nor _47878_ (_40296_, _40295_, _40279_);
  not _47879_ (_40297_, _38408_);
  and _47880_ (_40298_, _40297_, _40253_);
  and _47881_ (_40299_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _47882_ (_40300_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _47883_ (_40301_, _40300_, _40299_);
  and _47884_ (_40302_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _47885_ (_40303_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _47886_ (_40304_, _40303_, _40302_);
  and _47887_ (_40305_, _40304_, _40301_);
  nor _47888_ (_40306_, _40305_, _40189_);
  not _47889_ (_40307_, _38348_);
  and _47890_ (_40308_, _40189_, _40307_);
  nor _47891_ (_40309_, _40308_, _40306_);
  not _47892_ (_40310_, _40309_);
  and _47893_ (_40311_, _40310_, _40235_);
  nor _47894_ (_40312_, _40311_, _40298_);
  and _47895_ (_40313_, _40312_, _40296_);
  nor _47896_ (_40314_, _40313_, _40233_);
  nor _47897_ (_40315_, _40314_, _40276_);
  and _47898_ (_40316_, _24778_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _47899_ (_40317_, _40316_, _38936_);
  nor _47900_ (_40318_, _24018_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _47901_ (_40319_, _40318_, _40317_);
  not _47902_ (_40320_, _40319_);
  and _47903_ (_40321_, _40320_, _40315_);
  and _47904_ (_40322_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _47905_ (_40323_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _47906_ (_40324_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _47907_ (_40325_, _40324_, _40323_);
  and _47908_ (_40326_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _47909_ (_40327_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _47910_ (_40328_, _40327_, _40326_);
  and _47911_ (_40329_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _47912_ (_40330_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _47913_ (_40331_, _40330_, _40329_);
  and _47914_ (_40332_, _40331_, _40328_);
  and _47915_ (_40333_, _40332_, _40325_);
  nor _47916_ (_40334_, _40333_, _40213_);
  nor _47917_ (_40335_, _40334_, _40322_);
  not _47918_ (_40336_, _40335_);
  and _47919_ (_40337_, _40336_, _40256_);
  and _47920_ (_40338_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and _47921_ (_40339_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _47922_ (_40340_, _40339_, _40338_);
  and _47923_ (_40341_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _47924_ (_40342_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _47925_ (_40343_, _40342_, _40341_);
  and _47926_ (_40344_, _40343_, _40340_);
  nor _47927_ (_40345_, _40344_, _40189_);
  not _47928_ (_40346_, _38341_);
  and _47929_ (_40347_, _40189_, _40346_);
  nor _47930_ (_40348_, _40347_, _40345_);
  not _47931_ (_40349_, _40348_);
  and _47932_ (_40350_, _40349_, _40235_);
  nor _47933_ (_40351_, _40350_, _40337_);
  not _47934_ (_40352_, _38414_);
  and _47935_ (_40353_, _40352_, _40253_);
  not _47936_ (_40354_, _40167_);
  and _47937_ (_40355_, _40278_, _40354_);
  nor _47938_ (_40356_, _40355_, _40353_);
  and _47939_ (_40357_, _40356_, _40351_);
  not _47940_ (_40358_, _40357_);
  and _47941_ (_40359_, _40358_, _40234_);
  and _47942_ (_40360_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _47943_ (_40361_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _47944_ (_40362_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _47945_ (_40363_, _40362_, _40361_);
  and _47946_ (_40364_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _47947_ (_40365_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _47948_ (_40366_, _40365_, _40364_);
  and _47949_ (_40367_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _47950_ (_40368_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _47951_ (_40369_, _40368_, _40367_);
  and _47952_ (_40370_, _40369_, _40366_);
  and _47953_ (_40371_, _40370_, _40363_);
  nor _47954_ (_40372_, _40371_, _40213_);
  nor _47955_ (_40373_, _40372_, _40360_);
  not _47956_ (_40374_, _40373_);
  and _47957_ (_40375_, _40374_, _40256_);
  and _47958_ (_40376_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _47959_ (_40377_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _47960_ (_40378_, _40377_, _40376_);
  and _47961_ (_40379_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _47962_ (_40380_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _47963_ (_40381_, _40380_, _40379_);
  and _47964_ (_40382_, _40381_, _40378_);
  nor _47965_ (_40383_, _40382_, _40189_);
  and _47966_ (_40384_, _40189_, _38365_);
  nor _47967_ (_40385_, _40384_, _40383_);
  not _47968_ (_40386_, _40385_);
  and _47969_ (_40387_, _40386_, _40235_);
  nor _47970_ (_40388_, _40387_, _40375_);
  not _47971_ (_40389_, _38396_);
  and _47972_ (_40390_, _40389_, _40253_);
  and _47973_ (_40391_, _40278_, _34240_);
  nor _47974_ (_40392_, _40391_, _40390_);
  and _47975_ (_40393_, _40392_, _40388_);
  nor _47976_ (_40394_, _40393_, _40233_);
  nor _47977_ (_40395_, _40394_, _40359_);
  and _47978_ (_40396_, _40316_, _24942_);
  nor _47979_ (_40397_, _24265_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _47980_ (_40398_, _40397_, _40396_);
  not _47981_ (_40399_, _40398_);
  nor _47982_ (_40400_, _40399_, _40395_);
  nor _47983_ (_40401_, _40400_, _40321_);
  nor _47984_ (_40402_, _40320_, _40315_);
  not _47985_ (_40403_, _40402_);
  not _47986_ (_40404_, _38432_);
  and _47987_ (_40405_, _40404_, _40253_);
  not _47988_ (_40406_, _40405_);
  and _47989_ (_40407_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _47990_ (_40408_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _47991_ (_40409_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _47992_ (_40410_, _40409_, _40408_);
  and _47993_ (_40411_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _47994_ (_40412_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _47995_ (_40413_, _40412_, _40411_);
  and _47996_ (_40414_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _47997_ (_40415_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _47998_ (_40416_, _40415_, _40414_);
  and _47999_ (_40417_, _40416_, _40413_);
  and _48000_ (_40418_, _40417_, _40410_);
  nor _48001_ (_40419_, _40418_, _40213_);
  nor _48002_ (_40420_, _40419_, _40407_);
  not _48003_ (_40421_, _40420_);
  and _48004_ (_40422_, _40421_, _40256_);
  not _48005_ (_40423_, _40422_);
  and _48006_ (_40424_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and _48007_ (_40425_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _48008_ (_40426_, _40425_, _40424_);
  and _48009_ (_40427_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _48010_ (_40428_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _48011_ (_40429_, _40428_, _40427_);
  and _48012_ (_40430_, _40429_, _40426_);
  nor _48013_ (_40431_, _40430_, _40189_);
  not _48014_ (_40432_, _38217_);
  and _48015_ (_40433_, _40189_, _40432_);
  nor _48016_ (_40434_, _40433_, _40431_);
  not _48017_ (_40435_, _40434_);
  and _48018_ (_40436_, _40435_, _40235_);
  nor _48019_ (_40437_, _40436_, _40250_);
  and _48020_ (_40438_, _40437_, _40423_);
  and _48021_ (_40439_, _40438_, _40406_);
  and _48022_ (_40440_, _40439_, _40234_);
  nor _48023_ (_40441_, _40358_, _40234_);
  nor _48024_ (_40442_, _40441_, _40440_);
  nor _48025_ (_40443_, _40316_, _24942_);
  and _48026_ (_40444_, _40316_, _24494_);
  nor _48027_ (_40445_, _40444_, _40443_);
  not _48028_ (_40446_, _40445_);
  and _48029_ (_40447_, _40446_, _40442_);
  nor _48030_ (_40448_, _40446_, _40442_);
  nor _48031_ (_40449_, _40448_, _40447_);
  and _48032_ (_40450_, _40449_, _40403_);
  and _48033_ (_40451_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _48034_ (_40452_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _48035_ (_40453_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _48036_ (_40454_, _40453_, _40452_);
  and _48037_ (_40455_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _48038_ (_40456_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _48039_ (_40457_, _40456_, _40455_);
  and _48040_ (_40458_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _48041_ (_40459_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _48042_ (_40460_, _40459_, _40458_);
  and _48043_ (_40461_, _40460_, _40457_);
  and _48044_ (_40462_, _40461_, _40454_);
  nor _48045_ (_40463_, _40462_, _40213_);
  nor _48046_ (_40464_, _40463_, _40451_);
  not _48047_ (_40465_, _40464_);
  and _48048_ (_40466_, _40465_, _40256_);
  and _48049_ (_40467_, _38806_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _48050_ (_40468_, _40467_, _38900_);
  not _48051_ (_40469_, _40468_);
  and _48052_ (_40470_, _40469_, _40278_);
  nor _48053_ (_40471_, _40470_, _40466_);
  not _48054_ (_40472_, _38334_);
  and _48055_ (_40473_, _40189_, _40472_);
  and _48056_ (_40474_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and _48057_ (_40475_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _48058_ (_40476_, _40475_, _40474_);
  and _48059_ (_40477_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _48060_ (_40478_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _48061_ (_40479_, _40478_, _40477_);
  and _48062_ (_40480_, _40479_, _40476_);
  nor _48063_ (_40481_, _40480_, _40189_);
  nor _48064_ (_40482_, _40481_, _40473_);
  not _48065_ (_40483_, _40482_);
  and _48066_ (_40484_, _40483_, _40235_);
  not _48067_ (_40485_, _40484_);
  not _48068_ (_40486_, _38420_);
  and _48069_ (_40487_, _40486_, _40253_);
  not _48070_ (_40488_, _37932_);
  and _48071_ (_40489_, _40488_, _36788_);
  nor _48072_ (_40490_, _40489_, _40487_);
  and _48073_ (_40491_, _40490_, _40485_);
  and _48074_ (_40492_, _40491_, _40471_);
  not _48075_ (_40493_, _40492_);
  and _48076_ (_40494_, _40493_, _40234_);
  and _48077_ (_40495_, _40165_, _40488_);
  not _48078_ (_40496_, _38402_);
  and _48079_ (_40497_, _40496_, _40253_);
  nor _48080_ (_40498_, _40497_, _40495_);
  and _48081_ (_40499_, _40171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and _48082_ (_40500_, _40173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _48083_ (_40501_, _40500_, _40499_);
  and _48084_ (_40502_, _40168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _48085_ (_40503_, _40190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _48086_ (_40504_, _40503_, _40502_);
  and _48087_ (_40505_, _40504_, _40501_);
  nor _48088_ (_40506_, _40505_, _40189_);
  and _48089_ (_40507_, _40189_, _38356_);
  nor _48090_ (_40508_, _40507_, _40506_);
  not _48091_ (_40509_, _40508_);
  and _48092_ (_40510_, _40509_, _40235_);
  and _48093_ (_40511_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _48094_ (_40512_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _48095_ (_40513_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _48096_ (_40519_, _40513_, _40512_);
  and _48097_ (_40525_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _48098_ (_40531_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _48099_ (_40537_, _40531_, _40525_);
  and _48100_ (_40543_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _48101_ (_40546_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _48102_ (_40547_, _40546_, _40543_);
  and _48103_ (_40548_, _40547_, _40537_);
  and _48104_ (_40549_, _40548_, _40519_);
  nor _48105_ (_40550_, _40549_, _40213_);
  nor _48106_ (_40551_, _40550_, _40511_);
  not _48107_ (_40552_, _40551_);
  and _48108_ (_40553_, _40552_, _40256_);
  nor _48109_ (_40554_, _40553_, _40510_);
  and _48110_ (_40555_, _40278_, _34502_);
  not _48111_ (_40556_, _40555_);
  and _48112_ (_40557_, _40556_, _40554_);
  and _48113_ (_40558_, _40557_, _40498_);
  nor _48114_ (_40559_, _40558_, _40233_);
  nor _48115_ (_40561_, _40559_, _40494_);
  not _48116_ (_40564_, _25105_);
  and _48117_ (_40568_, _40316_, _40564_);
  nor _48118_ (_40571_, _24138_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _48119_ (_40572_, _40571_, _40568_);
  nand _48120_ (_40573_, _40572_, _40561_);
  or _48121_ (_40575_, _40572_, _40561_);
  and _48122_ (_40581_, _40575_, _40573_);
  not _48123_ (_40584_, _40581_);
  not _48124_ (_40585_, _40180_);
  and _48125_ (_40586_, _40399_, _40395_);
  nor _48126_ (_40590_, _40586_, _40585_);
  and _48127_ (_40596_, _40590_, _40584_);
  and _48128_ (_40597_, _40596_, _40450_);
  and _48129_ (_40598_, _40597_, _40401_);
  not _48130_ (_40600_, _40315_);
  and _48131_ (_40606_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not _48132_ (_40609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _48133_ (_40610_, _40395_, _40609_);
  or _48134_ (_40611_, _40610_, _40606_);
  and _48135_ (_40615_, _40611_, _40561_);
  not _48136_ (_40621_, _40561_);
  not _48137_ (_40622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _48138_ (_40623_, _40395_, _40622_);
  and _48139_ (_40626_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _48140_ (_40632_, _40626_, _40623_);
  and _48141_ (_40634_, _40632_, _40621_);
  or _48142_ (_40635_, _40634_, _40615_);
  or _48143_ (_40638_, _40635_, _40600_);
  not _48144_ (_40644_, _40442_);
  and _48145_ (_40646_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not _48146_ (_40647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor _48147_ (_40649_, _40395_, _40647_);
  or _48148_ (_40655_, _40649_, _40646_);
  and _48149_ (_40658_, _40655_, _40561_);
  not _48150_ (_40659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _48151_ (_40660_, _40395_, _40659_);
  and _48152_ (_40664_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _48153_ (_40670_, _40664_, _40660_);
  and _48154_ (_40671_, _40670_, _40621_);
  or _48155_ (_40672_, _40671_, _40658_);
  or _48156_ (_40675_, _40672_, _40315_);
  and _48157_ (_40681_, _40675_, _40644_);
  and _48158_ (_40683_, _40681_, _40638_);
  not _48159_ (_40684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _48160_ (_40687_, _40395_, _40684_);
  or _48161_ (_40693_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _48162_ (_40695_, _40693_, _40687_);
  and _48163_ (_40696_, _40695_, _40561_);
  or _48164_ (_40698_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not _48165_ (_40704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand _48166_ (_40707_, _40395_, _40704_);
  and _48167_ (_40708_, _40707_, _40698_);
  and _48168_ (_40709_, _40708_, _40621_);
  or _48169_ (_40715_, _40709_, _40696_);
  or _48170_ (_40719_, _40715_, _40600_);
  not _48171_ (_40720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _48172_ (_40721_, _40395_, _40720_);
  or _48173_ (_40726_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _48174_ (_40731_, _40726_, _40721_);
  and _48175_ (_40732_, _40731_, _40561_);
  or _48176_ (_40733_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not _48177_ (_40738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand _48178_ (_40743_, _40395_, _40738_);
  and _48179_ (_40744_, _40743_, _40733_);
  and _48180_ (_40745_, _40744_, _40621_);
  or _48181_ (_40750_, _40745_, _40732_);
  or _48182_ (_40754_, _40750_, _40315_);
  and _48183_ (_40755_, _40754_, _40442_);
  and _48184_ (_40756_, _40755_, _40719_);
  or _48185_ (_40757_, _40756_, _40683_);
  or _48186_ (_40758_, _40757_, _40598_);
  not _48187_ (_40759_, _40598_);
  or _48188_ (_40760_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and _48189_ (_40761_, _40760_, _41755_);
  and _48190_ (_42815_, _40761_, _40758_);
  nor _48191_ (_40762_, _40398_, _40585_);
  nor _48192_ (_40763_, _40572_, _40585_);
  and _48193_ (_40764_, _40763_, _40762_);
  and _48194_ (_40765_, _40445_, _40180_);
  nor _48195_ (_40766_, _40319_, _40585_);
  and _48196_ (_40767_, _40766_, _40765_);
  and _48197_ (_40768_, _40767_, _40764_);
  and _48198_ (_40769_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _48199_ (_40770_, _40769_, _25562_);
  nor _48200_ (_40771_, _40770_, _28510_);
  nand _48201_ (_40772_, _25562_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48202_ (_40773_, _17347_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48203_ (_40774_, _40773_, _40772_);
  nor _48204_ (_40775_, _38386_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _48205_ (_40776_, _40775_, _40774_);
  or _48206_ (_40777_, _40776_, _40771_);
  and _48207_ (_40778_, _40777_, _40180_);
  and _48208_ (_40779_, _40778_, _40768_);
  not _48209_ (_40780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _48210_ (_40781_, _40768_, _40780_);
  or _48211_ (_42826_, _40781_, _40779_);
  nor _48212_ (_40782_, _40766_, _40765_);
  nor _48213_ (_40783_, _40763_, _40762_);
  and _48214_ (_40784_, _40783_, _40180_);
  and _48215_ (_40785_, _40784_, _40782_);
  and _48216_ (_40786_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25551_);
  and _48217_ (_40787_, _40786_, _25595_);
  not _48218_ (_40788_, _40787_);
  nor _48219_ (_40789_, _40788_, _28510_);
  not _48220_ (_40790_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48221_ (_40791_, _38364_, _40790_);
  or _48222_ (_40792_, _16186_, _40790_);
  and _48223_ (_40793_, _40792_, _40788_);
  and _48224_ (_40794_, _40793_, _40791_);
  or _48225_ (_40795_, _40794_, _40789_);
  and _48226_ (_40796_, _40795_, _40785_);
  not _48227_ (_40797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _48228_ (_40798_, _40785_, _40797_);
  or _48229_ (_43082_, _40798_, _40796_);
  nand _48230_ (_40799_, _40786_, _25671_);
  nor _48231_ (_40800_, _40799_, _28510_);
  nor _48232_ (_40801_, _38355_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48233_ (_40802_, _40786_, _25627_);
  and _48234_ (_40803_, _40786_, _25562_);
  or _48235_ (_40804_, _40803_, _40769_);
  or _48236_ (_40805_, _40804_, _40802_);
  and _48237_ (_40806_, _40805_, _17173_);
  or _48238_ (_40807_, _40806_, _40801_);
  or _48239_ (_40808_, _40807_, _40800_);
  and _48240_ (_40809_, _40808_, _40785_);
  not _48241_ (_40810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _48242_ (_40811_, _40785_, _40810_);
  or _48243_ (_43088_, _40811_, _40809_);
  not _48244_ (_40812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _48245_ (_40813_, _40785_, _40812_);
  nand _48246_ (_40814_, _40786_, _25638_);
  nor _48247_ (_40815_, _40814_, _28510_);
  nor _48248_ (_40816_, _38348_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48249_ (_40817_, _40786_, _25660_);
  or _48250_ (_40818_, _40817_, _40804_);
  and _48251_ (_40819_, _40818_, _15824_);
  or _48252_ (_40820_, _40819_, _40816_);
  or _48253_ (_40821_, _40820_, _40815_);
  and _48254_ (_40822_, _40821_, _40785_);
  or _48255_ (_43094_, _40822_, _40813_);
  and _48256_ (_40823_, _40803_, _29134_);
  nor _48257_ (_40824_, _38341_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _48258_ (_40825_, _40802_, _40769_);
  or _48259_ (_40826_, _40825_, _40817_);
  and _48260_ (_40827_, _40826_, _16856_);
  or _48261_ (_40828_, _40827_, _40824_);
  or _48262_ (_40829_, _40828_, _40823_);
  and _48263_ (_40830_, _40829_, _40785_);
  not _48264_ (_40831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _48265_ (_40832_, _40785_, _40831_);
  or _48266_ (_43100_, _40832_, _40830_);
  nand _48267_ (_40833_, _40769_, _25595_);
  nor _48268_ (_40834_, _40833_, _28510_);
  nor _48269_ (_40835_, _38334_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48270_ (_40836_, _25595_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48271_ (_40837_, _16022_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48272_ (_40838_, _40837_, _40836_);
  or _48273_ (_40839_, _40838_, _40835_);
  or _48274_ (_40840_, _40839_, _40834_);
  and _48275_ (_40841_, _40840_, _40785_);
  not _48276_ (_40842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _48277_ (_40843_, _40785_, _40842_);
  or _48278_ (_43106_, _40843_, _40841_);
  nand _48279_ (_40844_, _40769_, _25671_);
  nor _48280_ (_40845_, _40844_, _28510_);
  nor _48281_ (_40846_, _38292_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48282_ (_40847_, _25671_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48283_ (_40848_, _17010_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48284_ (_40849_, _40848_, _40847_);
  or _48285_ (_40850_, _40849_, _40846_);
  or _48286_ (_40851_, _40850_, _40845_);
  and _48287_ (_40852_, _40851_, _40785_);
  not _48288_ (_40853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _48289_ (_40854_, _40785_, _40853_);
  or _48290_ (_43112_, _40854_, _40852_);
  nand _48291_ (_40855_, _40769_, _25638_);
  nor _48292_ (_40856_, _40855_, _28510_);
  nor _48293_ (_40857_, _38217_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _48294_ (_40858_, _25638_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _48295_ (_40859_, _16362_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _48296_ (_40860_, _40859_, _40858_);
  or _48297_ (_40861_, _40860_, _40857_);
  or _48298_ (_40862_, _40861_, _40856_);
  and _48299_ (_40863_, _40862_, _40785_);
  not _48300_ (_40864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _48301_ (_40865_, _40785_, _40864_);
  or _48302_ (_43118_, _40865_, _40863_);
  and _48303_ (_40866_, _40785_, _40777_);
  not _48304_ (_40867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _48305_ (_40868_, _40785_, _40867_);
  or _48306_ (_43121_, _40868_, _40866_);
  and _48307_ (_40869_, _40795_, _40180_);
  and _48308_ (_40870_, _40762_, _40572_);
  and _48309_ (_40871_, _40870_, _40782_);
  and _48310_ (_40872_, _40871_, _40869_);
  not _48311_ (_40873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _48312_ (_40874_, _40871_, _40873_);
  or _48313_ (_43129_, _40874_, _40872_);
  and _48314_ (_40875_, _40808_, _40180_);
  and _48315_ (_40876_, _40871_, _40875_);
  not _48316_ (_40877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _48317_ (_40878_, _40871_, _40877_);
  or _48318_ (_43133_, _40878_, _40876_);
  and _48319_ (_40879_, _40821_, _40180_);
  and _48320_ (_40880_, _40871_, _40879_);
  not _48321_ (_40881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _48322_ (_40882_, _40871_, _40881_);
  or _48323_ (_43137_, _40882_, _40880_);
  and _48324_ (_40883_, _40829_, _40180_);
  and _48325_ (_40884_, _40871_, _40883_);
  not _48326_ (_40885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _48327_ (_40886_, _40871_, _40885_);
  or _48328_ (_43141_, _40886_, _40884_);
  and _48329_ (_40887_, _40840_, _40180_);
  and _48330_ (_40888_, _40871_, _40887_);
  not _48331_ (_40889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _48332_ (_40890_, _40871_, _40889_);
  or _48333_ (_43145_, _40890_, _40888_);
  and _48334_ (_40891_, _40851_, _40180_);
  and _48335_ (_40892_, _40871_, _40891_);
  not _48336_ (_40893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _48337_ (_40894_, _40871_, _40893_);
  or _48338_ (_43149_, _40894_, _40892_);
  and _48339_ (_40895_, _40862_, _40180_);
  and _48340_ (_40896_, _40871_, _40895_);
  not _48341_ (_40897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _48342_ (_40898_, _40871_, _40897_);
  or _48343_ (_43153_, _40898_, _40896_);
  and _48344_ (_40899_, _40871_, _40778_);
  nor _48345_ (_40900_, _40871_, _40609_);
  or _48346_ (_43156_, _40900_, _40899_);
  and _48347_ (_40901_, _40763_, _40398_);
  and _48348_ (_40902_, _40901_, _40782_);
  and _48349_ (_40903_, _40902_, _40869_);
  not _48350_ (_40904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _48351_ (_40905_, _40902_, _40904_);
  or _48352_ (_43164_, _40905_, _40903_);
  and _48353_ (_40906_, _40902_, _40875_);
  not _48354_ (_40907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _48355_ (_40908_, _40902_, _40907_);
  or _48356_ (_43168_, _40908_, _40906_);
  and _48357_ (_40909_, _40902_, _40879_);
  not _48358_ (_40910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _48359_ (_40911_, _40902_, _40910_);
  or _48360_ (_43172_, _40911_, _40909_);
  and _48361_ (_40912_, _40902_, _40883_);
  not _48362_ (_40913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _48363_ (_40914_, _40902_, _40913_);
  or _48364_ (_43176_, _40914_, _40912_);
  and _48365_ (_40915_, _40902_, _40887_);
  not _48366_ (_40916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _48367_ (_40917_, _40902_, _40916_);
  or _48368_ (_43180_, _40917_, _40915_);
  and _48369_ (_40918_, _40902_, _40891_);
  not _48370_ (_40919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _48371_ (_40920_, _40902_, _40919_);
  or _48372_ (_43184_, _40920_, _40918_);
  and _48373_ (_40921_, _40902_, _40895_);
  not _48374_ (_40922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _48375_ (_40923_, _40902_, _40922_);
  or _48376_ (_43188_, _40923_, _40921_);
  and _48377_ (_40924_, _40902_, _40778_);
  not _48378_ (_40925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _48379_ (_40926_, _40902_, _40925_);
  or _48380_ (_43191_, _40926_, _40924_);
  and _48381_ (_40927_, _40782_, _40764_);
  and _48382_ (_40928_, _40927_, _40869_);
  not _48383_ (_40929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _48384_ (_40930_, _40927_, _40929_);
  or _48385_ (_43216_, _40930_, _40928_);
  and _48386_ (_40931_, _40927_, _40875_);
  not _48387_ (_40932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _48388_ (_40933_, _40927_, _40932_);
  or _48389_ (_43236_, _40933_, _40931_);
  and _48390_ (_40934_, _40927_, _40879_);
  not _48391_ (_40935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _48392_ (_40936_, _40927_, _40935_);
  or _48393_ (_43254_, _40936_, _40934_);
  and _48394_ (_40937_, _40927_, _40883_);
  not _48395_ (_40938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _48396_ (_40939_, _40927_, _40938_);
  or _48397_ (_43272_, _40939_, _40937_);
  and _48398_ (_40940_, _40927_, _40887_);
  not _48399_ (_40941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _48400_ (_40942_, _40927_, _40941_);
  or _48401_ (_43290_, _40942_, _40940_);
  and _48402_ (_40943_, _40927_, _40891_);
  not _48403_ (_40944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _48404_ (_40945_, _40927_, _40944_);
  or _48405_ (_43309_, _40945_, _40943_);
  and _48406_ (_40946_, _40927_, _40895_);
  not _48407_ (_40947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor _48408_ (_40948_, _40927_, _40947_);
  or _48409_ (_43326_, _40948_, _40946_);
  and _48410_ (_40949_, _40927_, _40778_);
  nor _48411_ (_40950_, _40927_, _40622_);
  or _48412_ (_43344_, _40950_, _40949_);
  and _48413_ (_40951_, _40766_, _40446_);
  and _48414_ (_40952_, _40951_, _40783_);
  and _48415_ (_40953_, _40952_, _40869_);
  not _48416_ (_40954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _48417_ (_40955_, _40952_, _40954_);
  or _48418_ (_43387_, _40955_, _40953_);
  and _48419_ (_40956_, _40952_, _40875_);
  not _48420_ (_40957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _48421_ (_40958_, _40952_, _40957_);
  or _48422_ (_43405_, _40958_, _40956_);
  and _48423_ (_40959_, _40952_, _40879_);
  not _48424_ (_40960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _48425_ (_40961_, _40952_, _40960_);
  or _48426_ (_43423_, _40961_, _40959_);
  and _48427_ (_40962_, _40952_, _40883_);
  not _48428_ (_40963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _48429_ (_40964_, _40952_, _40963_);
  or _48430_ (_43434_, _40964_, _40962_);
  and _48431_ (_40965_, _40952_, _40887_);
  not _48432_ (_40966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _48433_ (_40967_, _40952_, _40966_);
  or _48434_ (_43438_, _40967_, _40965_);
  and _48435_ (_40968_, _40952_, _40891_);
  not _48436_ (_40969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _48437_ (_40970_, _40952_, _40969_);
  or _48438_ (_43442_, _40970_, _40968_);
  and _48439_ (_40971_, _40952_, _40895_);
  not _48440_ (_40972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _48441_ (_40973_, _40952_, _40972_);
  or _48442_ (_43446_, _40973_, _40971_);
  and _48443_ (_40974_, _40952_, _40778_);
  not _48444_ (_40975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _48445_ (_40976_, _40952_, _40975_);
  or _48446_ (_43449_, _40976_, _40974_);
  and _48447_ (_40977_, _40951_, _40870_);
  and _48448_ (_40978_, _40977_, _40869_);
  not _48449_ (_40979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _48450_ (_40980_, _40977_, _40979_);
  or _48451_ (_43454_, _40980_, _40978_);
  and _48452_ (_40981_, _40977_, _40875_);
  not _48453_ (_40982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor _48454_ (_40983_, _40977_, _40982_);
  or _48455_ (_43458_, _40983_, _40981_);
  and _48456_ (_40984_, _40977_, _40879_);
  not _48457_ (_40985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _48458_ (_40986_, _40977_, _40985_);
  or _48459_ (_43462_, _40986_, _40984_);
  and _48460_ (_40987_, _40977_, _40883_);
  not _48461_ (_40988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _48462_ (_40989_, _40977_, _40988_);
  or _48463_ (_43465_, _40989_, _40987_);
  and _48464_ (_40990_, _40977_, _40887_);
  not _48465_ (_40991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _48466_ (_40992_, _40977_, _40991_);
  or _48467_ (_43469_, _40992_, _40990_);
  and _48468_ (_40993_, _40977_, _40891_);
  not _48469_ (_40994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _48470_ (_40995_, _40977_, _40994_);
  or _48471_ (_43473_, _40995_, _40993_);
  and _48472_ (_40996_, _40977_, _40895_);
  not _48473_ (_40997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _48474_ (_40998_, _40977_, _40997_);
  or _48475_ (_43477_, _40998_, _40996_);
  and _48476_ (_40999_, _40977_, _40778_);
  nor _48477_ (_41000_, _40977_, _40647_);
  or _48478_ (_43480_, _41000_, _40999_);
  and _48479_ (_41001_, _40951_, _40901_);
  and _48480_ (_41002_, _41001_, _40869_);
  not _48481_ (_41003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor _48482_ (_41004_, _41001_, _41003_);
  or _48483_ (_43485_, _41004_, _41002_);
  and _48484_ (_41005_, _41001_, _40875_);
  not _48485_ (_41006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _48486_ (_41007_, _41001_, _41006_);
  or _48487_ (_43489_, _41007_, _41005_);
  and _48488_ (_41008_, _41001_, _40879_);
  not _48489_ (_41009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _48490_ (_41010_, _41001_, _41009_);
  or _48491_ (_43493_, _41010_, _41008_);
  and _48492_ (_41011_, _41001_, _40883_);
  not _48493_ (_41012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor _48494_ (_41013_, _41001_, _41012_);
  or _48495_ (_43497_, _41013_, _41011_);
  and _48496_ (_41014_, _41001_, _40887_);
  not _48497_ (_41015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _48498_ (_41016_, _41001_, _41015_);
  or _48499_ (_43501_, _41016_, _41014_);
  and _48500_ (_41017_, _41001_, _40891_);
  not _48501_ (_41018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _48502_ (_41019_, _41001_, _41018_);
  or _48503_ (_43505_, _41019_, _41017_);
  and _48504_ (_41020_, _41001_, _40895_);
  not _48505_ (_41021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _48506_ (_41022_, _41001_, _41021_);
  or _48507_ (_43509_, _41022_, _41020_);
  and _48508_ (_41023_, _41001_, _40778_);
  not _48509_ (_41024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _48510_ (_41025_, _41001_, _41024_);
  or _48511_ (_43512_, _41025_, _41023_);
  and _48512_ (_41026_, _40951_, _40764_);
  and _48513_ (_41027_, _41026_, _40869_);
  not _48514_ (_41028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _48515_ (_41029_, _41026_, _41028_);
  or _48516_ (_43517_, _41029_, _41027_);
  and _48517_ (_41030_, _41026_, _40875_);
  not _48518_ (_41031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _48519_ (_41032_, _41026_, _41031_);
  or _48520_ (_43521_, _41032_, _41030_);
  and _48521_ (_41033_, _41026_, _40879_);
  not _48522_ (_41034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _48523_ (_41035_, _41026_, _41034_);
  or _48524_ (_43525_, _41035_, _41033_);
  and _48525_ (_41036_, _41026_, _40883_);
  not _48526_ (_41037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _48527_ (_41038_, _41026_, _41037_);
  or _48528_ (_43529_, _41038_, _41036_);
  and _48529_ (_41039_, _41026_, _40887_);
  not _48530_ (_41040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor _48531_ (_41041_, _41026_, _41040_);
  or _48532_ (_43533_, _41041_, _41039_);
  and _48533_ (_41042_, _41026_, _40891_);
  not _48534_ (_41043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor _48535_ (_41044_, _41026_, _41043_);
  or _48536_ (_43537_, _41044_, _41042_);
  and _48537_ (_41045_, _41026_, _40895_);
  not _48538_ (_41046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor _48539_ (_41047_, _41026_, _41046_);
  or _48540_ (_43541_, _41047_, _41045_);
  and _48541_ (_41048_, _41026_, _40778_);
  nor _48542_ (_41049_, _41026_, _40659_);
  or _48543_ (_43544_, _41049_, _41048_);
  and _48544_ (_41050_, _40765_, _40319_);
  and _48545_ (_41051_, _41050_, _40783_);
  and _48546_ (_41052_, _41051_, _40869_);
  not _48547_ (_41053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _48548_ (_41054_, _41051_, _41053_);
  or _48549_ (_43552_, _41054_, _41052_);
  and _48550_ (_41055_, _41051_, _40875_);
  not _48551_ (_41056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _48552_ (_41057_, _41051_, _41056_);
  or _48553_ (_43556_, _41057_, _41055_);
  and _48554_ (_41058_, _41051_, _40879_);
  not _48555_ (_41059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _48556_ (_41060_, _41051_, _41059_);
  or _48557_ (_43560_, _41060_, _41058_);
  and _48558_ (_41061_, _41051_, _40883_);
  not _48559_ (_41062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _48560_ (_41063_, _41051_, _41062_);
  or _48561_ (_43564_, _41063_, _41061_);
  and _48562_ (_41064_, _41051_, _40887_);
  not _48563_ (_41065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _48564_ (_41066_, _41051_, _41065_);
  or _48565_ (_43568_, _41066_, _41064_);
  and _48566_ (_41067_, _41051_, _40891_);
  not _48567_ (_41068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _48568_ (_41069_, _41051_, _41068_);
  or _48569_ (_43572_, _41069_, _41067_);
  and _48570_ (_41070_, _41051_, _40895_);
  not _48571_ (_41071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _48572_ (_41072_, _41051_, _41071_);
  or _48573_ (_43576_, _41072_, _41070_);
  and _48574_ (_41073_, _41051_, _40778_);
  nor _48575_ (_41074_, _41051_, _40684_);
  or _48576_ (_43579_, _41074_, _41073_);
  and _48577_ (_41075_, _41050_, _40870_);
  and _48578_ (_41076_, _41075_, _40869_);
  not _48579_ (_41077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _48580_ (_41078_, _41075_, _41077_);
  or _48581_ (_43584_, _41078_, _41076_);
  and _48582_ (_41079_, _41075_, _40875_);
  not _48583_ (_41080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor _48584_ (_41081_, _41075_, _41080_);
  or _48585_ (_43588_, _41081_, _41079_);
  and _48586_ (_41082_, _41075_, _40879_);
  not _48587_ (_41083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _48588_ (_41084_, _41075_, _41083_);
  or _48589_ (_43592_, _41084_, _41082_);
  and _48590_ (_41085_, _41075_, _40883_);
  not _48591_ (_41086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _48592_ (_41087_, _41075_, _41086_);
  or _48593_ (_43596_, _41087_, _41085_);
  and _48594_ (_41088_, _41075_, _40887_);
  not _48595_ (_41089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _48596_ (_41090_, _41075_, _41089_);
  or _48597_ (_43600_, _41090_, _41088_);
  and _48598_ (_41091_, _41075_, _40891_);
  not _48599_ (_41092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _48600_ (_41093_, _41075_, _41092_);
  or _48601_ (_43604_, _41093_, _41091_);
  and _48602_ (_41094_, _41075_, _40895_);
  not _48603_ (_41095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _48604_ (_41096_, _41075_, _41095_);
  or _48605_ (_43608_, _41096_, _41094_);
  and _48606_ (_41097_, _41075_, _40778_);
  not _48607_ (_41098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _48608_ (_41099_, _41075_, _41098_);
  or _48609_ (_43611_, _41099_, _41097_);
  and _48610_ (_41100_, _41050_, _40901_);
  and _48611_ (_41101_, _41100_, _40869_);
  not _48612_ (_41102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _48613_ (_41103_, _41100_, _41102_);
  or _48614_ (_43616_, _41103_, _41101_);
  and _48615_ (_41104_, _41100_, _40875_);
  not _48616_ (_41105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _48617_ (_41106_, _41100_, _41105_);
  or _48618_ (_43620_, _41106_, _41104_);
  and _48619_ (_41107_, _41100_, _40879_);
  not _48620_ (_41108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _48621_ (_41109_, _41100_, _41108_);
  or _48622_ (_43624_, _41109_, _41107_);
  and _48623_ (_41110_, _41100_, _40883_);
  not _48624_ (_41111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _48625_ (_41112_, _41100_, _41111_);
  or _48626_ (_43628_, _41112_, _41110_);
  and _48627_ (_41113_, _41100_, _40887_);
  not _48628_ (_41114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _48629_ (_41115_, _41100_, _41114_);
  or _48630_ (_43632_, _41115_, _41113_);
  and _48631_ (_41116_, _41100_, _40891_);
  not _48632_ (_41117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _48633_ (_41118_, _41100_, _41117_);
  or _48634_ (_43636_, _41118_, _41116_);
  and _48635_ (_41119_, _41100_, _40895_);
  not _48636_ (_41120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _48637_ (_41121_, _41100_, _41120_);
  or _48638_ (_43640_, _41121_, _41119_);
  and _48639_ (_41122_, _41100_, _40778_);
  nor _48640_ (_41123_, _41100_, _40704_);
  or _48641_ (_43643_, _41123_, _41122_);
  and _48642_ (_41124_, _41050_, _40764_);
  and _48643_ (_41125_, _41124_, _40869_);
  not _48644_ (_41126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _48645_ (_41127_, _41124_, _41126_);
  or _48646_ (_43648_, _41127_, _41125_);
  and _48647_ (_41128_, _41124_, _40875_);
  not _48648_ (_41129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _48649_ (_41130_, _41124_, _41129_);
  or _48650_ (_43652_, _41130_, _41128_);
  and _48651_ (_41131_, _41124_, _40879_);
  not _48652_ (_41132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _48653_ (_41133_, _41124_, _41132_);
  or _48654_ (_43656_, _41133_, _41131_);
  and _48655_ (_41134_, _41124_, _40883_);
  not _48656_ (_41135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _48657_ (_41136_, _41124_, _41135_);
  or _48658_ (_43660_, _41136_, _41134_);
  and _48659_ (_41137_, _41124_, _40887_);
  not _48660_ (_41138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _48661_ (_41139_, _41124_, _41138_);
  or _48662_ (_43664_, _41139_, _41137_);
  and _48663_ (_41140_, _41124_, _40891_);
  not _48664_ (_41141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _48665_ (_41142_, _41124_, _41141_);
  or _48666_ (_43668_, _41142_, _41140_);
  and _48667_ (_41143_, _41124_, _40895_);
  not _48668_ (_41144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _48669_ (_41145_, _41124_, _41144_);
  or _48670_ (_43672_, _41145_, _41143_);
  and _48671_ (_41146_, _41124_, _40778_);
  not _48672_ (_41147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _48673_ (_41148_, _41124_, _41147_);
  or _48674_ (_43675_, _41148_, _41146_);
  and _48675_ (_41149_, _40783_, _40767_);
  and _48676_ (_41150_, _41149_, _40869_);
  not _48677_ (_41151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _48678_ (_41152_, _41149_, _41151_);
  or _48679_ (_43681_, _41152_, _41150_);
  and _48680_ (_41153_, _41149_, _40875_);
  not _48681_ (_41154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _48682_ (_41156_, _41149_, _41154_);
  or _48683_ (_43685_, _41156_, _41153_);
  and _48684_ (_41159_, _41149_, _40879_);
  not _48685_ (_41161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _48686_ (_41163_, _41149_, _41161_);
  or _48687_ (_43689_, _41163_, _41159_);
  and _48688_ (_41166_, _41149_, _40883_);
  not _48689_ (_41168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _48690_ (_41170_, _41149_, _41168_);
  or _48691_ (_43693_, _41170_, _41166_);
  and _48692_ (_41173_, _41149_, _40887_);
  not _48693_ (_41175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _48694_ (_41177_, _41149_, _41175_);
  or _48695_ (_43697_, _41177_, _41173_);
  and _48696_ (_41180_, _41149_, _40891_);
  not _48697_ (_41182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _48698_ (_41184_, _41149_, _41182_);
  or _48699_ (_43701_, _41184_, _41180_);
  and _48700_ (_41187_, _41149_, _40895_);
  not _48701_ (_41189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _48702_ (_41191_, _41149_, _41189_);
  or _48703_ (_43705_, _41191_, _41187_);
  and _48704_ (_41194_, _41149_, _40778_);
  nor _48705_ (_41196_, _41149_, _40720_);
  or _48706_ (_43708_, _41196_, _41194_);
  and _48707_ (_41199_, _40870_, _40767_);
  and _48708_ (_41201_, _41199_, _40869_);
  not _48709_ (_41203_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _48710_ (_41204_, _41199_, _41203_);
  or _48711_ (_43713_, _41204_, _41201_);
  and _48712_ (_41205_, _41199_, _40875_);
  not _48713_ (_41206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _48714_ (_41207_, _41199_, _41206_);
  or _48715_ (_43717_, _41207_, _41205_);
  and _48716_ (_41208_, _41199_, _40879_);
  not _48717_ (_41209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _48718_ (_41210_, _41199_, _41209_);
  or _48719_ (_43721_, _41210_, _41208_);
  and _48720_ (_41211_, _41199_, _40883_);
  not _48721_ (_41212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _48722_ (_41213_, _41199_, _41212_);
  or _48723_ (_43725_, _41213_, _41211_);
  and _48724_ (_41214_, _41199_, _40887_);
  not _48725_ (_41215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _48726_ (_41216_, _41199_, _41215_);
  or _48727_ (_43729_, _41216_, _41214_);
  and _48728_ (_41217_, _41199_, _40891_);
  not _48729_ (_41218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor _48730_ (_41219_, _41199_, _41218_);
  or _48731_ (_43733_, _41219_, _41217_);
  and _48732_ (_41220_, _41199_, _40895_);
  not _48733_ (_41221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor _48734_ (_41222_, _41199_, _41221_);
  or _48735_ (_43737_, _41222_, _41220_);
  and _48736_ (_41223_, _41199_, _40778_);
  not _48737_ (_41224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor _48738_ (_41225_, _41199_, _41224_);
  or _48739_ (_43740_, _41225_, _41223_);
  and _48740_ (_41226_, _40901_, _40767_);
  and _48741_ (_41227_, _41226_, _40869_);
  not _48742_ (_41228_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _48743_ (_41229_, _41226_, _41228_);
  or _48744_ (_43745_, _41229_, _41227_);
  and _48745_ (_41230_, _41226_, _40875_);
  not _48746_ (_41231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _48747_ (_41232_, _41226_, _41231_);
  or _48748_ (_43749_, _41232_, _41230_);
  and _48749_ (_41233_, _41226_, _40879_);
  not _48750_ (_41234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _48751_ (_41235_, _41226_, _41234_);
  or _48752_ (_43753_, _41235_, _41233_);
  and _48753_ (_41236_, _41226_, _40883_);
  not _48754_ (_41237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _48755_ (_41238_, _41226_, _41237_);
  or _48756_ (_43757_, _41238_, _41236_);
  and _48757_ (_41239_, _41226_, _40887_);
  not _48758_ (_41240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _48759_ (_41241_, _41226_, _41240_);
  or _48760_ (_43761_, _41241_, _41239_);
  and _48761_ (_41242_, _41226_, _40891_);
  not _48762_ (_41243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _48763_ (_41244_, _41226_, _41243_);
  or _48764_ (_43765_, _41244_, _41242_);
  and _48765_ (_41245_, _41226_, _40895_);
  not _48766_ (_41246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _48767_ (_41247_, _41226_, _41246_);
  or _48768_ (_43767_, _41247_, _41245_);
  and _48769_ (_41248_, _41226_, _40778_);
  nor _48770_ (_41249_, _41226_, _40738_);
  or _48771_ (_43769_, _41249_, _41248_);
  and _48772_ (_41250_, _40869_, _40768_);
  not _48773_ (_41251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _48774_ (_41252_, _40768_, _41251_);
  or _48775_ (_43774_, _41252_, _41250_);
  and _48776_ (_41253_, _40875_, _40768_);
  not _48777_ (_41254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _48778_ (_41255_, _40768_, _41254_);
  or _48779_ (_43778_, _41255_, _41253_);
  and _48780_ (_41256_, _40879_, _40768_);
  not _48781_ (_41257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _48782_ (_41258_, _40768_, _41257_);
  or _48783_ (_43782_, _41258_, _41256_);
  and _48784_ (_41259_, _40883_, _40768_);
  not _48785_ (_41260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _48786_ (_41261_, _40768_, _41260_);
  or _48787_ (_43785_, _41261_, _41259_);
  and _48788_ (_41262_, _40887_, _40768_);
  not _48789_ (_41263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor _48790_ (_41264_, _40768_, _41263_);
  or _48791_ (_43788_, _41264_, _41262_);
  and _48792_ (_41265_, _40891_, _40768_);
  not _48793_ (_41266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _48794_ (_41267_, _40768_, _41266_);
  or _48795_ (_43792_, _41267_, _41265_);
  and _48796_ (_41268_, _40895_, _40768_);
  not _48797_ (_41269_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor _48798_ (_41270_, _40768_, _41269_);
  or _48799_ (_43796_, _41270_, _41268_);
  and _48800_ (_41271_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _48801_ (_41272_, _40395_, _40873_);
  or _48802_ (_41273_, _41272_, _41271_);
  and _48803_ (_41274_, _41273_, _40561_);
  nor _48804_ (_41275_, _40395_, _40929_);
  and _48805_ (_41276_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _48806_ (_41277_, _41276_, _41275_);
  and _48807_ (_41278_, _41277_, _40621_);
  or _48808_ (_41279_, _41278_, _41274_);
  or _48809_ (_41280_, _41279_, _40600_);
  and _48810_ (_41281_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _48811_ (_41282_, _40395_, _40979_);
  or _48812_ (_41283_, _41282_, _41281_);
  and _48813_ (_41284_, _41283_, _40561_);
  nor _48814_ (_41285_, _40395_, _41028_);
  and _48815_ (_41286_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _48816_ (_41287_, _41286_, _41285_);
  and _48817_ (_41288_, _41287_, _40621_);
  or _48818_ (_41289_, _41288_, _41284_);
  or _48819_ (_41290_, _41289_, _40315_);
  and _48820_ (_41291_, _41290_, _40644_);
  and _48821_ (_41292_, _41291_, _41280_);
  nand _48822_ (_41293_, _40395_, _41053_);
  or _48823_ (_41294_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _48824_ (_41295_, _41294_, _41293_);
  and _48825_ (_41296_, _41295_, _40561_);
  or _48826_ (_41297_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand _48827_ (_41298_, _40395_, _41102_);
  and _48828_ (_41299_, _41298_, _41297_);
  and _48829_ (_41300_, _41299_, _40621_);
  or _48830_ (_41301_, _41300_, _41296_);
  or _48831_ (_41302_, _41301_, _40600_);
  nand _48832_ (_41303_, _40395_, _41151_);
  or _48833_ (_41304_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _48834_ (_41305_, _41304_, _41303_);
  and _48835_ (_41306_, _41305_, _40561_);
  or _48836_ (_41307_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand _48837_ (_41308_, _40395_, _41228_);
  and _48838_ (_41309_, _41308_, _41307_);
  and _48839_ (_41310_, _41309_, _40621_);
  or _48840_ (_41311_, _41310_, _41306_);
  or _48841_ (_41312_, _41311_, _40315_);
  and _48842_ (_41313_, _41312_, _40442_);
  and _48843_ (_41314_, _41313_, _41302_);
  or _48844_ (_41315_, _41314_, _41292_);
  or _48845_ (_41316_, _41315_, _40598_);
  or _48846_ (_41317_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _48847_ (_41318_, _41317_, _41755_);
  and _48848_ (_01407_, _41318_, _41316_);
  and _48849_ (_41319_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _48850_ (_41320_, _40395_, _40877_);
  or _48851_ (_41321_, _41320_, _41319_);
  and _48852_ (_41322_, _41321_, _40561_);
  nor _48853_ (_41323_, _40395_, _40932_);
  and _48854_ (_41324_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _48855_ (_41325_, _41324_, _41323_);
  and _48856_ (_41326_, _41325_, _40621_);
  or _48857_ (_41327_, _41326_, _41322_);
  or _48858_ (_41328_, _41327_, _40600_);
  and _48859_ (_41329_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _48860_ (_41330_, _40395_, _40982_);
  or _48861_ (_41331_, _41330_, _41329_);
  and _48862_ (_41332_, _41331_, _40561_);
  nor _48863_ (_41333_, _40395_, _41031_);
  and _48864_ (_41334_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _48865_ (_41335_, _41334_, _41333_);
  and _48866_ (_41336_, _41335_, _40621_);
  or _48867_ (_41337_, _41336_, _41332_);
  or _48868_ (_41338_, _41337_, _40315_);
  and _48869_ (_41339_, _41338_, _40644_);
  and _48870_ (_41340_, _41339_, _41328_);
  nand _48871_ (_41341_, _40395_, _41056_);
  or _48872_ (_41342_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _48873_ (_41343_, _41342_, _41341_);
  and _48874_ (_41344_, _41343_, _40561_);
  or _48875_ (_41345_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand _48876_ (_41346_, _40395_, _41105_);
  and _48877_ (_41347_, _41346_, _41345_);
  and _48878_ (_41348_, _41347_, _40621_);
  or _48879_ (_41349_, _41348_, _41344_);
  or _48880_ (_41350_, _41349_, _40600_);
  nand _48881_ (_41351_, _40395_, _41154_);
  or _48882_ (_41352_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _48883_ (_41353_, _41352_, _41351_);
  and _48884_ (_41354_, _41353_, _40561_);
  or _48885_ (_41355_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand _48886_ (_41356_, _40395_, _41231_);
  and _48887_ (_41357_, _41356_, _41355_);
  and _48888_ (_41358_, _41357_, _40621_);
  or _48889_ (_41359_, _41358_, _41354_);
  or _48890_ (_41360_, _41359_, _40315_);
  and _48891_ (_41361_, _41360_, _40442_);
  and _48892_ (_41362_, _41361_, _41350_);
  or _48893_ (_41363_, _41362_, _41340_);
  or _48894_ (_41364_, _41363_, _40598_);
  or _48895_ (_41365_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and _48896_ (_41366_, _41365_, _41755_);
  and _48897_ (_01409_, _41366_, _41364_);
  and _48898_ (_41367_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _48899_ (_41368_, _40395_, _40881_);
  or _48900_ (_41369_, _41368_, _41367_);
  and _48901_ (_41370_, _41369_, _40561_);
  nor _48902_ (_41371_, _40395_, _40935_);
  and _48903_ (_41372_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _48904_ (_41373_, _41372_, _41371_);
  and _48905_ (_41374_, _41373_, _40621_);
  or _48906_ (_41375_, _41374_, _41370_);
  or _48907_ (_41376_, _41375_, _40600_);
  and _48908_ (_41377_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _48909_ (_41378_, _40395_, _40985_);
  or _48910_ (_41379_, _41378_, _41377_);
  and _48911_ (_41380_, _41379_, _40561_);
  nor _48912_ (_41381_, _40395_, _41034_);
  and _48913_ (_41382_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _48914_ (_41383_, _41382_, _41381_);
  and _48915_ (_41384_, _41383_, _40621_);
  or _48916_ (_41385_, _41384_, _41380_);
  or _48917_ (_41386_, _41385_, _40315_);
  and _48918_ (_41387_, _41386_, _40644_);
  and _48919_ (_41388_, _41387_, _41376_);
  nand _48920_ (_41389_, _40395_, _41059_);
  or _48921_ (_41390_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _48922_ (_41391_, _41390_, _41389_);
  and _48923_ (_41392_, _41391_, _40561_);
  or _48924_ (_41393_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand _48925_ (_41394_, _40395_, _41108_);
  and _48926_ (_41395_, _41394_, _41393_);
  and _48927_ (_41396_, _41395_, _40621_);
  or _48928_ (_41397_, _41396_, _41392_);
  or _48929_ (_41398_, _41397_, _40600_);
  nand _48930_ (_41399_, _40395_, _41161_);
  or _48931_ (_41400_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _48932_ (_41401_, _41400_, _41399_);
  and _48933_ (_41402_, _41401_, _40561_);
  or _48934_ (_41403_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand _48935_ (_41404_, _40395_, _41234_);
  and _48936_ (_41405_, _41404_, _41403_);
  and _48937_ (_41406_, _41405_, _40621_);
  or _48938_ (_41407_, _41406_, _41402_);
  or _48939_ (_41408_, _41407_, _40315_);
  and _48940_ (_41409_, _41408_, _40442_);
  and _48941_ (_41410_, _41409_, _41398_);
  or _48942_ (_41411_, _41410_, _41388_);
  or _48943_ (_41412_, _41411_, _40598_);
  or _48944_ (_41413_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _48945_ (_41414_, _41413_, _41755_);
  and _48946_ (_01411_, _41414_, _41412_);
  and _48947_ (_41415_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _48948_ (_41416_, _40395_, _40885_);
  or _48949_ (_41417_, _41416_, _41415_);
  and _48950_ (_41418_, _41417_, _40561_);
  nor _48951_ (_41419_, _40395_, _40938_);
  and _48952_ (_41420_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _48953_ (_41421_, _41420_, _41419_);
  and _48954_ (_41422_, _41421_, _40621_);
  or _48955_ (_41423_, _41422_, _41418_);
  or _48956_ (_41424_, _41423_, _40600_);
  and _48957_ (_41425_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _48958_ (_41426_, _40395_, _40988_);
  or _48959_ (_41427_, _41426_, _41425_);
  and _48960_ (_41428_, _41427_, _40561_);
  nor _48961_ (_41429_, _40395_, _41037_);
  and _48962_ (_41430_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _48963_ (_41431_, _41430_, _41429_);
  and _48964_ (_41432_, _41431_, _40621_);
  or _48965_ (_41433_, _41432_, _41428_);
  or _48966_ (_41434_, _41433_, _40315_);
  and _48967_ (_41435_, _41434_, _40644_);
  and _48968_ (_41436_, _41435_, _41424_);
  nand _48969_ (_41437_, _40395_, _41062_);
  or _48970_ (_41438_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _48971_ (_41439_, _41438_, _41437_);
  and _48972_ (_41440_, _41439_, _40561_);
  or _48973_ (_41441_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand _48974_ (_41442_, _40395_, _41111_);
  and _48975_ (_41443_, _41442_, _41441_);
  and _48976_ (_41444_, _41443_, _40621_);
  or _48977_ (_41445_, _41444_, _41440_);
  or _48978_ (_41446_, _41445_, _40600_);
  nand _48979_ (_41447_, _40395_, _41168_);
  or _48980_ (_41448_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _48981_ (_41449_, _41448_, _41447_);
  and _48982_ (_41450_, _41449_, _40561_);
  or _48983_ (_41451_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand _48984_ (_41452_, _40395_, _41237_);
  and _48985_ (_41453_, _41452_, _41451_);
  and _48986_ (_41454_, _41453_, _40621_);
  or _48987_ (_41455_, _41454_, _41450_);
  or _48988_ (_41456_, _41455_, _40315_);
  and _48989_ (_41457_, _41456_, _40442_);
  and _48990_ (_41458_, _41457_, _41446_);
  or _48991_ (_41459_, _41458_, _41436_);
  or _48992_ (_41460_, _41459_, _40598_);
  or _48993_ (_41461_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and _48994_ (_41462_, _41461_, _41755_);
  and _48995_ (_01413_, _41462_, _41460_);
  and _48996_ (_41463_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _48997_ (_41464_, _40395_, _40889_);
  or _48998_ (_41465_, _41464_, _41463_);
  and _48999_ (_41466_, _41465_, _40561_);
  nor _49000_ (_41467_, _40395_, _40941_);
  and _49001_ (_41468_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _49002_ (_41469_, _41468_, _41467_);
  and _49003_ (_41470_, _41469_, _40621_);
  or _49004_ (_41471_, _41470_, _41466_);
  or _49005_ (_41472_, _41471_, _40600_);
  and _49006_ (_41473_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _49007_ (_41474_, _40395_, _40991_);
  or _49008_ (_41475_, _41474_, _41473_);
  and _49009_ (_41476_, _41475_, _40561_);
  nor _49010_ (_41477_, _40395_, _41040_);
  and _49011_ (_41478_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _49012_ (_41479_, _41478_, _41477_);
  and _49013_ (_41480_, _41479_, _40621_);
  or _49014_ (_41481_, _41480_, _41476_);
  or _49015_ (_41482_, _41481_, _40315_);
  and _49016_ (_41483_, _41482_, _40644_);
  and _49017_ (_41484_, _41483_, _41472_);
  nand _49018_ (_41485_, _40395_, _41065_);
  or _49019_ (_41486_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _49020_ (_41487_, _41486_, _41485_);
  and _49021_ (_41488_, _41487_, _40561_);
  or _49022_ (_41489_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand _49023_ (_41490_, _40395_, _41114_);
  and _49024_ (_41491_, _41490_, _41489_);
  and _49025_ (_41492_, _41491_, _40621_);
  or _49026_ (_41493_, _41492_, _41488_);
  or _49027_ (_41494_, _41493_, _40600_);
  nand _49028_ (_41495_, _40395_, _41175_);
  or _49029_ (_41496_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and _49030_ (_41497_, _41496_, _41495_);
  and _49031_ (_41498_, _41497_, _40561_);
  or _49032_ (_41499_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand _49033_ (_41500_, _40395_, _41240_);
  and _49034_ (_41501_, _41500_, _41499_);
  and _49035_ (_41502_, _41501_, _40621_);
  or _49036_ (_41503_, _41502_, _41498_);
  or _49037_ (_41504_, _41503_, _40315_);
  and _49038_ (_41505_, _41504_, _40442_);
  and _49039_ (_41506_, _41505_, _41494_);
  or _49040_ (_41507_, _41506_, _41484_);
  or _49041_ (_41508_, _41507_, _40598_);
  or _49042_ (_41509_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and _49043_ (_41510_, _41509_, _41755_);
  and _49044_ (_01415_, _41510_, _41508_);
  and _49045_ (_41511_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _49046_ (_41512_, _40395_, _40893_);
  or _49047_ (_41513_, _41512_, _41511_);
  and _49048_ (_41514_, _41513_, _40561_);
  nor _49049_ (_41515_, _40395_, _40944_);
  and _49050_ (_41516_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _49051_ (_41517_, _41516_, _41515_);
  and _49052_ (_41518_, _41517_, _40621_);
  or _49053_ (_41519_, _41518_, _41514_);
  or _49054_ (_41520_, _41519_, _40600_);
  and _49055_ (_41521_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _49056_ (_41522_, _40395_, _40994_);
  or _49057_ (_41523_, _41522_, _41521_);
  and _49058_ (_41524_, _41523_, _40561_);
  nor _49059_ (_41525_, _40395_, _41043_);
  and _49060_ (_41526_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _49061_ (_41527_, _41526_, _41525_);
  and _49062_ (_41528_, _41527_, _40621_);
  or _49063_ (_41529_, _41528_, _41524_);
  or _49064_ (_41530_, _41529_, _40315_);
  and _49065_ (_41531_, _41530_, _40644_);
  and _49066_ (_41532_, _41531_, _41520_);
  nand _49067_ (_41533_, _40395_, _41068_);
  or _49068_ (_41534_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _49069_ (_41535_, _41534_, _41533_);
  and _49070_ (_41536_, _41535_, _40561_);
  or _49071_ (_41537_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _49072_ (_41538_, _40395_, _41117_);
  and _49073_ (_41539_, _41538_, _41537_);
  and _49074_ (_41540_, _41539_, _40621_);
  or _49075_ (_41541_, _41540_, _41536_);
  or _49076_ (_41542_, _41541_, _40600_);
  nand _49077_ (_41543_, _40395_, _41182_);
  or _49078_ (_41544_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _49079_ (_41545_, _41544_, _41543_);
  and _49080_ (_41546_, _41545_, _40561_);
  or _49081_ (_41547_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _49082_ (_41548_, _40395_, _41243_);
  and _49083_ (_41549_, _41548_, _41547_);
  and _49084_ (_41550_, _41549_, _40621_);
  or _49085_ (_41551_, _41550_, _41546_);
  or _49086_ (_41552_, _41551_, _40315_);
  and _49087_ (_41553_, _41552_, _40442_);
  and _49088_ (_41554_, _41553_, _41542_);
  or _49089_ (_41555_, _41554_, _41532_);
  or _49090_ (_41556_, _41555_, _40598_);
  or _49091_ (_41557_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _49092_ (_41558_, _41557_, _41755_);
  and _49093_ (_01416_, _41558_, _41556_);
  and _49094_ (_41559_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _49095_ (_41560_, _40395_, _40897_);
  or _49096_ (_41561_, _41560_, _41559_);
  and _49097_ (_41562_, _41561_, _40561_);
  nor _49098_ (_41563_, _40395_, _40947_);
  and _49099_ (_41564_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _49100_ (_41565_, _41564_, _41563_);
  and _49101_ (_41566_, _41565_, _40621_);
  or _49102_ (_41567_, _41566_, _41562_);
  or _49103_ (_41568_, _41567_, _40600_);
  and _49104_ (_41569_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _49105_ (_41570_, _40395_, _40997_);
  or _49106_ (_41571_, _41570_, _41569_);
  and _49107_ (_41572_, _41571_, _40561_);
  nor _49108_ (_41573_, _40395_, _41046_);
  and _49109_ (_41574_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _49110_ (_41575_, _41574_, _41573_);
  and _49111_ (_41576_, _41575_, _40621_);
  or _49112_ (_41577_, _41576_, _41572_);
  or _49113_ (_41578_, _41577_, _40315_);
  and _49114_ (_41579_, _41578_, _40644_);
  and _49115_ (_41580_, _41579_, _41568_);
  nand _49116_ (_41581_, _40395_, _41071_);
  or _49117_ (_41582_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _49118_ (_41583_, _41582_, _41581_);
  and _49119_ (_41584_, _41583_, _40561_);
  or _49120_ (_41585_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand _49121_ (_41586_, _40395_, _41120_);
  and _49122_ (_41587_, _41586_, _41585_);
  and _49123_ (_41588_, _41587_, _40621_);
  or _49124_ (_41589_, _41588_, _41584_);
  or _49125_ (_41590_, _41589_, _40600_);
  nand _49126_ (_41591_, _40395_, _41189_);
  or _49127_ (_41592_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _49128_ (_41593_, _41592_, _41591_);
  and _49129_ (_41594_, _41593_, _40561_);
  or _49130_ (_41595_, _40395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand _49131_ (_41596_, _40395_, _41246_);
  and _49132_ (_41597_, _41596_, _41595_);
  and _49133_ (_41598_, _41597_, _40621_);
  or _49134_ (_41599_, _41598_, _41594_);
  or _49135_ (_41600_, _41599_, _40315_);
  and _49136_ (_41601_, _41600_, _40442_);
  and _49137_ (_41602_, _41601_, _41590_);
  or _49138_ (_41603_, _41602_, _41580_);
  or _49139_ (_41604_, _41603_, _40598_);
  or _49140_ (_41605_, _40759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _49141_ (_41606_, _41605_, _41755_);
  and _49142_ (_01418_, _41606_, _41604_);
  or _49143_ (_41607_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not _49144_ (_41608_, \oc8051_gm_cxrom_1.cell0.valid );
  or _49145_ (_41609_, _41608_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand _49146_ (_41610_, _41609_, _41607_);
  nand _49147_ (_41611_, _41610_, _41755_);
  or _49148_ (_41612_, \oc8051_gm_cxrom_1.cell0.data [7], _41755_);
  and _49149_ (_01426_, _41612_, _41611_);
  or _49150_ (_41613_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or _49151_ (_41614_, \oc8051_gm_cxrom_1.cell0.data [0], _41608_);
  nand _49152_ (_41615_, _41614_, _41613_);
  nand _49153_ (_41616_, _41615_, _41755_);
  or _49154_ (_41617_, \oc8051_gm_cxrom_1.cell0.data [0], _41755_);
  and _49155_ (_01433_, _41617_, _41616_);
  or _49156_ (_41618_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or _49157_ (_41619_, \oc8051_gm_cxrom_1.cell0.data [1], _41608_);
  nand _49158_ (_41620_, _41619_, _41618_);
  nand _49159_ (_41621_, _41620_, _41755_);
  or _49160_ (_41622_, \oc8051_gm_cxrom_1.cell0.data [1], _41755_);
  and _49161_ (_01437_, _41622_, _41621_);
  or _49162_ (_41623_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or _49163_ (_41624_, \oc8051_gm_cxrom_1.cell0.data [2], _41608_);
  nand _49164_ (_41625_, _41624_, _41623_);
  nand _49165_ (_41626_, _41625_, _41755_);
  or _49166_ (_41627_, \oc8051_gm_cxrom_1.cell0.data [2], _41755_);
  and _49167_ (_01441_, _41627_, _41626_);
  or _49168_ (_41628_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or _49169_ (_41629_, \oc8051_gm_cxrom_1.cell0.data [3], _41608_);
  nand _49170_ (_41630_, _41629_, _41628_);
  nand _49171_ (_41631_, _41630_, _41755_);
  or _49172_ (_41632_, \oc8051_gm_cxrom_1.cell0.data [3], _41755_);
  and _49173_ (_01445_, _41632_, _41631_);
  or _49174_ (_41633_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or _49175_ (_41634_, \oc8051_gm_cxrom_1.cell0.data [4], _41608_);
  nand _49176_ (_41635_, _41634_, _41633_);
  nand _49177_ (_41636_, _41635_, _41755_);
  or _49178_ (_41637_, \oc8051_gm_cxrom_1.cell0.data [4], _41755_);
  and _49179_ (_01449_, _41637_, _41636_);
  or _49180_ (_41638_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or _49181_ (_41639_, \oc8051_gm_cxrom_1.cell0.data [5], _41608_);
  nand _49182_ (_41640_, _41639_, _41638_);
  nand _49183_ (_41641_, _41640_, _41755_);
  or _49184_ (_41642_, \oc8051_gm_cxrom_1.cell0.data [5], _41755_);
  and _49185_ (_01453_, _41642_, _41641_);
  or _49186_ (_41643_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or _49187_ (_41644_, \oc8051_gm_cxrom_1.cell0.data [6], _41608_);
  nand _49188_ (_41645_, _41644_, _41643_);
  nand _49189_ (_41646_, _41645_, _41755_);
  or _49190_ (_41647_, \oc8051_gm_cxrom_1.cell0.data [6], _41755_);
  and _49191_ (_01457_, _41647_, _41646_);
  or _49192_ (_41648_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not _49193_ (_41649_, \oc8051_gm_cxrom_1.cell1.valid );
  or _49194_ (_41650_, _41649_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand _49195_ (_41651_, _41650_, _41648_);
  nand _49196_ (_41652_, _41651_, _41755_);
  or _49197_ (_41653_, \oc8051_gm_cxrom_1.cell1.data [7], _41755_);
  and _49198_ (_01478_, _41653_, _41652_);
  or _49199_ (_41654_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or _49200_ (_41655_, \oc8051_gm_cxrom_1.cell1.data [0], _41649_);
  nand _49201_ (_41656_, _41655_, _41654_);
  nand _49202_ (_41657_, _41656_, _41755_);
  or _49203_ (_41658_, \oc8051_gm_cxrom_1.cell1.data [0], _41755_);
  and _49204_ (_01485_, _41658_, _41657_);
  or _49205_ (_41659_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or _49206_ (_41660_, \oc8051_gm_cxrom_1.cell1.data [1], _41649_);
  nand _49207_ (_41661_, _41660_, _41659_);
  nand _49208_ (_41662_, _41661_, _41755_);
  or _49209_ (_41663_, \oc8051_gm_cxrom_1.cell1.data [1], _41755_);
  and _49210_ (_01489_, _41663_, _41662_);
  or _49211_ (_41664_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or _49212_ (_41665_, \oc8051_gm_cxrom_1.cell1.data [2], _41649_);
  nand _49213_ (_41666_, _41665_, _41664_);
  nand _49214_ (_41667_, _41666_, _41755_);
  or _49215_ (_41668_, \oc8051_gm_cxrom_1.cell1.data [2], _41755_);
  and _49216_ (_01493_, _41668_, _41667_);
  or _49217_ (_41669_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or _49218_ (_41670_, \oc8051_gm_cxrom_1.cell1.data [3], _41649_);
  nand _49219_ (_41671_, _41670_, _41669_);
  nand _49220_ (_41672_, _41671_, _41755_);
  or _49221_ (_41673_, \oc8051_gm_cxrom_1.cell1.data [3], _41755_);
  and _49222_ (_01496_, _41673_, _41672_);
  or _49223_ (_41674_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or _49224_ (_41675_, \oc8051_gm_cxrom_1.cell1.data [4], _41649_);
  nand _49225_ (_41676_, _41675_, _41674_);
  nand _49226_ (_41677_, _41676_, _41755_);
  or _49227_ (_41678_, \oc8051_gm_cxrom_1.cell1.data [4], _41755_);
  and _49228_ (_01500_, _41678_, _41677_);
  or _49229_ (_41679_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or _49230_ (_41680_, \oc8051_gm_cxrom_1.cell1.data [5], _41649_);
  nand _49231_ (_41681_, _41680_, _41679_);
  nand _49232_ (_41682_, _41681_, _41755_);
  or _49233_ (_41683_, \oc8051_gm_cxrom_1.cell1.data [5], _41755_);
  and _49234_ (_01504_, _41683_, _41682_);
  or _49235_ (_41684_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or _49236_ (_41685_, \oc8051_gm_cxrom_1.cell1.data [6], _41649_);
  nand _49237_ (_41686_, _41685_, _41684_);
  nand _49238_ (_41687_, _41686_, _41755_);
  or _49239_ (_41688_, \oc8051_gm_cxrom_1.cell1.data [6], _41755_);
  and _49240_ (_01508_, _41688_, _41687_);
  or _49241_ (_41689_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not _49242_ (_41690_, \oc8051_gm_cxrom_1.cell2.valid );
  or _49243_ (_41691_, _41690_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand _49244_ (_41692_, _41691_, _41689_);
  nand _49245_ (_41693_, _41692_, _41755_);
  or _49246_ (_41694_, \oc8051_gm_cxrom_1.cell2.data [7], _41755_);
  and _49247_ (_01529_, _41694_, _41693_);
  or _49248_ (_41695_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or _49249_ (_41696_, \oc8051_gm_cxrom_1.cell2.data [0], _41690_);
  nand _49250_ (_41697_, _41696_, _41695_);
  nand _49251_ (_41699_, _41697_, _41755_);
  or _49252_ (_41700_, \oc8051_gm_cxrom_1.cell2.data [0], _41755_);
  and _49253_ (_01536_, _41700_, _41699_);
  or _49254_ (_41703_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or _49255_ (_41704_, \oc8051_gm_cxrom_1.cell2.data [1], _41690_);
  nand _49256_ (_41706_, _41704_, _41703_);
  nand _49257_ (_41708_, _41706_, _41755_);
  or _49258_ (_41710_, \oc8051_gm_cxrom_1.cell2.data [1], _41755_);
  and _49259_ (_01540_, _41710_, _41708_);
  or _49260_ (_41712_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or _49261_ (_41713_, \oc8051_gm_cxrom_1.cell2.data [2], _41690_);
  nand _49262_ (_41714_, _41713_, _41712_);
  nand _49263_ (_41715_, _41714_, _41755_);
  or _49264_ (_41716_, \oc8051_gm_cxrom_1.cell2.data [2], _41755_);
  and _49265_ (_01544_, _41716_, _41715_);
  or _49266_ (_41717_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or _49267_ (_41718_, \oc8051_gm_cxrom_1.cell2.data [3], _41690_);
  nand _49268_ (_41719_, _41718_, _41717_);
  nand _49269_ (_41720_, _41719_, _41755_);
  or _49270_ (_41721_, \oc8051_gm_cxrom_1.cell2.data [3], _41755_);
  and _49271_ (_01548_, _41721_, _41720_);
  or _49272_ (_41722_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or _49273_ (_41723_, \oc8051_gm_cxrom_1.cell2.data [4], _41690_);
  nand _49274_ (_41724_, _41723_, _41722_);
  nand _49275_ (_41725_, _41724_, _41755_);
  or _49276_ (_41726_, \oc8051_gm_cxrom_1.cell2.data [4], _41755_);
  and _49277_ (_01552_, _41726_, _41725_);
  or _49278_ (_41727_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or _49279_ (_41728_, \oc8051_gm_cxrom_1.cell2.data [5], _41690_);
  nand _49280_ (_41729_, _41728_, _41727_);
  nand _49281_ (_41730_, _41729_, _41755_);
  or _49282_ (_41731_, \oc8051_gm_cxrom_1.cell2.data [5], _41755_);
  and _49283_ (_01556_, _41731_, _41730_);
  or _49284_ (_41732_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or _49285_ (_41733_, \oc8051_gm_cxrom_1.cell2.data [6], _41690_);
  nand _49286_ (_41734_, _41733_, _41732_);
  nand _49287_ (_41735_, _41734_, _41755_);
  or _49288_ (_41736_, \oc8051_gm_cxrom_1.cell2.data [6], _41755_);
  and _49289_ (_01560_, _41736_, _41735_);
  or _49290_ (_41737_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not _49291_ (_41738_, \oc8051_gm_cxrom_1.cell3.valid );
  or _49292_ (_41739_, _41738_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand _49293_ (_41740_, _41739_, _41737_);
  nand _49294_ (_41741_, _41740_, _41755_);
  or _49295_ (_41742_, \oc8051_gm_cxrom_1.cell3.data [7], _41755_);
  and _49296_ (_01581_, _41742_, _41741_);
  or _49297_ (_41745_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or _49298_ (_41747_, \oc8051_gm_cxrom_1.cell3.data [0], _41738_);
  nand _49299_ (_41749_, _41747_, _41745_);
  nand _49300_ (_41751_, _41749_, _41755_);
  or _49301_ (_41753_, \oc8051_gm_cxrom_1.cell3.data [0], _41755_);
  and _49302_ (_01588_, _41753_, _41751_);
  or _49303_ (_41756_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or _49304_ (_41757_, \oc8051_gm_cxrom_1.cell3.data [1], _41738_);
  nand _49305_ (_41758_, _41757_, _41756_);
  nand _49306_ (_41759_, _41758_, _41755_);
  or _49307_ (_41760_, \oc8051_gm_cxrom_1.cell3.data [1], _41755_);
  and _49308_ (_01592_, _41760_, _41759_);
  or _49309_ (_41761_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or _49310_ (_41762_, \oc8051_gm_cxrom_1.cell3.data [2], _41738_);
  nand _49311_ (_41763_, _41762_, _41761_);
  nand _49312_ (_41764_, _41763_, _41755_);
  or _49313_ (_41765_, \oc8051_gm_cxrom_1.cell3.data [2], _41755_);
  and _49314_ (_01596_, _41765_, _41764_);
  or _49315_ (_41766_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or _49316_ (_41767_, \oc8051_gm_cxrom_1.cell3.data [3], _41738_);
  nand _49317_ (_41768_, _41767_, _41766_);
  nand _49318_ (_41769_, _41768_, _41755_);
  or _49319_ (_41770_, \oc8051_gm_cxrom_1.cell3.data [3], _41755_);
  and _49320_ (_01600_, _41770_, _41769_);
  or _49321_ (_41771_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or _49322_ (_41772_, \oc8051_gm_cxrom_1.cell3.data [4], _41738_);
  nand _49323_ (_41773_, _41772_, _41771_);
  nand _49324_ (_41774_, _41773_, _41755_);
  or _49325_ (_41775_, \oc8051_gm_cxrom_1.cell3.data [4], _41755_);
  and _49326_ (_01604_, _41775_, _41774_);
  or _49327_ (_41776_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or _49328_ (_41777_, \oc8051_gm_cxrom_1.cell3.data [5], _41738_);
  nand _49329_ (_41778_, _41777_, _41776_);
  nand _49330_ (_41779_, _41778_, _41755_);
  or _49331_ (_41780_, \oc8051_gm_cxrom_1.cell3.data [5], _41755_);
  and _49332_ (_01607_, _41780_, _41779_);
  or _49333_ (_41781_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or _49334_ (_41782_, \oc8051_gm_cxrom_1.cell3.data [6], _41738_);
  nand _49335_ (_41783_, _41782_, _41781_);
  nand _49336_ (_41784_, _41783_, _41755_);
  or _49337_ (_41785_, \oc8051_gm_cxrom_1.cell3.data [6], _41755_);
  and _49338_ (_01608_, _41785_, _41784_);
  or _49339_ (_41786_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not _49340_ (_41787_, \oc8051_gm_cxrom_1.cell4.valid );
  or _49341_ (_41788_, _41787_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand _49342_ (_41789_, _41788_, _41786_);
  nand _49343_ (_41790_, _41789_, _41755_);
  or _49344_ (_41791_, \oc8051_gm_cxrom_1.cell4.data [7], _41755_);
  and _49345_ (_01620_, _41791_, _41790_);
  or _49346_ (_41792_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or _49347_ (_41793_, \oc8051_gm_cxrom_1.cell4.data [0], _41787_);
  nand _49348_ (_41794_, _41793_, _41792_);
  nand _49349_ (_41795_, _41794_, _41755_);
  or _49350_ (_41796_, \oc8051_gm_cxrom_1.cell4.data [0], _41755_);
  and _49351_ (_01627_, _41796_, _41795_);
  or _49352_ (_41797_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or _49353_ (_41798_, \oc8051_gm_cxrom_1.cell4.data [1], _41787_);
  nand _49354_ (_41799_, _41798_, _41797_);
  nand _49355_ (_41800_, _41799_, _41755_);
  or _49356_ (_41801_, \oc8051_gm_cxrom_1.cell4.data [1], _41755_);
  and _49357_ (_01631_, _41801_, _41800_);
  or _49358_ (_41802_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or _49359_ (_41803_, \oc8051_gm_cxrom_1.cell4.data [2], _41787_);
  nand _49360_ (_41804_, _41803_, _41802_);
  nand _49361_ (_41805_, _41804_, _41755_);
  or _49362_ (_41806_, \oc8051_gm_cxrom_1.cell4.data [2], _41755_);
  and _49363_ (_01635_, _41806_, _41805_);
  or _49364_ (_41807_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or _49365_ (_41808_, \oc8051_gm_cxrom_1.cell4.data [3], _41787_);
  nand _49366_ (_41809_, _41808_, _41807_);
  nand _49367_ (_41810_, _41809_, _41755_);
  or _49368_ (_41811_, \oc8051_gm_cxrom_1.cell4.data [3], _41755_);
  and _49369_ (_01639_, _41811_, _41810_);
  or _49370_ (_41812_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or _49371_ (_41813_, \oc8051_gm_cxrom_1.cell4.data [4], _41787_);
  nand _49372_ (_41814_, _41813_, _41812_);
  nand _49373_ (_41815_, _41814_, _41755_);
  or _49374_ (_41816_, \oc8051_gm_cxrom_1.cell4.data [4], _41755_);
  and _49375_ (_01643_, _41816_, _41815_);
  or _49376_ (_41817_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or _49377_ (_41818_, \oc8051_gm_cxrom_1.cell4.data [5], _41787_);
  nand _49378_ (_41819_, _41818_, _41817_);
  nand _49379_ (_41820_, _41819_, _41755_);
  or _49380_ (_41821_, \oc8051_gm_cxrom_1.cell4.data [5], _41755_);
  and _49381_ (_01647_, _41821_, _41820_);
  or _49382_ (_41822_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or _49383_ (_41823_, \oc8051_gm_cxrom_1.cell4.data [6], _41787_);
  nand _49384_ (_41824_, _41823_, _41822_);
  nand _49385_ (_41825_, _41824_, _41755_);
  or _49386_ (_41826_, \oc8051_gm_cxrom_1.cell4.data [6], _41755_);
  and _49387_ (_01651_, _41826_, _41825_);
  or _49388_ (_41827_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not _49389_ (_41828_, \oc8051_gm_cxrom_1.cell5.valid );
  or _49390_ (_41829_, _41828_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand _49391_ (_41830_, _41829_, _41827_);
  nand _49392_ (_41831_, _41830_, _41755_);
  or _49393_ (_41832_, \oc8051_gm_cxrom_1.cell5.data [7], _41755_);
  and _49394_ (_01673_, _41832_, _41831_);
  or _49395_ (_41833_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or _49396_ (_41834_, \oc8051_gm_cxrom_1.cell5.data [0], _41828_);
  nand _49397_ (_41835_, _41834_, _41833_);
  nand _49398_ (_41836_, _41835_, _41755_);
  or _49399_ (_41837_, \oc8051_gm_cxrom_1.cell5.data [0], _41755_);
  and _49400_ (_01680_, _41837_, _41836_);
  or _49401_ (_41838_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or _49402_ (_41839_, \oc8051_gm_cxrom_1.cell5.data [1], _41828_);
  nand _49403_ (_41840_, _41839_, _41838_);
  nand _49404_ (_41841_, _41840_, _41755_);
  or _49405_ (_41842_, \oc8051_gm_cxrom_1.cell5.data [1], _41755_);
  and _49406_ (_01684_, _41842_, _41841_);
  or _49407_ (_41843_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or _49408_ (_41844_, \oc8051_gm_cxrom_1.cell5.data [2], _41828_);
  nand _49409_ (_41845_, _41844_, _41843_);
  nand _49410_ (_41846_, _41845_, _41755_);
  or _49411_ (_41847_, \oc8051_gm_cxrom_1.cell5.data [2], _41755_);
  and _49412_ (_01688_, _41847_, _41846_);
  or _49413_ (_41848_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or _49414_ (_41849_, \oc8051_gm_cxrom_1.cell5.data [3], _41828_);
  nand _49415_ (_41850_, _41849_, _41848_);
  nand _49416_ (_41851_, _41850_, _41755_);
  or _49417_ (_41852_, \oc8051_gm_cxrom_1.cell5.data [3], _41755_);
  and _49418_ (_01692_, _41852_, _41851_);
  or _49419_ (_41853_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or _49420_ (_41854_, \oc8051_gm_cxrom_1.cell5.data [4], _41828_);
  nand _49421_ (_41855_, _41854_, _41853_);
  nand _49422_ (_41856_, _41855_, _41755_);
  or _49423_ (_41857_, \oc8051_gm_cxrom_1.cell5.data [4], _41755_);
  and _49424_ (_01696_, _41857_, _41856_);
  or _49425_ (_41858_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or _49426_ (_41859_, \oc8051_gm_cxrom_1.cell5.data [5], _41828_);
  nand _49427_ (_41860_, _41859_, _41858_);
  nand _49428_ (_41861_, _41860_, _41755_);
  or _49429_ (_41862_, \oc8051_gm_cxrom_1.cell5.data [5], _41755_);
  and _49430_ (_01700_, _41862_, _41861_);
  or _49431_ (_41863_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or _49432_ (_41864_, \oc8051_gm_cxrom_1.cell5.data [6], _41828_);
  nand _49433_ (_41865_, _41864_, _41863_);
  nand _49434_ (_41866_, _41865_, _41755_);
  or _49435_ (_41867_, \oc8051_gm_cxrom_1.cell5.data [6], _41755_);
  and _49436_ (_01704_, _41867_, _41866_);
  or _49437_ (_41868_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not _49438_ (_41869_, \oc8051_gm_cxrom_1.cell6.valid );
  or _49439_ (_41870_, _41869_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand _49440_ (_41871_, _41870_, _41868_);
  nand _49441_ (_41872_, _41871_, _41755_);
  or _49442_ (_41873_, \oc8051_gm_cxrom_1.cell6.data [7], _41755_);
  and _49443_ (_01725_, _41873_, _41872_);
  or _49444_ (_41874_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or _49445_ (_41875_, \oc8051_gm_cxrom_1.cell6.data [0], _41869_);
  nand _49446_ (_41876_, _41875_, _41874_);
  nand _49447_ (_41877_, _41876_, _41755_);
  or _49448_ (_41878_, \oc8051_gm_cxrom_1.cell6.data [0], _41755_);
  and _49449_ (_01732_, _41878_, _41877_);
  or _49450_ (_41879_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or _49451_ (_41880_, \oc8051_gm_cxrom_1.cell6.data [1], _41869_);
  nand _49452_ (_41881_, _41880_, _41879_);
  nand _49453_ (_41882_, _41881_, _41755_);
  or _49454_ (_41883_, \oc8051_gm_cxrom_1.cell6.data [1], _41755_);
  and _49455_ (_01736_, _41883_, _41882_);
  or _49456_ (_41884_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or _49457_ (_41885_, \oc8051_gm_cxrom_1.cell6.data [2], _41869_);
  nand _49458_ (_41886_, _41885_, _41884_);
  nand _49459_ (_41887_, _41886_, _41755_);
  or _49460_ (_41888_, \oc8051_gm_cxrom_1.cell6.data [2], _41755_);
  and _49461_ (_01740_, _41888_, _41887_);
  or _49462_ (_41889_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or _49463_ (_41890_, \oc8051_gm_cxrom_1.cell6.data [3], _41869_);
  nand _49464_ (_41891_, _41890_, _41889_);
  nand _49465_ (_41892_, _41891_, _41755_);
  or _49466_ (_41893_, \oc8051_gm_cxrom_1.cell6.data [3], _41755_);
  and _49467_ (_01744_, _41893_, _41892_);
  or _49468_ (_41894_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or _49469_ (_41895_, \oc8051_gm_cxrom_1.cell6.data [4], _41869_);
  nand _49470_ (_41896_, _41895_, _41894_);
  nand _49471_ (_41897_, _41896_, _41755_);
  or _49472_ (_41898_, \oc8051_gm_cxrom_1.cell6.data [4], _41755_);
  and _49473_ (_01748_, _41898_, _41897_);
  or _49474_ (_41899_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or _49475_ (_41900_, \oc8051_gm_cxrom_1.cell6.data [5], _41869_);
  nand _49476_ (_41901_, _41900_, _41899_);
  nand _49477_ (_41902_, _41901_, _41755_);
  or _49478_ (_41903_, \oc8051_gm_cxrom_1.cell6.data [5], _41755_);
  and _49479_ (_01752_, _41903_, _41902_);
  or _49480_ (_41904_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or _49481_ (_41905_, \oc8051_gm_cxrom_1.cell6.data [6], _41869_);
  nand _49482_ (_41906_, _41905_, _41904_);
  nand _49483_ (_41907_, _41906_, _41755_);
  or _49484_ (_41908_, \oc8051_gm_cxrom_1.cell6.data [6], _41755_);
  and _49485_ (_01756_, _41908_, _41907_);
  or _49486_ (_41909_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not _49487_ (_41910_, \oc8051_gm_cxrom_1.cell7.valid );
  or _49488_ (_41911_, _41910_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand _49489_ (_41912_, _41911_, _41909_);
  nand _49490_ (_41913_, _41912_, _41755_);
  or _49491_ (_41914_, \oc8051_gm_cxrom_1.cell7.data [7], _41755_);
  and _49492_ (_01777_, _41914_, _41913_);
  or _49493_ (_41915_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or _49494_ (_41916_, \oc8051_gm_cxrom_1.cell7.data [0], _41910_);
  nand _49495_ (_41917_, _41916_, _41915_);
  nand _49496_ (_41918_, _41917_, _41755_);
  or _49497_ (_41919_, \oc8051_gm_cxrom_1.cell7.data [0], _41755_);
  and _49498_ (_01784_, _41919_, _41918_);
  or _49499_ (_41920_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or _49500_ (_41921_, \oc8051_gm_cxrom_1.cell7.data [1], _41910_);
  nand _49501_ (_41922_, _41921_, _41920_);
  nand _49502_ (_41923_, _41922_, _41755_);
  or _49503_ (_41924_, \oc8051_gm_cxrom_1.cell7.data [1], _41755_);
  and _49504_ (_01788_, _41924_, _41923_);
  or _49505_ (_41925_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or _49506_ (_41926_, \oc8051_gm_cxrom_1.cell7.data [2], _41910_);
  nand _49507_ (_41927_, _41926_, _41925_);
  nand _49508_ (_41928_, _41927_, _41755_);
  or _49509_ (_41929_, \oc8051_gm_cxrom_1.cell7.data [2], _41755_);
  and _49510_ (_01792_, _41929_, _41928_);
  or _49511_ (_41930_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or _49512_ (_41931_, \oc8051_gm_cxrom_1.cell7.data [3], _41910_);
  nand _49513_ (_41932_, _41931_, _41930_);
  nand _49514_ (_41933_, _41932_, _41755_);
  or _49515_ (_41934_, \oc8051_gm_cxrom_1.cell7.data [3], _41755_);
  and _49516_ (_01795_, _41934_, _41933_);
  or _49517_ (_41935_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or _49518_ (_41936_, \oc8051_gm_cxrom_1.cell7.data [4], _41910_);
  nand _49519_ (_41937_, _41936_, _41935_);
  nand _49520_ (_41938_, _41937_, _41755_);
  or _49521_ (_41939_, \oc8051_gm_cxrom_1.cell7.data [4], _41755_);
  and _49522_ (_01799_, _41939_, _41938_);
  or _49523_ (_41940_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or _49524_ (_41941_, \oc8051_gm_cxrom_1.cell7.data [5], _41910_);
  nand _49525_ (_41942_, _41941_, _41940_);
  nand _49526_ (_41943_, _41942_, _41755_);
  or _49527_ (_41944_, \oc8051_gm_cxrom_1.cell7.data [5], _41755_);
  and _49528_ (_01803_, _41944_, _41943_);
  or _49529_ (_41945_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or _49530_ (_41946_, \oc8051_gm_cxrom_1.cell7.data [6], _41910_);
  nand _49531_ (_41947_, _41946_, _41945_);
  nand _49532_ (_41948_, _41947_, _41755_);
  or _49533_ (_41949_, \oc8051_gm_cxrom_1.cell7.data [6], _41755_);
  and _49534_ (_01807_, _41949_, _41948_);
  or _49535_ (_41950_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not _49536_ (_41951_, \oc8051_gm_cxrom_1.cell8.valid );
  or _49537_ (_41952_, _41951_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand _49538_ (_41953_, _41952_, _41950_);
  nand _49539_ (_41954_, _41953_, _41755_);
  or _49540_ (_41955_, \oc8051_gm_cxrom_1.cell8.data [7], _41755_);
  and _49541_ (_01828_, _41955_, _41954_);
  or _49542_ (_41956_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or _49543_ (_41957_, \oc8051_gm_cxrom_1.cell8.data [0], _41951_);
  nand _49544_ (_41958_, _41957_, _41956_);
  nand _49545_ (_41959_, _41958_, _41755_);
  or _49546_ (_41960_, \oc8051_gm_cxrom_1.cell8.data [0], _41755_);
  and _49547_ (_01835_, _41960_, _41959_);
  or _49548_ (_41961_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or _49549_ (_41962_, \oc8051_gm_cxrom_1.cell8.data [1], _41951_);
  nand _49550_ (_41963_, _41962_, _41961_);
  nand _49551_ (_41964_, _41963_, _41755_);
  or _49552_ (_41965_, \oc8051_gm_cxrom_1.cell8.data [1], _41755_);
  and _49553_ (_01839_, _41965_, _41964_);
  or _49554_ (_41966_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or _49555_ (_41967_, \oc8051_gm_cxrom_1.cell8.data [2], _41951_);
  nand _49556_ (_41968_, _41967_, _41966_);
  nand _49557_ (_41969_, _41968_, _41755_);
  or _49558_ (_41970_, \oc8051_gm_cxrom_1.cell8.data [2], _41755_);
  and _49559_ (_01843_, _41970_, _41969_);
  or _49560_ (_41971_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or _49561_ (_41972_, \oc8051_gm_cxrom_1.cell8.data [3], _41951_);
  nand _49562_ (_41973_, _41972_, _41971_);
  nand _49563_ (_41974_, _41973_, _41755_);
  or _49564_ (_41975_, \oc8051_gm_cxrom_1.cell8.data [3], _41755_);
  and _49565_ (_01847_, _41975_, _41974_);
  or _49566_ (_41976_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or _49567_ (_41977_, \oc8051_gm_cxrom_1.cell8.data [4], _41951_);
  nand _49568_ (_41978_, _41977_, _41976_);
  nand _49569_ (_41979_, _41978_, _41755_);
  or _49570_ (_41980_, \oc8051_gm_cxrom_1.cell8.data [4], _41755_);
  and _49571_ (_01851_, _41980_, _41979_);
  or _49572_ (_41981_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or _49573_ (_41982_, \oc8051_gm_cxrom_1.cell8.data [5], _41951_);
  nand _49574_ (_41983_, _41982_, _41981_);
  nand _49575_ (_41984_, _41983_, _41755_);
  or _49576_ (_41985_, \oc8051_gm_cxrom_1.cell8.data [5], _41755_);
  and _49577_ (_01855_, _41985_, _41984_);
  or _49578_ (_41986_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or _49579_ (_41987_, \oc8051_gm_cxrom_1.cell8.data [6], _41951_);
  nand _49580_ (_41988_, _41987_, _41986_);
  nand _49581_ (_41989_, _41988_, _41755_);
  or _49582_ (_41990_, \oc8051_gm_cxrom_1.cell8.data [6], _41755_);
  and _49583_ (_01859_, _41990_, _41989_);
  or _49584_ (_41991_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not _49585_ (_41992_, \oc8051_gm_cxrom_1.cell9.valid );
  or _49586_ (_41993_, _41992_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand _49587_ (_41994_, _41993_, _41991_);
  nand _49588_ (_41995_, _41994_, _41755_);
  or _49589_ (_41996_, \oc8051_gm_cxrom_1.cell9.data [7], _41755_);
  and _49590_ (_01881_, _41996_, _41995_);
  or _49591_ (_41997_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or _49592_ (_41998_, \oc8051_gm_cxrom_1.cell9.data [0], _41992_);
  nand _49593_ (_41999_, _41998_, _41997_);
  nand _49594_ (_42000_, _41999_, _41755_);
  or _49595_ (_42001_, \oc8051_gm_cxrom_1.cell9.data [0], _41755_);
  and _49596_ (_01887_, _42001_, _42000_);
  or _49597_ (_42002_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or _49598_ (_42003_, \oc8051_gm_cxrom_1.cell9.data [1], _41992_);
  nand _49599_ (_42004_, _42003_, _42002_);
  nand _49600_ (_42005_, _42004_, _41755_);
  or _49601_ (_42006_, \oc8051_gm_cxrom_1.cell9.data [1], _41755_);
  and _49602_ (_01891_, _42006_, _42005_);
  or _49603_ (_42007_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or _49604_ (_42008_, \oc8051_gm_cxrom_1.cell9.data [2], _41992_);
  nand _49605_ (_42009_, _42008_, _42007_);
  nand _49606_ (_42010_, _42009_, _41755_);
  or _49607_ (_42011_, \oc8051_gm_cxrom_1.cell9.data [2], _41755_);
  and _49608_ (_01895_, _42011_, _42010_);
  or _49609_ (_42012_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or _49610_ (_42013_, \oc8051_gm_cxrom_1.cell9.data [3], _41992_);
  nand _49611_ (_42014_, _42013_, _42012_);
  nand _49612_ (_42015_, _42014_, _41755_);
  or _49613_ (_42016_, \oc8051_gm_cxrom_1.cell9.data [3], _41755_);
  and _49614_ (_01899_, _42016_, _42015_);
  or _49615_ (_42017_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or _49616_ (_42018_, \oc8051_gm_cxrom_1.cell9.data [4], _41992_);
  nand _49617_ (_42019_, _42018_, _42017_);
  nand _49618_ (_42020_, _42019_, _41755_);
  or _49619_ (_42021_, \oc8051_gm_cxrom_1.cell9.data [4], _41755_);
  and _49620_ (_01903_, _42021_, _42020_);
  or _49621_ (_42022_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or _49622_ (_42023_, \oc8051_gm_cxrom_1.cell9.data [5], _41992_);
  nand _49623_ (_42024_, _42023_, _42022_);
  nand _49624_ (_42025_, _42024_, _41755_);
  or _49625_ (_42026_, \oc8051_gm_cxrom_1.cell9.data [5], _41755_);
  and _49626_ (_01907_, _42026_, _42025_);
  or _49627_ (_42027_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or _49628_ (_42028_, \oc8051_gm_cxrom_1.cell9.data [6], _41992_);
  nand _49629_ (_42029_, _42028_, _42027_);
  nand _49630_ (_42030_, _42029_, _41755_);
  or _49631_ (_42031_, \oc8051_gm_cxrom_1.cell9.data [6], _41755_);
  and _49632_ (_01911_, _42031_, _42030_);
  or _49633_ (_42032_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not _49634_ (_42033_, \oc8051_gm_cxrom_1.cell10.valid );
  or _49635_ (_42034_, _42033_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand _49636_ (_42035_, _42034_, _42032_);
  nand _49637_ (_42036_, _42035_, _41755_);
  or _49638_ (_42037_, \oc8051_gm_cxrom_1.cell10.data [7], _41755_);
  and _49639_ (_01933_, _42037_, _42036_);
  or _49640_ (_42038_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or _49641_ (_42039_, \oc8051_gm_cxrom_1.cell10.data [0], _42033_);
  nand _49642_ (_42040_, _42039_, _42038_);
  nand _49643_ (_42041_, _42040_, _41755_);
  or _49644_ (_42042_, \oc8051_gm_cxrom_1.cell10.data [0], _41755_);
  and _49645_ (_01940_, _42042_, _42041_);
  or _49646_ (_42043_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or _49647_ (_42044_, \oc8051_gm_cxrom_1.cell10.data [1], _42033_);
  nand _49648_ (_42045_, _42044_, _42043_);
  nand _49649_ (_42046_, _42045_, _41755_);
  or _49650_ (_42047_, \oc8051_gm_cxrom_1.cell10.data [1], _41755_);
  and _49651_ (_01943_, _42047_, _42046_);
  or _49652_ (_42048_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or _49653_ (_42049_, \oc8051_gm_cxrom_1.cell10.data [2], _42033_);
  nand _49654_ (_42050_, _42049_, _42048_);
  nand _49655_ (_42051_, _42050_, _41755_);
  or _49656_ (_42052_, \oc8051_gm_cxrom_1.cell10.data [2], _41755_);
  and _49657_ (_01947_, _42052_, _42051_);
  or _49658_ (_42053_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or _49659_ (_42054_, \oc8051_gm_cxrom_1.cell10.data [3], _42033_);
  nand _49660_ (_42055_, _42054_, _42053_);
  nand _49661_ (_42056_, _42055_, _41755_);
  or _49662_ (_42057_, \oc8051_gm_cxrom_1.cell10.data [3], _41755_);
  and _49663_ (_01951_, _42057_, _42056_);
  or _49664_ (_42058_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or _49665_ (_42059_, \oc8051_gm_cxrom_1.cell10.data [4], _42033_);
  nand _49666_ (_42060_, _42059_, _42058_);
  nand _49667_ (_42061_, _42060_, _41755_);
  or _49668_ (_42062_, \oc8051_gm_cxrom_1.cell10.data [4], _41755_);
  and _49669_ (_01955_, _42062_, _42061_);
  or _49670_ (_42063_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or _49671_ (_42064_, \oc8051_gm_cxrom_1.cell10.data [5], _42033_);
  nand _49672_ (_42065_, _42064_, _42063_);
  nand _49673_ (_42066_, _42065_, _41755_);
  or _49674_ (_42067_, \oc8051_gm_cxrom_1.cell10.data [5], _41755_);
  and _49675_ (_01959_, _42067_, _42066_);
  or _49676_ (_42068_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or _49677_ (_42069_, \oc8051_gm_cxrom_1.cell10.data [6], _42033_);
  nand _49678_ (_42070_, _42069_, _42068_);
  nand _49679_ (_42071_, _42070_, _41755_);
  or _49680_ (_42072_, \oc8051_gm_cxrom_1.cell10.data [6], _41755_);
  and _49681_ (_01963_, _42072_, _42071_);
  or _49682_ (_42073_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not _49683_ (_42074_, \oc8051_gm_cxrom_1.cell11.valid );
  or _49684_ (_42075_, _42074_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand _49685_ (_42076_, _42075_, _42073_);
  nand _49686_ (_42077_, _42076_, _41755_);
  or _49687_ (_42078_, \oc8051_gm_cxrom_1.cell11.data [7], _41755_);
  and _49688_ (_01985_, _42078_, _42077_);
  or _49689_ (_42079_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or _49690_ (_42080_, \oc8051_gm_cxrom_1.cell11.data [0], _42074_);
  nand _49691_ (_42081_, _42080_, _42079_);
  nand _49692_ (_42082_, _42081_, _41755_);
  or _49693_ (_42083_, \oc8051_gm_cxrom_1.cell11.data [0], _41755_);
  and _49694_ (_01992_, _42083_, _42082_);
  or _49695_ (_42084_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or _49696_ (_42085_, \oc8051_gm_cxrom_1.cell11.data [1], _42074_);
  nand _49697_ (_42086_, _42085_, _42084_);
  nand _49698_ (_42087_, _42086_, _41755_);
  or _49699_ (_42088_, \oc8051_gm_cxrom_1.cell11.data [1], _41755_);
  and _49700_ (_01996_, _42088_, _42087_);
  or _49701_ (_42089_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or _49702_ (_42090_, \oc8051_gm_cxrom_1.cell11.data [2], _42074_);
  nand _49703_ (_42091_, _42090_, _42089_);
  nand _49704_ (_42092_, _42091_, _41755_);
  or _49705_ (_42093_, \oc8051_gm_cxrom_1.cell11.data [2], _41755_);
  and _49706_ (_01999_, _42093_, _42092_);
  or _49707_ (_42094_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or _49708_ (_42095_, \oc8051_gm_cxrom_1.cell11.data [3], _42074_);
  nand _49709_ (_42096_, _42095_, _42094_);
  nand _49710_ (_42097_, _42096_, _41755_);
  or _49711_ (_42098_, \oc8051_gm_cxrom_1.cell11.data [3], _41755_);
  and _49712_ (_02003_, _42098_, _42097_);
  or _49713_ (_42099_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or _49714_ (_42100_, \oc8051_gm_cxrom_1.cell11.data [4], _42074_);
  nand _49715_ (_42101_, _42100_, _42099_);
  nand _49716_ (_42102_, _42101_, _41755_);
  or _49717_ (_42103_, \oc8051_gm_cxrom_1.cell11.data [4], _41755_);
  and _49718_ (_02007_, _42103_, _42102_);
  or _49719_ (_42104_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or _49720_ (_42105_, \oc8051_gm_cxrom_1.cell11.data [5], _42074_);
  nand _49721_ (_42106_, _42105_, _42104_);
  nand _49722_ (_42107_, _42106_, _41755_);
  or _49723_ (_42108_, \oc8051_gm_cxrom_1.cell11.data [5], _41755_);
  and _49724_ (_02011_, _42108_, _42107_);
  or _49725_ (_42109_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or _49726_ (_42110_, \oc8051_gm_cxrom_1.cell11.data [6], _42074_);
  nand _49727_ (_42111_, _42110_, _42109_);
  nand _49728_ (_42112_, _42111_, _41755_);
  or _49729_ (_42113_, \oc8051_gm_cxrom_1.cell11.data [6], _41755_);
  and _49730_ (_02015_, _42113_, _42112_);
  or _49731_ (_42114_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not _49732_ (_42115_, \oc8051_gm_cxrom_1.cell12.valid );
  or _49733_ (_42116_, _42115_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand _49734_ (_42117_, _42116_, _42114_);
  nand _49735_ (_42118_, _42117_, _41755_);
  or _49736_ (_42119_, \oc8051_gm_cxrom_1.cell12.data [7], _41755_);
  and _49737_ (_02037_, _42119_, _42118_);
  or _49738_ (_42120_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or _49739_ (_42121_, \oc8051_gm_cxrom_1.cell12.data [0], _42115_);
  nand _49740_ (_42122_, _42121_, _42120_);
  nand _49741_ (_42123_, _42122_, _41755_);
  or _49742_ (_42124_, \oc8051_gm_cxrom_1.cell12.data [0], _41755_);
  and _49743_ (_02044_, _42124_, _42123_);
  or _49744_ (_42125_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or _49745_ (_42126_, \oc8051_gm_cxrom_1.cell12.data [1], _42115_);
  nand _49746_ (_42127_, _42126_, _42125_);
  nand _49747_ (_42128_, _42127_, _41755_);
  or _49748_ (_42129_, \oc8051_gm_cxrom_1.cell12.data [1], _41755_);
  and _49749_ (_02048_, _42129_, _42128_);
  or _49750_ (_42130_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or _49751_ (_42131_, \oc8051_gm_cxrom_1.cell12.data [2], _42115_);
  nand _49752_ (_42132_, _42131_, _42130_);
  nand _49753_ (_42133_, _42132_, _41755_);
  or _49754_ (_42134_, \oc8051_gm_cxrom_1.cell12.data [2], _41755_);
  and _49755_ (_02052_, _42134_, _42133_);
  or _49756_ (_42135_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or _49757_ (_42136_, \oc8051_gm_cxrom_1.cell12.data [3], _42115_);
  nand _49758_ (_42137_, _42136_, _42135_);
  nand _49759_ (_42138_, _42137_, _41755_);
  or _49760_ (_42139_, \oc8051_gm_cxrom_1.cell12.data [3], _41755_);
  and _49761_ (_02055_, _42139_, _42138_);
  or _49762_ (_42140_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or _49763_ (_42141_, \oc8051_gm_cxrom_1.cell12.data [4], _42115_);
  nand _49764_ (_42142_, _42141_, _42140_);
  nand _49765_ (_42143_, _42142_, _41755_);
  or _49766_ (_42144_, \oc8051_gm_cxrom_1.cell12.data [4], _41755_);
  and _49767_ (_02059_, _42144_, _42143_);
  or _49768_ (_42145_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or _49769_ (_42146_, \oc8051_gm_cxrom_1.cell12.data [5], _42115_);
  nand _49770_ (_42147_, _42146_, _42145_);
  nand _49771_ (_42148_, _42147_, _41755_);
  or _49772_ (_42149_, \oc8051_gm_cxrom_1.cell12.data [5], _41755_);
  and _49773_ (_02063_, _42149_, _42148_);
  or _49774_ (_42150_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or _49775_ (_42151_, \oc8051_gm_cxrom_1.cell12.data [6], _42115_);
  nand _49776_ (_42152_, _42151_, _42150_);
  nand _49777_ (_42153_, _42152_, _41755_);
  or _49778_ (_42154_, \oc8051_gm_cxrom_1.cell12.data [6], _41755_);
  and _49779_ (_02067_, _42154_, _42153_);
  or _49780_ (_42155_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not _49781_ (_42156_, \oc8051_gm_cxrom_1.cell13.valid );
  or _49782_ (_42157_, _42156_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand _49783_ (_42158_, _42157_, _42155_);
  nand _49784_ (_42159_, _42158_, _41755_);
  or _49785_ (_42160_, \oc8051_gm_cxrom_1.cell13.data [7], _41755_);
  and _49786_ (_02089_, _42160_, _42159_);
  or _49787_ (_42161_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or _49788_ (_42162_, \oc8051_gm_cxrom_1.cell13.data [0], _42156_);
  nand _49789_ (_42163_, _42162_, _42161_);
  nand _49790_ (_42164_, _42163_, _41755_);
  or _49791_ (_42165_, \oc8051_gm_cxrom_1.cell13.data [0], _41755_);
  and _49792_ (_02096_, _42165_, _42164_);
  or _49793_ (_42166_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or _49794_ (_42167_, \oc8051_gm_cxrom_1.cell13.data [1], _42156_);
  nand _49795_ (_42168_, _42167_, _42166_);
  nand _49796_ (_42169_, _42168_, _41755_);
  or _49797_ (_42170_, \oc8051_gm_cxrom_1.cell13.data [1], _41755_);
  and _49798_ (_02100_, _42170_, _42169_);
  or _49799_ (_42171_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or _49800_ (_42172_, \oc8051_gm_cxrom_1.cell13.data [2], _42156_);
  nand _49801_ (_42173_, _42172_, _42171_);
  nand _49802_ (_42174_, _42173_, _41755_);
  or _49803_ (_42175_, \oc8051_gm_cxrom_1.cell13.data [2], _41755_);
  and _49804_ (_02104_, _42175_, _42174_);
  or _49805_ (_42176_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or _49806_ (_42177_, \oc8051_gm_cxrom_1.cell13.data [3], _42156_);
  nand _49807_ (_42178_, _42177_, _42176_);
  nand _49808_ (_42179_, _42178_, _41755_);
  or _49809_ (_42180_, \oc8051_gm_cxrom_1.cell13.data [3], _41755_);
  and _49810_ (_02108_, _42180_, _42179_);
  or _49811_ (_42181_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or _49812_ (_42182_, \oc8051_gm_cxrom_1.cell13.data [4], _42156_);
  nand _49813_ (_42183_, _42182_, _42181_);
  nand _49814_ (_42184_, _42183_, _41755_);
  or _49815_ (_42185_, \oc8051_gm_cxrom_1.cell13.data [4], _41755_);
  and _49816_ (_02111_, _42185_, _42184_);
  or _49817_ (_42186_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or _49818_ (_42187_, \oc8051_gm_cxrom_1.cell13.data [5], _42156_);
  nand _49819_ (_42188_, _42187_, _42186_);
  nand _49820_ (_42189_, _42188_, _41755_);
  or _49821_ (_42190_, \oc8051_gm_cxrom_1.cell13.data [5], _41755_);
  and _49822_ (_02115_, _42190_, _42189_);
  or _49823_ (_42191_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or _49824_ (_42192_, \oc8051_gm_cxrom_1.cell13.data [6], _42156_);
  nand _49825_ (_42193_, _42192_, _42191_);
  nand _49826_ (_42194_, _42193_, _41755_);
  or _49827_ (_42195_, \oc8051_gm_cxrom_1.cell13.data [6], _41755_);
  and _49828_ (_02119_, _42195_, _42194_);
  or _49829_ (_42196_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not _49830_ (_42197_, \oc8051_gm_cxrom_1.cell14.valid );
  or _49831_ (_42198_, _42197_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand _49832_ (_42199_, _42198_, _42196_);
  nand _49833_ (_42200_, _42199_, _41755_);
  or _49834_ (_42201_, \oc8051_gm_cxrom_1.cell14.data [7], _41755_);
  and _49835_ (_02141_, _42201_, _42200_);
  or _49836_ (_42202_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or _49837_ (_42203_, \oc8051_gm_cxrom_1.cell14.data [0], _42197_);
  nand _49838_ (_42204_, _42203_, _42202_);
  nand _49839_ (_42205_, _42204_, _41755_);
  or _49840_ (_42206_, \oc8051_gm_cxrom_1.cell14.data [0], _41755_);
  and _49841_ (_02148_, _42206_, _42205_);
  or _49842_ (_42207_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or _49843_ (_42208_, \oc8051_gm_cxrom_1.cell14.data [1], _42197_);
  nand _49844_ (_42209_, _42208_, _42207_);
  nand _49845_ (_42210_, _42209_, _41755_);
  or _49846_ (_42211_, \oc8051_gm_cxrom_1.cell14.data [1], _41755_);
  and _49847_ (_02152_, _42211_, _42210_);
  or _49848_ (_42212_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or _49849_ (_42213_, \oc8051_gm_cxrom_1.cell14.data [2], _42197_);
  nand _49850_ (_42214_, _42213_, _42212_);
  nand _49851_ (_42215_, _42214_, _41755_);
  or _49852_ (_42216_, \oc8051_gm_cxrom_1.cell14.data [2], _41755_);
  and _49853_ (_02156_, _42216_, _42215_);
  or _49854_ (_42217_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or _49855_ (_42218_, \oc8051_gm_cxrom_1.cell14.data [3], _42197_);
  nand _49856_ (_42219_, _42218_, _42217_);
  nand _49857_ (_42220_, _42219_, _41755_);
  or _49858_ (_42221_, \oc8051_gm_cxrom_1.cell14.data [3], _41755_);
  and _49859_ (_02160_, _42221_, _42220_);
  or _49860_ (_42222_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or _49861_ (_42223_, \oc8051_gm_cxrom_1.cell14.data [4], _42197_);
  nand _49862_ (_42224_, _42223_, _42222_);
  nand _49863_ (_42225_, _42224_, _41755_);
  or _49864_ (_42226_, \oc8051_gm_cxrom_1.cell14.data [4], _41755_);
  and _49865_ (_02164_, _42226_, _42225_);
  or _49866_ (_42227_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or _49867_ (_42228_, \oc8051_gm_cxrom_1.cell14.data [5], _42197_);
  nand _49868_ (_42229_, _42228_, _42227_);
  nand _49869_ (_42230_, _42229_, _41755_);
  or _49870_ (_42231_, \oc8051_gm_cxrom_1.cell14.data [5], _41755_);
  and _49871_ (_02167_, _42231_, _42230_);
  or _49872_ (_42232_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or _49873_ (_42233_, \oc8051_gm_cxrom_1.cell14.data [6], _42197_);
  nand _49874_ (_42234_, _42233_, _42232_);
  nand _49875_ (_42235_, _42234_, _41755_);
  or _49876_ (_42236_, \oc8051_gm_cxrom_1.cell14.data [6], _41755_);
  and _49877_ (_02171_, _42236_, _42235_);
  or _49878_ (_42237_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not _49879_ (_42238_, \oc8051_gm_cxrom_1.cell15.valid );
  or _49880_ (_42239_, _42238_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand _49881_ (_42240_, _42239_, _42237_);
  nand _49882_ (_42241_, _42240_, _41755_);
  or _49883_ (_42242_, \oc8051_gm_cxrom_1.cell15.data [7], _41755_);
  and _49884_ (_02193_, _42242_, _42241_);
  or _49885_ (_42243_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or _49886_ (_42244_, \oc8051_gm_cxrom_1.cell15.data [0], _42238_);
  nand _49887_ (_42245_, _42244_, _42243_);
  nand _49888_ (_42246_, _42245_, _41755_);
  or _49889_ (_42247_, \oc8051_gm_cxrom_1.cell15.data [0], _41755_);
  and _49890_ (_02200_, _42247_, _42246_);
  or _49891_ (_42248_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or _49892_ (_42249_, \oc8051_gm_cxrom_1.cell15.data [1], _42238_);
  nand _49893_ (_42250_, _42249_, _42248_);
  nand _49894_ (_42251_, _42250_, _41755_);
  or _49895_ (_42252_, \oc8051_gm_cxrom_1.cell15.data [1], _41755_);
  and _49896_ (_02204_, _42252_, _42251_);
  or _49897_ (_42253_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or _49898_ (_42254_, \oc8051_gm_cxrom_1.cell15.data [2], _42238_);
  nand _49899_ (_42255_, _42254_, _42253_);
  nand _49900_ (_42256_, _42255_, _41755_);
  or _49901_ (_42257_, \oc8051_gm_cxrom_1.cell15.data [2], _41755_);
  and _49902_ (_02208_, _42257_, _42256_);
  or _49903_ (_42258_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or _49904_ (_42259_, \oc8051_gm_cxrom_1.cell15.data [3], _42238_);
  nand _49905_ (_42260_, _42259_, _42258_);
  nand _49906_ (_42261_, _42260_, _41755_);
  or _49907_ (_42262_, \oc8051_gm_cxrom_1.cell15.data [3], _41755_);
  and _49908_ (_02212_, _42262_, _42261_);
  or _49909_ (_42263_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or _49910_ (_42264_, \oc8051_gm_cxrom_1.cell15.data [4], _42238_);
  nand _49911_ (_42265_, _42264_, _42263_);
  nand _49912_ (_42266_, _42265_, _41755_);
  or _49913_ (_42267_, \oc8051_gm_cxrom_1.cell15.data [4], _41755_);
  and _49914_ (_02216_, _42267_, _42266_);
  or _49915_ (_42268_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or _49916_ (_42269_, \oc8051_gm_cxrom_1.cell15.data [5], _42238_);
  nand _49917_ (_42270_, _42269_, _42268_);
  nand _49918_ (_42271_, _42270_, _41755_);
  or _49919_ (_42272_, \oc8051_gm_cxrom_1.cell15.data [5], _41755_);
  and _49920_ (_02220_, _42272_, _42271_);
  or _49921_ (_42273_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or _49922_ (_42274_, \oc8051_gm_cxrom_1.cell15.data [6], _42238_);
  nand _49923_ (_42275_, _42274_, _42273_);
  nand _49924_ (_42276_, _42275_, _41755_);
  or _49925_ (_42277_, \oc8051_gm_cxrom_1.cell15.data [6], _41755_);
  and _49926_ (_02223_, _42277_, _42276_);
  nor _49927_ (_05997_, _37910_, rst);
  and _49928_ (_42278_, _33793_, _41755_);
  nand _49929_ (_42279_, _42278_, _36328_);
  nor _49930_ (_42280_, _36174_, _35004_);
  or _49931_ (_06000_, _42280_, _42279_);
  not _49932_ (_42281_, _34447_);
  and _49933_ (_42282_, _34938_, _34698_);
  and _49934_ (_42283_, _42282_, _42281_);
  not _49935_ (_42284_, _34185_);
  nor _49936_ (_42285_, _35213_, _35455_);
  not _49937_ (_42286_, _35701_);
  and _49938_ (_42287_, _35932_, _42286_);
  and _49939_ (_42288_, _42287_, _42285_);
  nor _49940_ (_42289_, _42288_, _42284_);
  and _49941_ (_42290_, _35932_, _35701_);
  not _49942_ (_42291_, _35455_);
  and _49943_ (_42292_, _35213_, _42291_);
  and _49944_ (_42293_, _42292_, _42290_);
  nor _49945_ (_42294_, _35213_, _42291_);
  and _49946_ (_42295_, _42294_, _42287_);
  nor _49947_ (_42296_, _42295_, _42293_);
  nand _49948_ (_42297_, _42296_, _42289_);
  and _49949_ (_42298_, _42297_, _42283_);
  nor _49950_ (_42299_, _42284_, _34447_);
  and _49951_ (_42300_, _42299_, _42282_);
  not _49952_ (_42301_, _35932_);
  and _49953_ (_42302_, _42301_, _35701_);
  and _49954_ (_42303_, _42302_, _42294_);
  and _49955_ (_42304_, _42303_, _42300_);
  and _49956_ (_42305_, _42302_, _42292_);
  not _49957_ (_42306_, _34938_);
  not _49958_ (_42307_, _34698_);
  and _49959_ (_42308_, _42307_, _34447_);
  nor _49960_ (_42309_, _42308_, _42306_);
  not _49961_ (_42310_, _42309_);
  and _49962_ (_42311_, _42310_, _42305_);
  nor _49963_ (_42312_, _42311_, _42304_);
  not _49964_ (_42313_, _42312_);
  or _49965_ (_42314_, _42313_, _42298_);
  not _49966_ (_42315_, _35213_);
  and _49967_ (_42316_, _34938_, _42307_);
  and _49968_ (_42317_, _42316_, _42299_);
  and _49969_ (_42318_, _42317_, _42315_);
  and _49970_ (_42319_, _42318_, _42302_);
  nor _49971_ (_42320_, _42294_, _42292_);
  and _49972_ (_42321_, _42320_, _42290_);
  and _49973_ (_42322_, _42321_, _42300_);
  nor _49974_ (_42323_, _35932_, _35701_);
  and _49975_ (_42324_, _42323_, _35455_);
  and _49976_ (_42325_, _42324_, _35213_);
  and _49977_ (_42326_, _42316_, _42281_);
  and _49978_ (_42327_, _42326_, _42284_);
  and _49979_ (_42328_, _42327_, _42325_);
  nor _49980_ (_42329_, _42328_, _42322_);
  not _49981_ (_42330_, _42329_);
  or _49982_ (_42331_, _42330_, _42319_);
  or _49983_ (_42332_, _42331_, _42314_);
  and _49984_ (_42333_, _42282_, _34447_);
  and _49985_ (_42334_, _42333_, _34185_);
  and _49986_ (_42335_, _42290_, _35455_);
  and _49987_ (_42336_, _42335_, _42334_);
  and _49988_ (_42337_, _34698_, _34447_);
  and _49989_ (_42338_, _42323_, _42291_);
  and _49990_ (_42339_, _42338_, _42337_);
  and _49991_ (_42340_, _42339_, _34938_);
  or _49992_ (_42341_, _42340_, _42336_);
  and _49993_ (_42342_, _42341_, _35213_);
  and _49994_ (_42343_, _35213_, _35455_);
  nand _49995_ (_42344_, _42334_, _42290_);
  or _49996_ (_42345_, _42344_, _42343_);
  and _49997_ (_42346_, _42338_, _42300_);
  and _49998_ (_42347_, _42292_, _42287_);
  and _49999_ (_42348_, _42333_, _42284_);
  and _50000_ (_42349_, _42348_, _42347_);
  and _50001_ (_42350_, _42325_, _42306_);
  or _50002_ (_42351_, _42350_, _42349_);
  nor _50003_ (_42352_, _42351_, _42346_);
  and _50004_ (_42353_, _42352_, _42345_);
  and _50005_ (_42354_, _42300_, _35213_);
  and _50006_ (_42355_, _42354_, _42287_);
  not _50007_ (_42356_, _42355_);
  nor _50008_ (_42357_, _35213_, _42306_);
  and _50009_ (_42358_, _42357_, _42339_);
  and _50010_ (_42359_, _42302_, _35455_);
  and _50011_ (_42360_, _42348_, _42359_);
  and _50012_ (_42361_, _42326_, _42305_);
  or _50013_ (_42362_, _42361_, _42360_);
  nor _50014_ (_42363_, _42362_, _42358_);
  and _50015_ (_42364_, _42363_, _42356_);
  nand _50016_ (_42365_, _42364_, _42353_);
  or _50017_ (_42366_, _42365_, _42342_);
  or _50018_ (_42367_, _42366_, _42332_);
  and _50019_ (_42368_, _42367_, _33804_);
  not _50020_ (_42369_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _50021_ (_42370_, _33782_, _15507_);
  and _50022_ (_42371_, _42370_, _36678_);
  nor _50023_ (_42372_, _42371_, _42369_);
  or _50024_ (_42373_, _42372_, rst);
  or _50025_ (_06003_, _42373_, _42368_);
  nand _50026_ (_42374_, _35932_, _33739_);
  or _50027_ (_42375_, _33739_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _50028_ (_42376_, _42375_, _41755_);
  and _50029_ (_06006_, _42376_, _42374_);
  and _50030_ (_42377_, \oc8051_top_1.oc8051_sfr1.wait_data , _41755_);
  and _50031_ (_42378_, _42377_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _50032_ (_42379_, _35015_, _37431_);
  and _50033_ (_42380_, _37811_, _36875_);
  or _50034_ (_42381_, _42380_, _42379_);
  and _50035_ (_42382_, _37431_, _36174_);
  or _50036_ (_42383_, _42382_, _37635_);
  or _50037_ (_42384_, _42383_, _37373_);
  and _50038_ (_42385_, _37372_, _35015_);
  and _50039_ (_42386_, _36218_, _35004_);
  or _50040_ (_42387_, _42386_, _42385_);
  or _50041_ (_42388_, _42387_, _42384_);
  or _50042_ (_42389_, _42388_, _37180_);
  or _50043_ (_42390_, _42389_, _42381_);
  and _50044_ (_42391_, _42390_, _42278_);
  or _50045_ (_06009_, _42391_, _42378_);
  and _50046_ (_42392_, _36174_, _36075_);
  or _50047_ (_42393_, _42392_, _36031_);
  and _50048_ (_42394_, _36995_, _36207_);
  or _50049_ (_42395_, _42394_, _36448_);
  and _50050_ (_42396_, _36842_, _34491_);
  and _50051_ (_42397_, _42396_, _37372_);
  or _50052_ (_42398_, _42397_, _42395_);
  or _50053_ (_42399_, _42398_, _42393_);
  and _50054_ (_42400_, _42399_, _33793_);
  and _50055_ (_42401_, \oc8051_top_1.oc8051_decoder1.state [0], _15507_);
  and _50056_ (_42402_, _42401_, _42369_);
  not _50057_ (_42403_, _37844_);
  and _50058_ (_42404_, _42403_, _42402_);
  and _50059_ (_42405_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50060_ (_42406_, _42405_, _42404_);
  or _50061_ (_42407_, _42406_, _42400_);
  and _50062_ (_06012_, _42407_, _41755_);
  and _50063_ (_42408_, _42377_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _50064_ (_42409_, _37811_, _37016_);
  nor _50065_ (_42410_, _37016_, _36218_);
  nor _50066_ (_42411_, _42410_, _37082_);
  or _50067_ (_42412_, _42411_, _42409_);
  and _50068_ (_42413_, _42396_, _37136_);
  or _50069_ (_42414_, _42413_, _42412_);
  and _50070_ (_42415_, _37136_, _36459_);
  nor _50071_ (_42416_, _42410_, _34982_);
  nor _50072_ (_42417_, _42416_, _42415_);
  nor _50073_ (_42418_, _35257_, _34982_);
  and _50074_ (_42419_, _42418_, _36009_);
  nor _50075_ (_42420_, _42419_, _36557_);
  nand _50076_ (_42421_, _42420_, _42417_);
  and _50077_ (_42422_, _37811_, _36897_);
  or _50078_ (_42423_, _42422_, _42393_);
  or _50079_ (_42424_, _42423_, _42421_);
  or _50080_ (_42425_, _42424_, _42414_);
  and _50081_ (_42426_, _42425_, _42278_);
  or _50082_ (_06015_, _42426_, _42408_);
  and _50083_ (_42427_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50084_ (_42428_, _37530_, _33793_);
  or _50085_ (_42429_, _42428_, _42427_);
  or _50086_ (_42430_, _42429_, _42404_);
  and _50087_ (_06018_, _42430_, _41755_);
  and _50088_ (_42431_, _35015_, _36064_);
  not _50089_ (_42432_, _36875_);
  nor _50090_ (_42433_, _42280_, _42432_);
  nor _50091_ (_42434_, _42433_, _42431_);
  not _50092_ (_42435_, _42434_);
  and _50093_ (_42436_, _42435_, _42402_);
  or _50094_ (_42437_, _42436_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50095_ (_42438_, _37136_, _36361_);
  and _50096_ (_42439_, _36853_, _34993_);
  and _50097_ (_42440_, _42439_, _36042_);
  or _50098_ (_42441_, _42440_, _42438_);
  or _50099_ (_42442_, _42441_, _42379_);
  and _50100_ (_42443_, _42441_, _36700_);
  or _50101_ (_42444_, _42443_, _37888_);
  and _50102_ (_42445_, _42444_, _42442_);
  or _50103_ (_42446_, _42445_, _42437_);
  or _50104_ (_42447_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15507_);
  and _50105_ (_42448_, _42447_, _41755_);
  and _50106_ (_06021_, _42448_, _42446_);
  and _50107_ (_42449_, _42377_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _50108_ (_42450_, _37372_, _37136_);
  and _50109_ (_42451_, _42450_, _36251_);
  and _50110_ (_42452_, _36218_, _36459_);
  or _50111_ (_42453_, _42452_, _42415_);
  or _50112_ (_42454_, _42453_, _42451_);
  and _50113_ (_42455_, _36361_, _36009_);
  or _50114_ (_42456_, _42413_, _42386_);
  or _50115_ (_42457_, _42456_, _42455_);
  or _50116_ (_42458_, _42394_, _37409_);
  or _50117_ (_42459_, _37318_, _36031_);
  or _50118_ (_42460_, _42459_, _42458_);
  or _50119_ (_42461_, _42460_, _42457_);
  or _50120_ (_42462_, _42461_, _42454_);
  and _50121_ (_42463_, _42462_, _42278_);
  or _50122_ (_06024_, _42463_, _42449_);
  and _50123_ (_42464_, _42377_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not _50124_ (_42465_, _42417_);
  or _50125_ (_42466_, _42397_, _37279_);
  and _50126_ (_42467_, _35015_, _36372_);
  and _50127_ (_42468_, _42396_, _36951_);
  or _50128_ (_42469_, _42468_, _42467_);
  or _50129_ (_42470_, _42469_, _42466_);
  or _50130_ (_42471_, _42470_, _42465_);
  and _50131_ (_42472_, _37811_, _37224_);
  or _50132_ (_42473_, _37310_, _37235_);
  or _50133_ (_42474_, _42473_, _42472_);
  and _50134_ (_42475_, _36196_, _36262_);
  or _50135_ (_42476_, _36405_, _42475_);
  and _50136_ (_42477_, _36218_, _36251_);
  or _50137_ (_42478_, _42477_, _42476_);
  or _50138_ (_42479_, _42478_, _42474_);
  or _50139_ (_42480_, _42479_, _42471_);
  and _50140_ (_42481_, _36995_, _36196_);
  and _50141_ (_42482_, _36995_, _36097_);
  or _50142_ (_42483_, _42482_, _42481_);
  not _50143_ (_42484_, _37356_);
  or _50144_ (_42485_, _36962_, _36525_);
  or _50145_ (_42486_, _42485_, _42484_);
  or _50146_ (_42487_, _42486_, _42483_);
  or _50147_ (_42488_, _42487_, _42414_);
  or _50148_ (_42489_, _42488_, _42480_);
  and _50149_ (_42490_, _42489_, _42278_);
  or _50150_ (_06027_, _42490_, _42464_);
  and _50151_ (_42491_, _42396_, _36383_);
  or _50152_ (_42492_, _42491_, _36492_);
  and _50153_ (_42493_, _42418_, _36064_);
  or _50154_ (_42494_, _42493_, _36601_);
  and _50155_ (_42495_, _36383_, _36459_);
  or _50156_ (_42496_, _42495_, _42494_);
  or _50157_ (_42497_, _42496_, _42492_);
  and _50158_ (_42498_, _42396_, _36075_);
  or _50159_ (_42499_, _42498_, _42497_);
  and _50160_ (_42500_, _42499_, _33793_);
  nor _50161_ (_42501_, _37844_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50162_ (_42502_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _50163_ (_42503_, _42502_, _42501_);
  or _50164_ (_42504_, _42503_, _42500_);
  and _50165_ (_06030_, _42504_, _41755_);
  or _50166_ (_42505_, _37497_, _37409_);
  not _50167_ (_42506_, _37541_);
  or _50168_ (_42507_, _42411_, _42506_);
  or _50169_ (_42508_, _42507_, _42505_);
  and _50170_ (_42509_, _36086_, _36042_);
  and _50171_ (_42510_, _42509_, _36864_);
  or _50172_ (_42511_, _42510_, _37257_);
  or _50173_ (_42512_, _42511_, _37235_);
  or _50174_ (_42513_, _42512_, _42438_);
  nand _50175_ (_42514_, _37374_, _36973_);
  or _50176_ (_42515_, _42514_, _42513_);
  or _50177_ (_42516_, _42515_, _42508_);
  and _50178_ (_42517_, _37431_, _36459_);
  and _50179_ (_42518_, _37431_, _36251_);
  or _50180_ (_42519_, _42440_, _42518_);
  or _50181_ (_42520_, _42519_, _42517_);
  or _50182_ (_42521_, _42520_, _37453_);
  and _50183_ (_42522_, _42509_, _36251_);
  or _50184_ (_42523_, _42522_, _36525_);
  or _50185_ (_42524_, _42523_, _36809_);
  and _50186_ (_42525_, _42418_, _36086_);
  or _50187_ (_42526_, _42525_, _37006_);
  or _50188_ (_42527_, _42526_, _42395_);
  or _50189_ (_42528_, _42527_, _42524_);
  or _50190_ (_42529_, _42528_, _42465_);
  or _50191_ (_42530_, _42529_, _42521_);
  or _50192_ (_42531_, _42530_, _42516_);
  and _50193_ (_42532_, _42531_, _33793_);
  or _50194_ (_42533_, _42443_, _42404_);
  and _50195_ (_42534_, _37690_, _36700_);
  or _50196_ (_42535_, _42534_, _42533_);
  and _50197_ (_42536_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50198_ (_42537_, _42536_, _42535_);
  or _50199_ (_42538_, _42537_, _42532_);
  and _50200_ (_06033_, _42538_, _41755_);
  nor _50201_ (_06092_, _36766_, rst);
  nor _50202_ (_06094_, _37756_, rst);
  not _50203_ (_42539_, _42278_);
  or _50204_ (_06097_, _42434_, _42539_);
  and _50205_ (_42540_, _36328_, _36174_);
  nor _50206_ (_42541_, _42540_, _42431_);
  or _50207_ (_06100_, _42541_, _42539_);
  and _50208_ (_42542_, _42290_, _42291_);
  and _50209_ (_42543_, _42334_, _42542_);
  or _50210_ (_42544_, _42360_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _50211_ (_42545_, _42544_, _42543_);
  or _50212_ (_42546_, _42545_, _42319_);
  and _50213_ (_42547_, _42546_, _42371_);
  nor _50214_ (_42548_, _42370_, _36678_);
  or _50215_ (_42549_, _42548_, rst);
  or _50216_ (_06103_, _42549_, _42547_);
  nand _50217_ (_42550_, _34185_, _33739_);
  or _50218_ (_42551_, _33739_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _50219_ (_42552_, _42551_, _41755_);
  and _50220_ (_06106_, _42552_, _42550_);
  not _50221_ (_42553_, _33739_);
  or _50222_ (_42554_, _34447_, _42553_);
  or _50223_ (_42555_, _33739_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _50224_ (_42556_, _42555_, _41755_);
  and _50225_ (_06109_, _42556_, _42554_);
  nand _50226_ (_42557_, _34698_, _33739_);
  or _50227_ (_42558_, _33739_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _50228_ (_42559_, _42558_, _41755_);
  and _50229_ (_06112_, _42559_, _42557_);
  nand _50230_ (_42560_, _34938_, _33739_);
  or _50231_ (_42561_, _33739_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _50232_ (_42562_, _42561_, _41755_);
  and _50233_ (_06115_, _42562_, _42560_);
  or _50234_ (_42563_, _35213_, _42553_);
  or _50235_ (_42564_, _33739_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _50236_ (_42565_, _42564_, _41755_);
  and _50237_ (_06118_, _42565_, _42563_);
  nand _50238_ (_42566_, _35455_, _33739_);
  or _50239_ (_42567_, _33739_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _50240_ (_42568_, _42567_, _41755_);
  and _50241_ (_06121_, _42568_, _42566_);
  nand _50242_ (_42569_, _35701_, _33739_);
  or _50243_ (_42570_, _33739_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _50244_ (_42571_, _42570_, _41755_);
  and _50245_ (_06124_, _42571_, _42569_);
  and _50246_ (_42572_, _42396_, _37224_);
  or _50247_ (_42573_, _42572_, _42392_);
  nor _50248_ (_42574_, _37071_, _34982_);
  or _50249_ (_42575_, _42574_, _42573_);
  or _50250_ (_42576_, _42396_, _36459_);
  or _50251_ (_42577_, _36875_, _36951_);
  and _50252_ (_42578_, _42577_, _42576_);
  or _50253_ (_42579_, _42578_, _42575_);
  and _50254_ (_42580_, _36951_, _36251_);
  or _50255_ (_42581_, _36031_, _42580_);
  or _50256_ (_42582_, _42494_, _42467_);
  or _50257_ (_42583_, _42582_, _42581_);
  or _50258_ (_42584_, _36218_, _36514_);
  and _50259_ (_42585_, _42584_, _37811_);
  and _50260_ (_42586_, _36075_, _36251_);
  or _50261_ (_42587_, _42491_, _42586_);
  and _50262_ (_42588_, _36995_, _36306_);
  or _50263_ (_42589_, _42588_, _42498_);
  or _50264_ (_42590_, _42589_, _42587_);
  or _50265_ (_42591_, _42590_, _42585_);
  or _50266_ (_42592_, _42591_, _42583_);
  and _50267_ (_42593_, _36579_, _36842_);
  and _50268_ (_42594_, _37811_, _36108_);
  and _50269_ (_42595_, _36328_, _36042_);
  and _50270_ (_42596_, _42595_, _37811_);
  or _50271_ (_42597_, _42596_, _42594_);
  nor _50272_ (_42598_, _42597_, _42593_);
  nand _50273_ (_42599_, _42598_, _36350_);
  or _50274_ (_42600_, _42599_, _42592_);
  or _50275_ (_42601_, _42600_, _42579_);
  and _50276_ (_42602_, _42601_, _33793_);
  and _50277_ (_42603_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50278_ (_42604_, _42603_, _42436_);
  or _50279_ (_42605_, _42604_, _42602_);
  and _50280_ (_30491_, _42605_, _41755_);
  and _50281_ (_42606_, _42377_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _50282_ (_42607_, _37224_, _36951_);
  and _50283_ (_42608_, _42607_, _36361_);
  or _50284_ (_42609_, _42573_, _42483_);
  or _50285_ (_42610_, _42609_, _42608_);
  nor _50286_ (_42611_, _42419_, _36536_);
  not _50287_ (_42612_, _42611_);
  nor _50288_ (_42613_, _42612_, _42422_);
  nand _50289_ (_42614_, _42613_, _37420_);
  or _50290_ (_42615_, _42614_, _42381_);
  not _50291_ (_42616_, _36951_);
  nand _50292_ (_42617_, _37071_, _42616_);
  and _50293_ (_42618_, _42617_, _37811_);
  or _50294_ (_42619_, _42618_, _42478_);
  or _50295_ (_42620_, _42619_, _42615_);
  or _50296_ (_42621_, _42620_, _42610_);
  and _50297_ (_42622_, _42621_, _42278_);
  or _50298_ (_30494_, _42622_, _42606_);
  or _50299_ (_42623_, _42521_, _42516_);
  and _50300_ (_42624_, _42623_, _33793_);
  and _50301_ (_42625_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50302_ (_42626_, _42625_, _42535_);
  or _50303_ (_42627_, _42626_, _42624_);
  and _50304_ (_30496_, _42627_, _41755_);
  and _50305_ (_42628_, _36940_, _35257_);
  or _50306_ (_42629_, _42628_, _36448_);
  or _50307_ (_42630_, _42629_, _42524_);
  or _50308_ (_42631_, _42630_, _42441_);
  and _50309_ (_42632_, _42631_, _33793_);
  and _50310_ (_42633_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50311_ (_42634_, _42633_, _42533_);
  or _50312_ (_42635_, _42634_, _42632_);
  and _50313_ (_30498_, _42635_, _41755_);
  or _50314_ (_42636_, _42574_, _42467_);
  or _50315_ (_42637_, _42494_, _36590_);
  or _50316_ (_42638_, _42607_, _36108_);
  and _50317_ (_42639_, _42638_, _37811_);
  or _50318_ (_42640_, _42639_, _42637_);
  or _50319_ (_42641_, _42640_, _42636_);
  and _50320_ (_42642_, _37811_, _37372_);
  or _50321_ (_42643_, _42596_, _37822_);
  or _50322_ (_42644_, _42643_, _42642_);
  and _50323_ (_42645_, _42396_, _37268_);
  or _50324_ (_42646_, _42645_, _42498_);
  or _50325_ (_42647_, _42646_, _42380_);
  or _50326_ (_42648_, _42647_, _42585_);
  or _50327_ (_42649_, _42648_, _42644_);
  and _50328_ (_42650_, _36108_, _35015_);
  and _50329_ (_42651_, _42491_, _35257_);
  or _50330_ (_42652_, _42651_, _42650_);
  or _50331_ (_42653_, _42525_, _42586_);
  or _50332_ (_42654_, _42653_, _42522_);
  and _50333_ (_42655_, _36579_, _36361_);
  and _50334_ (_42656_, _42595_, _36864_);
  or _50335_ (_42657_, _42656_, _42655_);
  or _50336_ (_42658_, _42657_, _42654_);
  or _50337_ (_42659_, _42658_, _42652_);
  and _50338_ (_42660_, _42396_, _37126_);
  or _50339_ (_42661_, _42660_, _42431_);
  and _50340_ (_42662_, _42396_, _36579_);
  or _50341_ (_42663_, _42662_, _37833_);
  or _50342_ (_42664_, _42663_, _42661_);
  or _50343_ (_42665_, _42664_, _42441_);
  or _50344_ (_42666_, _42665_, _42659_);
  or _50345_ (_42667_, _42666_, _42649_);
  or _50346_ (_42668_, _42667_, _42641_);
  and _50347_ (_42669_, _42668_, _33793_);
  and _50348_ (_42670_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50349_ (_42671_, _42436_, _37899_);
  or _50350_ (_42672_, _42671_, _42670_);
  or _50351_ (_42673_, _42672_, _42669_);
  and _50352_ (_30500_, _42673_, _41755_);
  and _50353_ (_42674_, _42418_, _36328_);
  and _50354_ (_42675_, _42595_, _36251_);
  or _50355_ (_42676_, _42675_, _37453_);
  or _50356_ (_42677_, _42676_, _42674_);
  or _50357_ (_42679_, _42677_, _42637_);
  or _50358_ (_42681_, _42679_, _42636_);
  or _50359_ (_42683_, _37833_, _42586_);
  or _50360_ (_42685_, _42510_, _42392_);
  or _50361_ (_42687_, _42685_, _42683_);
  or _50362_ (_42689_, _42687_, _36141_);
  and _50363_ (_42691_, _42607_, _35015_);
  or _50364_ (_42693_, _42691_, _37093_);
  or _50365_ (_42695_, _42693_, _42689_);
  or _50366_ (_42697_, _42695_, _42649_);
  or _50367_ (_42699_, _42697_, _42681_);
  and _50368_ (_42701_, _42699_, _33793_);
  and _50369_ (_42703_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50370_ (_42705_, _42703_, _42671_);
  or _50371_ (_42707_, _42705_, _42701_);
  and _50372_ (_30502_, _42707_, _41755_);
  and _50373_ (_42710_, _42377_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _50374_ (_42712_, _35015_, _36218_);
  and _50375_ (_42714_, _35015_, _36514_);
  and _50376_ (_42716_, _42714_, _36042_);
  or _50377_ (_42718_, _42716_, _42712_);
  or _50378_ (_42720_, _36240_, _36459_);
  or _50379_ (_42722_, _42720_, _35015_);
  and _50380_ (_42724_, _35015_, _37268_);
  or _50381_ (_42726_, _42724_, _37126_);
  and _50382_ (_42728_, _42726_, _42722_);
  not _50383_ (_42730_, _40223_);
  or _50384_ (_42732_, _42498_, _42730_);
  or _50385_ (_42734_, _42732_, _42728_);
  or _50386_ (_42736_, _42734_, _42718_);
  not _50387_ (_42738_, _40222_);
  or _50388_ (_42739_, _42459_, _42738_);
  and _50389_ (_42740_, _37811_, _36218_);
  or _50390_ (_42741_, _42740_, _42413_);
  or _50391_ (_42742_, _42741_, _42505_);
  or _50392_ (_42743_, _42742_, _42739_);
  or _50393_ (_42744_, _42493_, _42394_);
  or _50394_ (_42745_, _42744_, _42660_);
  or _50395_ (_42746_, _37519_, _42586_);
  or _50396_ (_42747_, _42746_, _42745_);
  or _50397_ (_42748_, _42747_, _42454_);
  or _50398_ (_42749_, _42748_, _42743_);
  or _50399_ (_42750_, _42749_, _42736_);
  and _50400_ (_42751_, _42750_, _42278_);
  or _50401_ (_30504_, _42751_, _42710_);
  or _50402_ (_42752_, _37349_, _36031_);
  or _50403_ (_42753_, _42477_, _42397_);
  or _50404_ (_42754_, _42753_, _42752_);
  or _50405_ (_42755_, _42754_, _42474_);
  or _50406_ (_42756_, _42755_, _42664_);
  and _50407_ (_42757_, _37126_, _35015_);
  or _50408_ (_42758_, _42740_, _42757_);
  or _50409_ (_42759_, _42716_, _42652_);
  or _50410_ (_42760_, _42759_, _42758_);
  or _50411_ (_42761_, _42481_, _40199_);
  or _50412_ (_42762_, _42761_, _42475_);
  or _50413_ (_42763_, _42762_, _36612_);
  not _50414_ (_42764_, _37464_);
  or _50415_ (_42765_, _42574_, _42764_);
  or _50416_ (_42766_, _42765_, _42763_);
  or _50417_ (_42767_, _42766_, _42760_);
  or _50418_ (_42768_, _42767_, _42756_);
  or _50419_ (_42769_, _37833_, _37888_);
  or _50420_ (_42770_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15507_);
  and _50421_ (_42771_, _42770_, _41755_);
  and _50422_ (_42772_, _42771_, _42769_);
  and _50423_ (_30506_, _42772_, _42768_);
  or _50424_ (_42773_, _37341_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _50425_ (_42774_, _42773_, _37833_);
  or _50426_ (_42775_, _42774_, _42647_);
  and _50427_ (_42776_, _35004_, _37268_);
  or _50428_ (_42777_, _42776_, _42596_);
  and _50429_ (_42778_, _42418_, _36306_);
  or _50430_ (_42779_, _42778_, _36590_);
  or _50431_ (_42780_, _42779_, _42777_);
  or _50432_ (_42781_, _42780_, _42775_);
  not _50433_ (_42782_, _37442_);
  nor _50434_ (_42783_, _42662_, _37453_);
  and _50435_ (_42784_, _42783_, _42782_);
  or _50436_ (_42785_, _42586_, _36448_);
  or _50437_ (_42786_, _42397_, _42785_);
  and _50438_ (_42787_, _35015_, _36383_);
  or _50439_ (_42788_, _42744_, _42787_);
  nor _50440_ (_42789_, _42788_, _42786_);
  nand _50441_ (_42790_, _42789_, _42784_);
  or _50442_ (_42791_, _42790_, _42781_);
  or _50443_ (_42792_, _42421_, _42414_);
  or _50444_ (_42793_, _42792_, _42791_);
  or _50445_ (_42794_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15507_);
  and _50446_ (_42795_, _42794_, _41755_);
  and _50447_ (_42796_, _42795_, _42769_);
  and _50448_ (_30508_, _42796_, _42793_);
  not _50449_ (_42797_, _42783_);
  or _50450_ (_42798_, _42797_, _42777_);
  or _50451_ (_42799_, _42798_, _42779_);
  or _50452_ (_42800_, _36448_, _36525_);
  nor _50453_ (_42801_, _42800_, _42714_);
  nand _50454_ (_42802_, _42801_, _40223_);
  or _50455_ (_42803_, _42741_, _42458_);
  or _50456_ (_42804_, _42803_, _42802_);
  or _50457_ (_42805_, _42465_, _42412_);
  or _50458_ (_42806_, _42805_, _42804_);
  or _50459_ (_42807_, _42806_, _42799_);
  and _50460_ (_42808_, _42807_, _33793_);
  and _50461_ (_42809_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _50462_ (_42810_, _37822_, _15507_);
  or _50463_ (_42811_, _42810_, _42809_);
  or _50464_ (_42812_, _42811_, _42808_);
  and _50465_ (_30510_, _42812_, _41755_);
  and _50466_ (_42813_, _42377_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor _50467_ (_42814_, _42385_, _37486_);
  nand _50468_ (_42816_, _42814_, _40222_);
  not _50469_ (_42817_, _34993_);
  or _50470_ (_42818_, _35015_, _42817_);
  and _50471_ (_42819_, _42818_, _37268_);
  or _50472_ (_42820_, _42819_, _42758_);
  or _50473_ (_42821_, _42820_, _42816_);
  or _50474_ (_42822_, _42732_, _42497_);
  or _50475_ (_42823_, _42822_, _42718_);
  or _50476_ (_42824_, _42823_, _42821_);
  and _50477_ (_42825_, _42824_, _42278_);
  or _50478_ (_30512_, _42825_, _42813_);
  nor _50479_ (_38759_, _35932_, rst);
  nor _50480_ (_38761_, _40215_, rst);
  and _50481_ (_42827_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _50482_ (_42828_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _50483_ (_42829_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _50484_ (_42830_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _50485_ (_42831_, _42830_, _42829_);
  and _50486_ (_42832_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _50487_ (_42833_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _50488_ (_42834_, _42833_, _42832_);
  and _50489_ (_42835_, _42834_, _42831_);
  and _50490_ (_42836_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _50491_ (_42837_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _50492_ (_42838_, _42837_, _42836_);
  and _50493_ (_42839_, _42838_, _42835_);
  nor _50494_ (_42840_, _42839_, _33870_);
  nor _50495_ (_42841_, _42840_, _42828_);
  nor _50496_ (_42842_, _42841_, _40199_);
  nor _50497_ (_42843_, _42842_, _42827_);
  nor _50498_ (_38762_, _42843_, rst);
  nor _50499_ (_38774_, _34185_, rst);
  and _50500_ (_38775_, _34447_, _41755_);
  nor _50501_ (_38776_, _34698_, rst);
  nor _50502_ (_38777_, _34938_, rst);
  and _50503_ (_38778_, _35213_, _41755_);
  nor _50504_ (_38779_, _35455_, rst);
  nor _50505_ (_38780_, _35701_, rst);
  nor _50506_ (_38781_, _40373_, rst);
  nor _50507_ (_38783_, _40551_, rst);
  nor _50508_ (_38784_, _40293_, rst);
  nor _50509_ (_38785_, _40335_, rst);
  nor _50510_ (_38786_, _40464_, rst);
  nor _50511_ (_38787_, _40270_, rst);
  nor _50512_ (_38789_, _40420_, rst);
  and _50513_ (_42844_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _50514_ (_42845_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _50515_ (_42846_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _50516_ (_42847_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _50517_ (_42848_, _42847_, _42846_);
  and _50518_ (_42849_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _50519_ (_42850_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _50520_ (_42851_, _42850_, _42849_);
  and _50521_ (_42852_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _50522_ (_42853_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _50523_ (_42854_, _42853_, _42852_);
  and _50524_ (_42855_, _42854_, _42851_);
  and _50525_ (_42856_, _42855_, _42848_);
  nor _50526_ (_42857_, _42856_, _33870_);
  nor _50527_ (_42858_, _42857_, _42845_);
  nor _50528_ (_42859_, _42858_, _40199_);
  nor _50529_ (_42860_, _42859_, _42844_);
  nor _50530_ (_38790_, _42860_, rst);
  and _50531_ (_42861_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _50532_ (_42862_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _50533_ (_42863_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _50534_ (_42864_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _50535_ (_42865_, _42864_, _42863_);
  and _50536_ (_42866_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _50537_ (_42867_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _50538_ (_42868_, _42867_, _42866_);
  and _50539_ (_42869_, _42868_, _42865_);
  and _50540_ (_42870_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _50541_ (_42871_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _50542_ (_42872_, _42871_, _42870_);
  and _50543_ (_42873_, _42872_, _42869_);
  nor _50544_ (_42874_, _42873_, _33870_);
  nor _50545_ (_42875_, _42874_, _42862_);
  nor _50546_ (_42876_, _42875_, _40199_);
  nor _50547_ (_42877_, _42876_, _42861_);
  nor _50548_ (_38791_, _42877_, rst);
  and _50549_ (_42878_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _50550_ (_42879_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _50551_ (_42880_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _50552_ (_42881_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _50553_ (_42882_, _42881_, _42880_);
  and _50554_ (_42883_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _50555_ (_42884_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _50556_ (_42885_, _42884_, _42883_);
  and _50557_ (_42886_, _42885_, _42882_);
  and _50558_ (_42887_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _50559_ (_42888_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _50560_ (_42889_, _42888_, _42887_);
  and _50561_ (_42890_, _42889_, _42886_);
  nor _50562_ (_42891_, _42890_, _33870_);
  nor _50563_ (_42892_, _42891_, _42879_);
  nor _50564_ (_42893_, _42892_, _40199_);
  nor _50565_ (_42894_, _42893_, _42878_);
  nor _50566_ (_38792_, _42894_, rst);
  and _50567_ (_42895_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _50568_ (_42896_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _50569_ (_42897_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _50570_ (_42898_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _50571_ (_42899_, _42898_, _42897_);
  and _50572_ (_42900_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _50573_ (_42901_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _50574_ (_42902_, _42901_, _42900_);
  and _50575_ (_42903_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _50576_ (_42904_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _50577_ (_42905_, _42904_, _42903_);
  and _50578_ (_42906_, _42905_, _42902_);
  and _50579_ (_42907_, _42906_, _42899_);
  nor _50580_ (_42908_, _42907_, _33870_);
  nor _50581_ (_42909_, _42908_, _42896_);
  nor _50582_ (_42910_, _42909_, _40199_);
  nor _50583_ (_42911_, _42910_, _42895_);
  nor _50584_ (_38793_, _42911_, rst);
  and _50585_ (_42912_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _50586_ (_42913_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _50587_ (_42914_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _50588_ (_42915_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _50589_ (_42916_, _42915_, _42914_);
  and _50590_ (_42917_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _50591_ (_42918_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _50592_ (_42919_, _42918_, _42917_);
  and _50593_ (_42920_, _42919_, _42916_);
  and _50594_ (_42921_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _50595_ (_42922_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _50596_ (_42923_, _42922_, _42921_);
  and _50597_ (_42924_, _42923_, _42920_);
  nor _50598_ (_42925_, _42924_, _33870_);
  nor _50599_ (_42926_, _42925_, _42913_);
  nor _50600_ (_42927_, _42926_, _40199_);
  nor _50601_ (_42928_, _42927_, _42912_);
  nor _50602_ (_38795_, _42928_, rst);
  and _50603_ (_42929_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _50604_ (_42930_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _50605_ (_42931_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _50606_ (_42932_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _50607_ (_42933_, _42932_, _42931_);
  and _50608_ (_42934_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _50609_ (_42935_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _50610_ (_42936_, _42935_, _42934_);
  and _50611_ (_42937_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _50612_ (_42938_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _50613_ (_42939_, _42938_, _42937_);
  and _50614_ (_42940_, _42939_, _42936_);
  and _50615_ (_42941_, _42940_, _42933_);
  nor _50616_ (_42942_, _42941_, _33870_);
  nor _50617_ (_42943_, _42942_, _42930_);
  nor _50618_ (_42944_, _42943_, _40199_);
  nor _50619_ (_42945_, _42944_, _42929_);
  nor _50620_ (_38796_, _42945_, rst);
  and _50621_ (_42946_, _40199_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _50622_ (_42947_, _33870_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _50623_ (_42948_, _34088_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _50624_ (_42949_, _33957_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _50625_ (_42950_, _42949_, _42948_);
  and _50626_ (_42951_, _34022_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _50627_ (_42952_, _33913_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _50628_ (_42953_, _42952_, _42951_);
  and _50629_ (_42954_, _42953_, _42950_);
  and _50630_ (_42955_, _34000_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _50631_ (_42956_, _34055_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _50632_ (_42957_, _42956_, _42955_);
  and _50633_ (_42958_, _42957_, _42954_);
  nor _50634_ (_42959_, _42958_, _33870_);
  nor _50635_ (_42960_, _42959_, _42947_);
  nor _50636_ (_42961_, _42960_, _40199_);
  nor _50637_ (_42962_, _42961_, _42946_);
  nor _50638_ (_38797_, _42962_, rst);
  and _50639_ (_42963_, _33804_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _50640_ (_42964_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _50641_ (_42965_, _42963_, _38515_);
  and _50642_ (_42966_, _42965_, _41755_);
  and _50643_ (_38821_, _42966_, _42964_);
  not _50644_ (_42967_, _42963_);
  or _50645_ (_42968_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _50646_ (_00000_, _42963_, _41755_);
  and _50647_ (_42969_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _41755_);
  or _50648_ (_42970_, _42969_, _00000_);
  and _50649_ (_38823_, _42970_, _42968_);
  nor _50650_ (_38859_, _40220_, rst);
  nor _50651_ (_38861_, _40468_, rst);
  nor _50652_ (_38862_, _40195_, rst);
  nor _50653_ (_42971_, _40220_, _24778_);
  and _50654_ (_42972_, _40220_, _24778_);
  nor _50655_ (_42973_, _42972_, _42971_);
  nor _50656_ (_42974_, _40357_, _24931_);
  and _50657_ (_42975_, _40357_, _24931_);
  nor _50658_ (_42976_, _42975_, _42974_);
  nor _50659_ (_42977_, _40492_, _25105_);
  and _50660_ (_42978_, _40492_, _25105_);
  nor _50661_ (_42979_, _42978_, _42977_);
  nor _50662_ (_42980_, _42979_, _42976_);
  nor _50663_ (_42981_, _40274_, _24626_);
  and _50664_ (_42982_, _40274_, _24626_);
  nor _50665_ (_42983_, _42982_, _42981_);
  nor _50666_ (_42984_, _40439_, _24494_);
  and _50667_ (_42985_, _40439_, _24494_);
  nor _50668_ (_42986_, _42985_, _42984_);
  nor _50669_ (_42987_, _42986_, _42983_);
  nand _50670_ (_42988_, _42987_, _42980_);
  nor _50671_ (_42989_, _42988_, _42973_);
  nor _50672_ (_42990_, _37169_, _42401_);
  and _50673_ (_42991_, _38764_, _27918_);
  and _50674_ (_42992_, _42991_, _42990_);
  and _50675_ (_42993_, _42992_, _42989_);
  and _50676_ (_42994_, _30064_, _28706_);
  nand _50677_ (_42995_, _42994_, _30732_);
  nor _50678_ (_42996_, _42995_, _31496_);
  and _50679_ (_42997_, _42996_, _32291_);
  and _50680_ (_42998_, _42997_, _26722_);
  nor _50681_ (_42999_, _42990_, _37646_);
  and _50682_ (_43000_, _42999_, _42998_);
  and _50683_ (_43001_, _43000_, _33042_);
  and _50684_ (_43002_, _43001_, _26908_);
  and _50685_ (_43003_, _42990_, _25845_);
  not _50686_ (_43004_, _37646_);
  nor _50687_ (_43005_, _42990_, _35510_);
  nor _50688_ (_43006_, _43005_, _43004_);
  and _50689_ (_43007_, _43006_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _50690_ (_43008_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _50691_ (_43009_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _50692_ (_43010_, _43009_, _43008_);
  nor _50693_ (_43011_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _50694_ (_43012_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _50695_ (_43013_, _43012_, _43011_);
  and _50696_ (_43014_, _43013_, _43010_);
  and _50697_ (_43015_, _43014_, _36722_);
  or _50698_ (_43016_, _43015_, _43007_);
  or _50699_ (_43017_, _43016_, _43003_);
  nor _50700_ (_43018_, _43017_, _43002_);
  nor _50701_ (_43019_, _42645_, _37318_);
  nor _50702_ (_43020_, _42612_, _42452_);
  nand _50703_ (_43021_, _43020_, _43019_);
  or _50704_ (_43022_, _37126_, _36108_);
  or _50705_ (_43023_, _43022_, _36579_);
  and _50706_ (_43024_, _43023_, _36174_);
  or _50707_ (_43025_, _43024_, _43021_);
  and _50708_ (_43026_, _43025_, _43018_);
  nand _50709_ (_43027_, _37635_, _35257_);
  and _50710_ (_43028_, _43027_, _37701_);
  nor _50711_ (_43029_, _43028_, _43018_);
  or _50712_ (_43030_, _42382_, _42650_);
  or _50713_ (_43031_, _43030_, _43029_);
  or _50714_ (_43032_, _43031_, _43026_);
  and _50715_ (_43033_, _43032_, _36700_);
  and _50716_ (_43034_, _36361_, _36514_);
  nor _50717_ (_43035_, _43034_, _42439_);
  nor _50718_ (_43036_, _43035_, _33750_);
  nor _50719_ (_43037_, _43036_, _36733_);
  not _50720_ (_43038_, _43037_);
  nor _50721_ (_43039_, _43038_, _43033_);
  nor _50722_ (_43040_, _38763_, _38788_);
  and _50723_ (_43041_, _43040_, _38806_);
  not _50724_ (_43042_, _43041_);
  and _50725_ (_43043_, _43042_, _43006_);
  not _50726_ (_43044_, _39022_);
  and _50727_ (_43045_, _43044_, _36722_);
  nor _50728_ (_43046_, _43045_, _43043_);
  not _50729_ (_43047_, _43046_);
  nor _50730_ (_43048_, _43047_, _43039_);
  not _50731_ (_43049_, _43048_);
  nor _50732_ (_43050_, _43049_, _42993_);
  nor _50733_ (_43051_, _40393_, _29802_);
  and _50734_ (_43052_, _40393_, _29802_);
  nor _50735_ (_43053_, _40313_, _24018_);
  and _50736_ (_43054_, _40313_, _24018_);
  nor _50737_ (_43055_, _43054_, _43053_);
  or _50738_ (_43056_, _43055_, _43052_);
  nor _50739_ (_43057_, _43056_, _43051_);
  nor _50740_ (_43058_, _40558_, _24138_);
  and _50741_ (_43059_, _40558_, _24138_);
  nor _50742_ (_43060_, _43059_, _43058_);
  nor _50743_ (_43061_, _43060_, _27907_);
  and _50744_ (_43062_, _43061_, _42989_);
  and _50745_ (_43063_, _43062_, _43057_);
  nor _50746_ (_43064_, _24778_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _50747_ (_43065_, _43064_, _43063_);
  not _50748_ (_43066_, _43065_);
  and _50749_ (_43067_, _43066_, _43050_);
  and _50750_ (_43068_, _43067_, _37624_);
  and _50751_ (_38866_, _43068_, _41755_);
  and _50752_ (_38867_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _41755_);
  and _50753_ (_38868_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _41755_);
  not _50754_ (_43069_, _42843_);
  and _50755_ (_43070_, _42611_, _37169_);
  and _50756_ (_43071_, _43070_, _43019_);
  nor _50757_ (_43072_, _43071_, _37657_);
  not _50758_ (_43073_, _43072_);
  and _50759_ (_43074_, _43034_, _37888_);
  and _50760_ (_43075_, _37104_, _37888_);
  nor _50761_ (_43076_, _43075_, _43074_);
  and _50762_ (_43077_, _43076_, _37624_);
  and _50763_ (_43078_, _43077_, _43073_);
  nor _50764_ (_43079_, _43078_, _43069_);
  and _50765_ (_43080_, _43078_, _40215_);
  nor _50766_ (_43081_, _43080_, _43079_);
  and _50767_ (_43083_, _43081_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _50768_ (_43084_, _43081_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _50769_ (_43085_, _42962_);
  nor _50770_ (_43086_, _43078_, _43085_);
  and _50771_ (_43087_, _43078_, _40420_);
  nor _50772_ (_43089_, _43087_, _43086_);
  and _50773_ (_43090_, _43089_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _50774_ (_43091_, _43089_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _50775_ (_43092_, _43091_, _43090_);
  not _50776_ (_43093_, _42945_);
  nor _50777_ (_43095_, _43078_, _43093_);
  and _50778_ (_43096_, _43078_, _40270_);
  nor _50779_ (_43097_, _43096_, _43095_);
  and _50780_ (_43098_, _43097_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _50781_ (_43099_, _43097_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not _50782_ (_43101_, _42928_);
  nor _50783_ (_43102_, _43078_, _43101_);
  and _50784_ (_43103_, _43078_, _40464_);
  nor _50785_ (_43104_, _43103_, _43102_);
  nand _50786_ (_43105_, _43104_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not _50787_ (_43107_, _42911_);
  nor _50788_ (_43108_, _43078_, _43107_);
  and _50789_ (_43109_, _43078_, _40335_);
  nor _50790_ (_43110_, _43109_, _43108_);
  and _50791_ (_43111_, _43110_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _50792_ (_43113_, _43110_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _50793_ (_43114_, _42894_);
  nor _50794_ (_43115_, _43078_, _43114_);
  and _50795_ (_43116_, _43078_, _40293_);
  nor _50796_ (_43117_, _43116_, _43115_);
  and _50797_ (_43119_, _43117_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _50798_ (_43120_, _42877_);
  nor _50799_ (_43122_, _43078_, _43120_);
  and _50800_ (_43123_, _43078_, _40551_);
  nor _50801_ (_43124_, _43123_, _43122_);
  and _50802_ (_43125_, _43124_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _50803_ (_43126_, _42860_);
  nor _50804_ (_43127_, _43078_, _43126_);
  and _50805_ (_43128_, _43078_, _40373_);
  nor _50806_ (_43130_, _43128_, _43127_);
  and _50807_ (_43131_, _43130_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _50808_ (_43132_, _43124_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _50809_ (_43134_, _43132_, _43125_);
  and _50810_ (_43135_, _43134_, _43131_);
  nor _50811_ (_43136_, _43135_, _43125_);
  not _50812_ (_43138_, _43136_);
  nor _50813_ (_43139_, _43117_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _50814_ (_43140_, _43139_, _43119_);
  and _50815_ (_43142_, _43140_, _43138_);
  nor _50816_ (_43143_, _43142_, _43119_);
  nor _50817_ (_43144_, _43143_, _43113_);
  or _50818_ (_43146_, _43144_, _43111_);
  or _50819_ (_43147_, _43104_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _50820_ (_43148_, _43147_, _43105_);
  nand _50821_ (_43150_, _43148_, _43146_);
  and _50822_ (_43151_, _43150_, _43105_);
  nor _50823_ (_43152_, _43151_, _43099_);
  or _50824_ (_43154_, _43152_, _43098_);
  and _50825_ (_43155_, _43154_, _43092_);
  nor _50826_ (_43157_, _43155_, _43090_);
  nor _50827_ (_43158_, _43157_, _43084_);
  or _50828_ (_43159_, _43158_, _43083_);
  and _50829_ (_43160_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _50830_ (_43161_, _43160_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _50831_ (_43162_, _43161_, _43159_);
  and _50832_ (_43163_, _43162_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _50833_ (_43165_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _50834_ (_43166_, _43165_, _43163_);
  nor _50835_ (_43167_, _43166_, _43081_);
  not _50836_ (_43169_, _43081_);
  nor _50837_ (_43170_, _43159_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _50838_ (_43171_, _43170_, _38493_);
  and _50839_ (_43173_, _43171_, _38498_);
  and _50840_ (_43174_, _43173_, _38483_);
  nor _50841_ (_43175_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _50842_ (_43177_, _43175_, _43174_);
  nor _50843_ (_43178_, _43177_, _43169_);
  nor _50844_ (_43179_, _43178_, _43167_);
  or _50845_ (_43181_, _43081_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _50846_ (_43182_, _43081_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _50847_ (_43183_, _43182_, _43181_);
  and _50848_ (_43185_, _43183_, _43179_);
  nand _50849_ (_43186_, _43185_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _50850_ (_43187_, _43185_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _50851_ (_43189_, _36700_, _42650_);
  nor _50852_ (_43190_, _43189_, _43036_);
  not _50853_ (_43192_, _43190_);
  and _50854_ (_43193_, _43192_, _43078_);
  or _50855_ (_43197_, _37635_, _37180_);
  or _50856_ (_43202_, _43030_, _43197_);
  or _50857_ (_43215_, _43202_, _43021_);
  and _50858_ (_43220_, _43215_, _36700_);
  nor _50859_ (_43221_, _43220_, _43075_);
  nor _50860_ (_43235_, _43221_, _43193_);
  and _50861_ (_43240_, _43235_, _43187_);
  and _50862_ (_43241_, _43240_, _43186_);
  and _50863_ (_43253_, _36744_, _27852_);
  not _50864_ (_43260_, _43189_);
  nor _50865_ (_43261_, _43260_, _38526_);
  and _50866_ (_43271_, _43221_, _43193_);
  and _50867_ (_43280_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _50868_ (_43281_, _43280_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _50869_ (_43289_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _50870_ (_43298_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _50871_ (_43299_, _43298_, _43289_);
  and _50872_ (_43308_, _43299_, _43281_);
  and _50873_ (_43316_, _43308_, _43161_);
  and _50874_ (_43317_, _43316_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _50875_ (_43325_, _43317_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _50876_ (_43332_, _43325_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _50877_ (_43333_, _43332_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _50878_ (_43348_, _43333_, _38515_);
  or _50879_ (_43349_, _43333_, _38515_);
  and _50880_ (_43354_, _43349_, _43348_);
  and _50881_ (_43362_, _43354_, _43271_);
  and _50882_ (_43368_, _43074_, _40216_);
  and _50883_ (_43372_, _43190_, _43078_);
  and _50884_ (_43386_, _43372_, _43221_);
  and _50885_ (_43391_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _50886_ (_43392_, _43391_, _43368_);
  or _50887_ (_43404_, _43392_, _43362_);
  nor _50888_ (_43411_, _43404_, _43261_);
  nand _50889_ (_43412_, _43411_, _43067_);
  or _50890_ (_43422_, _43412_, _43253_);
  or _50891_ (_43431_, _43422_, _43241_);
  not _50892_ (_43432_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _50893_ (_43433_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _50894_ (_43435_, _43433_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _50895_ (_43436_, _43435_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _50896_ (_43437_, _43436_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _50897_ (_43439_, _43437_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _50898_ (_43440_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _50899_ (_43441_, _43440_, _43439_);
  and _50900_ (_43443_, _43441_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _50901_ (_43444_, _43443_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _50902_ (_43445_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _50903_ (_43447_, _34077_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _50904_ (_43448_, _43447_, _40199_);
  nor _50905_ (_43450_, _43448_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _50906_ (_43451_, _43450_);
  and _50907_ (_43452_, _43451_, _43445_);
  and _50908_ (_43453_, _43452_, _43444_);
  nand _50909_ (_43455_, _43453_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _50910_ (_43456_, _43455_, _43432_);
  or _50911_ (_43457_, _43455_, _43432_);
  and _50912_ (_43459_, _43457_, _43456_);
  or _50913_ (_43460_, _43459_, _43067_);
  and _50914_ (_43461_, _43460_, _41755_);
  and _50915_ (_38870_, _43461_, _43431_);
  and _50916_ (_43463_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _41755_);
  and _50917_ (_43464_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _50918_ (_43466_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _50919_ (_43467_, _33793_, _43466_);
  not _50920_ (_43468_, _43467_);
  not _50921_ (_43470_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _50922_ (_43471_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _50923_ (_43472_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not _50924_ (_43474_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _50925_ (_43475_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _50926_ (_43476_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _50927_ (_43478_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _50928_ (_43479_, _43478_, _43476_);
  and _50929_ (_43481_, _43479_, _43475_);
  and _50930_ (_43482_, _43481_, _43474_);
  nor _50931_ (_43483_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _50932_ (_43484_, _43483_, _43482_);
  and _50933_ (_43486_, _43484_, _43472_);
  and _50934_ (_43487_, _43486_, _43471_);
  nor _50935_ (_43488_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _50936_ (_43490_, _43488_, _43487_);
  and _50937_ (_43491_, _43490_, _43470_);
  nor _50938_ (_43492_, _43491_, _43432_);
  and _50939_ (_43494_, _43491_, _43432_);
  nor _50940_ (_43495_, _43494_, _43492_);
  nor _50941_ (_43496_, _43490_, _43470_);
  or _50942_ (_43498_, _43496_, _43491_);
  not _50943_ (_43499_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _50944_ (_43500_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _50945_ (_43502_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _50946_ (_43503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _50947_ (_43504_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _50948_ (_43506_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _50949_ (_43507_, _43506_, _43503_);
  and _50950_ (_43508_, _43507_, _43504_);
  nor _50951_ (_43510_, _43508_, _43503_);
  nor _50952_ (_43511_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _50953_ (_43513_, _43511_, _43502_);
  not _50954_ (_43514_, _43513_);
  nor _50955_ (_43515_, _43514_, _43510_);
  nor _50956_ (_43516_, _43515_, _43502_);
  not _50957_ (_43518_, _43516_);
  and _50958_ (_43519_, _43518_, _43487_);
  and _50959_ (_43520_, _43519_, _43500_);
  and _50960_ (_43522_, _43520_, _43499_);
  and _50961_ (_43523_, _43522_, _43498_);
  nor _50962_ (_43524_, _43522_, _43498_);
  or _50963_ (_43526_, _43524_, _43523_);
  not _50964_ (_43527_, _43526_);
  and _50965_ (_43528_, _43516_, _43490_);
  and _50966_ (_43530_, _43516_, _43487_);
  and _50967_ (_43531_, _43530_, _43500_);
  nor _50968_ (_43532_, _43531_, _43499_);
  nor _50969_ (_43534_, _43532_, _43528_);
  not _50970_ (_43535_, _43534_);
  nor _50971_ (_43536_, _43530_, _43500_);
  nor _50972_ (_43538_, _43536_, _43531_);
  not _50973_ (_43539_, _43538_);
  and _50974_ (_43540_, _43516_, _43484_);
  and _50975_ (_43542_, _43540_, _43472_);
  nor _50976_ (_43543_, _43542_, _43471_);
  nor _50977_ (_43545_, _43543_, _43530_);
  not _50978_ (_43546_, _43545_);
  nor _50979_ (_43547_, _43540_, _43472_);
  nor _50980_ (_43548_, _43547_, _43542_);
  not _50981_ (_43549_, _43548_);
  not _50982_ (_43550_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _50983_ (_43551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _50984_ (_43553_, _43516_, _43482_);
  and _50985_ (_43554_, _43553_, _43551_);
  nor _50986_ (_43555_, _43554_, _43550_);
  nor _50987_ (_43557_, _43555_, _43540_);
  not _50988_ (_43558_, _43557_);
  and _50989_ (_43559_, _43516_, _43481_);
  nor _50990_ (_43561_, _43559_, _43474_);
  nor _50991_ (_43562_, _43561_, _43553_);
  not _50992_ (_43563_, _43562_);
  and _50993_ (_43565_, _43516_, _43479_);
  nor _50994_ (_43566_, _43565_, _43475_);
  nor _50995_ (_43567_, _43566_, _43559_);
  not _50996_ (_43569_, _43567_);
  and _50997_ (_43570_, _43516_, _43478_);
  nor _50998_ (_43571_, _43570_, _43476_);
  nor _50999_ (_43573_, _43571_, _43565_);
  not _51000_ (_43574_, _43573_);
  not _51001_ (_43575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _51002_ (_43577_, _43516_, _43575_);
  nor _51003_ (_43578_, _43516_, _43575_);
  nor _51004_ (_43580_, _43578_, _43577_);
  not _51005_ (_43581_, _43580_);
  and _51006_ (_43582_, _42334_, _42302_);
  and _51007_ (_43583_, _43582_, _42320_);
  not _51008_ (_43585_, _43583_);
  or _51009_ (_43586_, _42347_, _42303_);
  and _51010_ (_43587_, _43586_, _42327_);
  and _51011_ (_43589_, _42302_, _42285_);
  nor _51012_ (_43590_, _42347_, _43589_);
  nor _51013_ (_43591_, _43590_, _34938_);
  nor _51014_ (_43593_, _43591_, _43587_);
  and _51015_ (_43594_, _43593_, _43585_);
  and _51016_ (_43595_, _42343_, _42287_);
  not _51017_ (_43597_, _43595_);
  nor _51018_ (_43598_, _42334_, _42326_);
  nor _51019_ (_43599_, _43598_, _43597_);
  not _51020_ (_43601_, _42327_);
  and _51021_ (_43602_, _42323_, _42292_);
  nor _51022_ (_43603_, _43602_, _42295_);
  nor _51023_ (_43605_, _43603_, _43601_);
  nor _51024_ (_43606_, _43605_, _43599_);
  not _51025_ (_43607_, _42334_);
  and _51026_ (_43609_, _42323_, _42294_);
  nor _51027_ (_43610_, _43609_, _42305_);
  nor _51028_ (_43612_, _43610_, _43607_);
  not _51029_ (_43613_, _42300_);
  nor _51030_ (_43614_, _42324_, _43589_);
  nor _51031_ (_43615_, _43614_, _43613_);
  nor _51032_ (_43617_, _43615_, _43612_);
  and _51033_ (_43618_, _43617_, _43606_);
  and _51034_ (_43619_, _43618_, _43594_);
  and _51035_ (_43621_, _42317_, _42305_);
  not _51036_ (_43622_, _43621_);
  and _51037_ (_43623_, _43622_, _42329_);
  and _51038_ (_43625_, _42317_, _42295_);
  nor _51039_ (_43626_, _43625_, _42334_);
  not _51040_ (_43627_, _42295_);
  nor _51041_ (_43629_, _42347_, _42325_);
  and _51042_ (_43630_, _43629_, _43627_);
  nor _51043_ (_43631_, _43630_, _43626_);
  not _51044_ (_43633_, _43631_);
  and _51045_ (_43634_, _43633_, _43623_);
  and _51046_ (_43635_, _43634_, _43619_);
  and _51047_ (_43637_, _42327_, _42305_);
  and _51048_ (_43638_, _43595_, _42348_);
  nor _51049_ (_43639_, _43638_, _43637_);
  and _51050_ (_43641_, _42318_, _42542_);
  and _51051_ (_43642_, _42343_, _42302_);
  or _51052_ (_43644_, _43642_, _42288_);
  and _51053_ (_43645_, _42333_, _42288_);
  or _51054_ (_43646_, _43645_, _42326_);
  and _51055_ (_43647_, _43646_, _43644_);
  nor _51056_ (_43649_, _43647_, _43641_);
  and _51057_ (_43650_, _43649_, _43639_);
  and _51058_ (_43651_, _42356_, _42312_);
  and _51059_ (_43653_, _42302_, _42354_);
  nor _51060_ (_43654_, _43653_, _42298_);
  and _51061_ (_43655_, _43654_, _43651_);
  and _51062_ (_43657_, _42317_, _42293_);
  and _51063_ (_43658_, _42323_, _42285_);
  nor _51064_ (_43659_, _43658_, _42290_);
  nor _51065_ (_43661_, _43659_, _43601_);
  nor _51066_ (_43662_, _43661_, _43657_);
  and _51067_ (_43663_, _43609_, _42327_);
  and _51068_ (_43665_, _42347_, _42317_);
  nor _51069_ (_43666_, _43665_, _43663_);
  and _51070_ (_43667_, _43666_, _43662_);
  and _51071_ (_43669_, _42303_, _42306_);
  and _51072_ (_43670_, _42308_, _34938_);
  and _51073_ (_43671_, _43670_, _42347_);
  nor _51074_ (_43673_, _43671_, _43669_);
  and _51075_ (_43674_, _42348_, _42295_);
  and _51076_ (_43676_, _42334_, _42303_);
  nor _51077_ (_43677_, _43676_, _43674_);
  and _51078_ (_43678_, _43677_, _43673_);
  not _51079_ (_43679_, _42336_);
  and _51080_ (_43680_, _42308_, _42302_);
  and _51081_ (_43682_, _43680_, _42357_);
  nor _51082_ (_43683_, _43682_, _42350_);
  and _51083_ (_43684_, _43683_, _43679_);
  and _51084_ (_43686_, _43684_, _43678_);
  and _51085_ (_43687_, _43686_, _43667_);
  and _51086_ (_43688_, _43687_, _43655_);
  and _51087_ (_43690_, _43688_, _43650_);
  and _51088_ (_43691_, _43690_, _43635_);
  nor _51089_ (_43692_, _43507_, _43504_);
  nor _51090_ (_43694_, _43692_, _43508_);
  not _51091_ (_43695_, _43694_);
  nor _51092_ (_43696_, _43695_, _43691_);
  not _51093_ (_43698_, _43696_);
  nand _51094_ (_43699_, _43639_, _43623_);
  or _51095_ (_43700_, _42336_, _42311_);
  or _51096_ (_43702_, _43700_, _43587_);
  and _51097_ (_43703_, _42300_, _42293_);
  or _51098_ (_43704_, _43674_, _43703_);
  and _51099_ (_43706_, _42348_, _42288_);
  and _51100_ (_43707_, _43642_, _42300_);
  or _51101_ (_43709_, _43707_, _43706_);
  or _51102_ (_43710_, _43709_, _43704_);
  or _51103_ (_43711_, _43710_, _43702_);
  or _51104_ (_43712_, _43711_, _43699_);
  nor _51105_ (_43714_, _43712_, _43691_);
  not _51106_ (_43715_, _43714_);
  nor _51107_ (_43716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _51108_ (_43718_, _43716_, _43504_);
  and _51109_ (_43719_, _43718_, _43715_);
  and _51110_ (_43720_, _43695_, _43691_);
  nor _51111_ (_43722_, _43720_, _43696_);
  nand _51112_ (_43723_, _43722_, _43719_);
  and _51113_ (_43724_, _43723_, _43698_);
  not _51114_ (_43726_, _43724_);
  and _51115_ (_43727_, _43514_, _43510_);
  nor _51116_ (_43728_, _43727_, _43515_);
  and _51117_ (_43730_, _43728_, _43726_);
  and _51118_ (_43731_, _43730_, _43581_);
  not _51119_ (_43732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _51120_ (_43734_, _43577_, _43732_);
  or _51121_ (_43735_, _43734_, _43570_);
  and _51122_ (_43736_, _43735_, _43731_);
  and _51123_ (_43738_, _43736_, _43574_);
  and _51124_ (_43739_, _43738_, _43569_);
  and _51125_ (_43741_, _43739_, _43563_);
  nor _51126_ (_43742_, _43553_, _43551_);
  or _51127_ (_43743_, _43742_, _43554_);
  and _51128_ (_43744_, _43743_, _43741_);
  and _51129_ (_43746_, _43744_, _43558_);
  and _51130_ (_43747_, _43746_, _43549_);
  and _51131_ (_43748_, _43747_, _43546_);
  and _51132_ (_43750_, _43748_, _43539_);
  and _51133_ (_43751_, _43750_, _43535_);
  and _51134_ (_43752_, _43751_, _43527_);
  or _51135_ (_43754_, _43752_, _43523_);
  nor _51136_ (_43755_, _43754_, _43495_);
  and _51137_ (_43756_, _43754_, _43495_);
  or _51138_ (_43758_, _43756_, _43755_);
  or _51139_ (_43759_, _43758_, _43468_);
  or _51140_ (_43760_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _51141_ (_43762_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _51142_ (_43763_, _43762_, _43760_);
  and _51143_ (_43764_, _43763_, _43759_);
  or _51144_ (_38871_, _43764_, _43464_);
  nor _51145_ (_43766_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _51146_ (_38872_, _43766_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _51147_ (_38873_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _41755_);
  nor _51148_ (_43768_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _51149_ (_43770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _51150_ (_43771_, _43770_, _43768_);
  nor _51151_ (_43772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _51152_ (_43773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _51153_ (_43775_, _43773_, _43772_);
  and _51154_ (_43776_, _43775_, _43771_);
  nor _51155_ (_43777_, _43776_, rst);
  and _51156_ (_43779_, \oc8051_top_1.oc8051_rom1.ea_int , _33760_);
  nand _51157_ (_43780_, _43779_, _33793_);
  and _51158_ (_43781_, _43780_, _38873_);
  or _51159_ (_38875_, _43781_, _43777_);
  and _51160_ (_43783_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _51161_ (_43784_, _43783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _51162_ (_38876_, _43784_, _41755_);
  nor _51163_ (_43786_, _43450_, _40199_);
  or _51164_ (_43787_, _43691_, _33935_);
  nor _51165_ (_43789_, _43714_, _33901_);
  nand _51166_ (_43790_, _43691_, _33935_);
  and _51167_ (_43791_, _43790_, _43787_);
  nand _51168_ (_43793_, _43791_, _43789_);
  and _51169_ (_43794_, _43793_, _43787_);
  nor _51170_ (_43795_, _43794_, _40199_);
  and _51171_ (_43797_, _43795_, _33880_);
  nor _51172_ (_43798_, _43795_, _33880_);
  nor _51173_ (_43799_, _43798_, _43797_);
  nor _51174_ (_43800_, _43799_, _43786_);
  and _51175_ (_43801_, _33946_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _51176_ (_43802_, _43801_, _43786_);
  and _51177_ (_43803_, _43802_, _43712_);
  or _51178_ (_43804_, _43803_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _51179_ (_43805_, _43804_, _43800_);
  and _51180_ (_38877_, _43805_, _41755_);
  nor _51181_ (_43806_, _35147_, _34382_);
  and _51182_ (_43807_, _35888_, _35657_);
  and _51183_ (_43808_, _43807_, _43806_);
  and _51184_ (_43809_, _33804_, _41755_);
  nand _51185_ (_43810_, _43809_, _34654_);
  nor _51186_ (_43811_, _43810_, _34895_);
  not _51187_ (_43812_, _34142_);
  and _51188_ (_43813_, _43812_, _35411_);
  and _51189_ (_43814_, _43813_, _43811_);
  and _51190_ (_38880_, _43814_, _43808_);
  nor _51191_ (_43815_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _51192_ (_43816_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _51193_ (_43817_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _51194_ (_38883_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _41755_);
  and _51195_ (_43818_, _38883_, _43817_);
  or _51196_ (_38882_, _43818_, _43816_);
  not _51197_ (_43819_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _51198_ (_43820_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _51199_ (_43821_, _43820_, _43819_);
  and _51200_ (_43822_, _43820_, _43819_);
  nor _51201_ (_43823_, _43822_, _43821_);
  not _51202_ (_43824_, _43823_);
  and _51203_ (_43825_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _51204_ (_43826_, _43825_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _51205_ (_43827_, _43825_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _51206_ (_43828_, _43827_, _43826_);
  or _51207_ (_43829_, _43828_, _43820_);
  and _51208_ (_43830_, _43829_, _43824_);
  nor _51209_ (_43831_, _43821_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _51210_ (_43832_, _43821_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _51211_ (_43833_, _43832_, _43831_);
  or _51212_ (_43834_, _43826_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _51213_ (_38885_, _43834_, _41755_);
  and _51214_ (_43835_, _38885_, _43833_);
  and _51215_ (_38884_, _43835_, _43830_);
  not _51216_ (_43836_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _51217_ (_43837_, _43450_, _43836_);
  and _51218_ (_43838_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _51219_ (_43839_, _43837_);
  and _51220_ (_43840_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _51221_ (_43841_, _43840_, _43838_);
  and _51222_ (_38886_, _43841_, _41755_);
  and _51223_ (_43842_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _51224_ (_43843_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _51225_ (_43844_, _43843_, _43842_);
  and _51226_ (_38887_, _43844_, _41755_);
  and _51227_ (_43845_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _51228_ (_43846_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _51229_ (_43847_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _43846_);
  and _51230_ (_43848_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _51231_ (_43849_, _43848_, _43845_);
  and _51232_ (_38889_, _43849_, _41755_);
  and _51233_ (_43850_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _51234_ (_43851_, _43850_, _43847_);
  and _51235_ (_38890_, _43851_, _41755_);
  or _51236_ (_43852_, _43846_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _51237_ (_38891_, _43852_, _41755_);
  not _51238_ (_43853_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _51239_ (_43854_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _51240_ (_43855_, _43854_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _51241_ (_43856_, _43846_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _51242_ (_43857_, _43856_, _41755_);
  and _51243_ (_38892_, _43857_, _43855_);
  or _51244_ (_43858_, _43846_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _51245_ (_38893_, _43858_, _41755_);
  nor _51246_ (_43859_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _51247_ (_43860_, _43859_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _51248_ (_43861_, _43860_, _41755_);
  and _51249_ (_43862_, _38883_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _51250_ (_38894_, _43862_, _43861_);
  and _51251_ (_43863_, _43836_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _51252_ (_43864_, _43863_, _43860_);
  and _51253_ (_38895_, _43864_, _41755_);
  nand _51254_ (_43865_, _43860_, _38526_);
  or _51255_ (_43866_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _51256_ (_43867_, _43866_, _41755_);
  and _51257_ (_38896_, _43867_, _43865_);
  and _51258_ (_38897_, _37943_, _40164_);
  or _51259_ (_43868_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _51260_ (_43869_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand _51261_ (_43870_, _42963_, _43869_);
  and _51262_ (_43871_, _43870_, _41755_);
  and _51263_ (_38933_, _43871_, _43868_);
  or _51264_ (_43872_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _51265_ (_43873_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _41755_);
  or _51266_ (_43874_, _43873_, _00000_);
  and _51267_ (_38934_, _43874_, _43872_);
  or _51268_ (_43875_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _51269_ (_43876_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _51270_ (_43877_, _42963_, _43876_);
  and _51271_ (_43878_, _43877_, _41755_);
  and _51272_ (_38935_, _43878_, _43875_);
  or _51273_ (_43879_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _51274_ (_43880_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _51275_ (_43881_, _42963_, _43880_);
  and _51276_ (_43882_, _43881_, _41755_);
  and _51277_ (_38937_, _43882_, _43879_);
  or _51278_ (_43883_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not _51279_ (_43884_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _51280_ (_43885_, _42963_, _43884_);
  and _51281_ (_43886_, _43885_, _41755_);
  and _51282_ (_38938_, _43886_, _43883_);
  or _51283_ (_43887_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _51284_ (_43888_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _51285_ (_43889_, _42963_, _43888_);
  and _51286_ (_43890_, _43889_, _41755_);
  and _51287_ (_38939_, _43890_, _43887_);
  or _51288_ (_43891_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _51289_ (_43892_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6], _41755_);
  or _51290_ (_43893_, _43892_, _00000_);
  and _51291_ (_38940_, _43893_, _43891_);
  or _51292_ (_43894_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _51293_ (_43895_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _51294_ (_43896_, _42963_, _43895_);
  and _51295_ (_43897_, _43896_, _41755_);
  and _51296_ (_38941_, _43897_, _43894_);
  or _51297_ (_43898_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _51298_ (_43899_, _42963_, _38487_);
  and _51299_ (_43900_, _43899_, _41755_);
  and _51300_ (_38942_, _43900_, _43898_);
  or _51301_ (_43901_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _51302_ (_43902_, _42963_, _38493_);
  and _51303_ (_43903_, _43902_, _41755_);
  and _51304_ (_38943_, _43903_, _43901_);
  or _51305_ (_43904_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _51306_ (_43905_, _42963_, _38498_);
  and _51307_ (_43906_, _43905_, _41755_);
  and _51308_ (_38944_, _43906_, _43904_);
  or _51309_ (_43907_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _51310_ (_43908_, _42963_, _38483_);
  and _51311_ (_43909_, _43908_, _41755_);
  and _51312_ (_38945_, _43909_, _43907_);
  or _51313_ (_43910_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _51314_ (_43911_, _42963_, _38504_);
  and _51315_ (_43912_, _43911_, _41755_);
  and _51316_ (_38946_, _43912_, _43910_);
  or _51317_ (_43913_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _51318_ (_43914_, _42963_, _38479_);
  and _51319_ (_43915_, _43914_, _41755_);
  and _51320_ (_38948_, _43915_, _43913_);
  or _51321_ (_43916_, _42963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _51322_ (_43917_, _42963_, _38510_);
  and _51323_ (_43918_, _43917_, _41755_);
  and _51324_ (_38949_, _43918_, _43916_);
  or _51325_ (_43919_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _51326_ (_43920_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _41755_);
  or _51327_ (_43921_, _43920_, _00000_);
  and _51328_ (_38953_, _43921_, _43919_);
  or _51329_ (_43922_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _51330_ (_43923_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _41755_);
  or _51331_ (_43924_, _43923_, _00000_);
  and _51332_ (_38954_, _43924_, _43922_);
  or _51333_ (_43925_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _51334_ (_43926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _41755_);
  or _51335_ (_43927_, _43926_, _00000_);
  and _51336_ (_38955_, _43927_, _43925_);
  or _51337_ (_43928_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _51338_ (_43929_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _41755_);
  or _51339_ (_43930_, _43929_, _00000_);
  and _51340_ (_38956_, _43930_, _43928_);
  or _51341_ (_43931_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _51342_ (_43932_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _41755_);
  or _51343_ (_43933_, _43932_, _00000_);
  and _51344_ (_38957_, _43933_, _43931_);
  or _51345_ (_43934_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _51346_ (_43935_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _41755_);
  or _51347_ (_43936_, _43935_, _00000_);
  and _51348_ (_38958_, _43936_, _43934_);
  or _51349_ (_43937_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _51350_ (_43938_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _41755_);
  or _51351_ (_43939_, _43938_, _00000_);
  and _51352_ (_38959_, _43939_, _43937_);
  or _51353_ (_43940_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _51354_ (_43941_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _41755_);
  or _51355_ (_43942_, _43941_, _00000_);
  and _51356_ (_38960_, _43942_, _43940_);
  or _51357_ (_43943_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _51358_ (_43944_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _41755_);
  or _51359_ (_43945_, _43944_, _00000_);
  and _51360_ (_38962_, _43945_, _43943_);
  or _51361_ (_43946_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _51362_ (_43947_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _41755_);
  or _51363_ (_43948_, _43947_, _00000_);
  and _51364_ (_38963_, _43948_, _43946_);
  or _51365_ (_43949_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _51366_ (_43950_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _41755_);
  or _51367_ (_43951_, _43950_, _00000_);
  and _51368_ (_38964_, _43951_, _43949_);
  or _51369_ (_43952_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _51370_ (_43953_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _41755_);
  or _51371_ (_43954_, _43953_, _00000_);
  and _51372_ (_38965_, _43954_, _43952_);
  or _51373_ (_43955_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _51374_ (_43956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _41755_);
  or _51375_ (_43957_, _43956_, _00000_);
  and _51376_ (_38966_, _43957_, _43955_);
  or _51377_ (_43958_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _51378_ (_43959_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _41755_);
  or _51379_ (_43960_, _43959_, _00000_);
  and _51380_ (_38967_, _43960_, _43958_);
  or _51381_ (_43961_, _42967_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _51382_ (_43962_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _41755_);
  or _51383_ (_43963_, _43962_, _00000_);
  and _51384_ (_38968_, _43963_, _43961_);
  and _51385_ (_43964_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _51386_ (_43965_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _51387_ (_43966_, _43965_, _43964_);
  and _51388_ (_39145_, _43966_, _41755_);
  and _51389_ (_43967_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _51390_ (_43968_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or _51391_ (_43969_, _43968_, _43967_);
  and _51392_ (_39146_, _43969_, _41755_);
  and _51393_ (_43970_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _51394_ (_43971_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _51395_ (_43972_, _43971_, _43970_);
  and _51396_ (_39147_, _43972_, _41755_);
  and _51397_ (_43973_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _51398_ (_43974_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or _51399_ (_43975_, _43974_, _43973_);
  and _51400_ (_39148_, _43975_, _41755_);
  and _51401_ (_43976_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _51402_ (_43977_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _51403_ (_43978_, _43977_, _43976_);
  and _51404_ (_39149_, _43978_, _41755_);
  and _51405_ (_43979_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _51406_ (_43980_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or _51407_ (_43981_, _43980_, _43979_);
  and _51408_ (_39150_, _43981_, _41755_);
  and _51409_ (_43982_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _51410_ (_43983_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or _51411_ (_43984_, _43983_, _43982_);
  and _51412_ (_39151_, _43984_, _41755_);
  and _51413_ (_43985_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _51414_ (_43986_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _51415_ (_43987_, _43986_, _43985_);
  and _51416_ (_39152_, _43987_, _41755_);
  and _51417_ (_43988_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _51418_ (_43989_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _51419_ (_43990_, _43989_, _43988_);
  and _51420_ (_39153_, _43990_, _41755_);
  and _51421_ (_43991_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _51422_ (_43992_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _51423_ (_43993_, _43992_, _43991_);
  and _51424_ (_39154_, _43993_, _41755_);
  and _51425_ (_43994_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _51426_ (_43995_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _51427_ (_43996_, _43995_, _43994_);
  and _51428_ (_39155_, _43996_, _41755_);
  and _51429_ (_43997_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _51430_ (_43998_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _51431_ (_43999_, _43998_, _43997_);
  and _51432_ (_39156_, _43999_, _41755_);
  and _51433_ (_44000_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _51434_ (_44001_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _51435_ (_44002_, _44001_, _44000_);
  and _51436_ (_39157_, _44002_, _41755_);
  and _51437_ (_44003_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _51438_ (_44004_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _51439_ (_44005_, _44004_, _44003_);
  and _51440_ (_39158_, _44005_, _41755_);
  and _51441_ (_44006_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _51442_ (_00006_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _51443_ (_00007_, _00006_, _44006_);
  and _51444_ (_39159_, _00007_, _41755_);
  and _51445_ (_00008_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _51446_ (_00009_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _51447_ (_00010_, _00009_, _00008_);
  and _51448_ (_39160_, _00010_, _41755_);
  and _51449_ (_00011_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _51450_ (_00012_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _51451_ (_00013_, _00012_, _00011_);
  and _51452_ (_39162_, _00013_, _41755_);
  and _51453_ (_00014_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _51454_ (_00015_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _51455_ (_00016_, _00015_, _00014_);
  and _51456_ (_39163_, _00016_, _41755_);
  and _51457_ (_00017_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _51458_ (_00018_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _51459_ (_00019_, _00018_, _00017_);
  and _51460_ (_39164_, _00019_, _41755_);
  and _51461_ (_00020_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _51462_ (_00021_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _51463_ (_00022_, _00021_, _00020_);
  and _51464_ (_39165_, _00022_, _41755_);
  and _51465_ (_00023_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _51466_ (_00024_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _51467_ (_00025_, _00024_, _00023_);
  and _51468_ (_39166_, _00025_, _41755_);
  and _51469_ (_00026_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _51470_ (_00027_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _51471_ (_00028_, _00027_, _00026_);
  and _51472_ (_39167_, _00028_, _41755_);
  and _51473_ (_00029_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _51474_ (_00030_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _51475_ (_00031_, _00030_, _00029_);
  and _51476_ (_39168_, _00031_, _41755_);
  and _51477_ (_00032_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _51478_ (_00033_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _51479_ (_00034_, _00033_, _00032_);
  and _51480_ (_39169_, _00034_, _41755_);
  and _51481_ (_00035_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _51482_ (_00036_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _51483_ (_00037_, _00036_, _00035_);
  and _51484_ (_39170_, _00037_, _41755_);
  and _51485_ (_00038_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _51486_ (_00039_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _51487_ (_00040_, _00039_, _00038_);
  and _51488_ (_39171_, _00040_, _41755_);
  and _51489_ (_00041_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _51490_ (_00042_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _51491_ (_00043_, _00042_, _00041_);
  and _51492_ (_39173_, _00043_, _41755_);
  and _51493_ (_00044_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _51494_ (_00045_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _51495_ (_00046_, _00045_, _00044_);
  and _51496_ (_39174_, _00046_, _41755_);
  and _51497_ (_00047_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _51498_ (_00048_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _51499_ (_00049_, _00048_, _00047_);
  and _51500_ (_39175_, _00049_, _41755_);
  and _51501_ (_00050_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _51502_ (_00051_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _51503_ (_00052_, _00051_, _00050_);
  and _51504_ (_39176_, _00052_, _41755_);
  and _51505_ (_00053_, _43837_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _51506_ (_00054_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _51507_ (_00055_, _00054_, _00053_);
  and _51508_ (_39177_, _00055_, _41755_);
  nor _51509_ (_39178_, _34229_, rst);
  nor _51510_ (_39179_, _34491_, rst);
  nor _51511_ (_39180_, _34742_, rst);
  nor _51512_ (_39181_, _40167_, rst);
  nor _51513_ (_39183_, _40385_, rst);
  nor _51514_ (_39184_, _40508_, rst);
  nor _51515_ (_39185_, _40309_, rst);
  nor _51516_ (_39186_, _40348_, rst);
  nor _51517_ (_39187_, _40482_, rst);
  nor _51518_ (_39189_, _40246_, rst);
  nor _51519_ (_39190_, _40434_, rst);
  and _51520_ (_39206_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _41755_);
  and _51521_ (_39207_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _41755_);
  and _51522_ (_39208_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _41755_);
  and _51523_ (_39210_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _41755_);
  and _51524_ (_39211_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _41755_);
  and _51525_ (_39212_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _41755_);
  and _51526_ (_39213_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _41755_);
  nor _51527_ (_00056_, _43386_, _43189_);
  nor _51528_ (_00057_, _00056_, _29046_);
  and _51529_ (_00058_, _43074_, _43126_);
  and _51530_ (_00059_, _43271_, _40374_);
  or _51531_ (_00060_, _00059_, _00058_);
  and _51532_ (_00061_, _37613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _51533_ (_00062_, _00061_, _00060_);
  or _51534_ (_00063_, _00062_, _00057_);
  and _51535_ (_00064_, _36174_, _37888_);
  and _51536_ (_00065_, _00064_, _36383_);
  nor _51537_ (_00066_, _43220_, _00065_);
  nor _51538_ (_00067_, _00066_, _43193_);
  nor _51539_ (_00068_, _43130_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _51540_ (_00069_, _00068_, _43131_);
  nand _51541_ (_00070_, _00069_, _00067_);
  nand _51542_ (_00071_, _00070_, _43067_);
  or _51543_ (_00072_, _00071_, _00063_);
  or _51544_ (_00073_, _43067_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _51545_ (_00074_, _00073_, _41755_);
  and _51546_ (_39214_, _00074_, _00072_);
  not _51547_ (_00075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _51548_ (_00076_, _43068_, _00075_);
  and _51549_ (_00077_, _43074_, _43120_);
  and _51550_ (_00078_, _43271_, _40552_);
  or _51551_ (_00079_, _00078_, _00077_);
  or _51552_ (_00080_, _43134_, _43131_);
  not _51553_ (_00081_, _00067_);
  nor _51554_ (_00082_, _00081_, _43135_);
  and _51555_ (_00083_, _00082_, _00080_);
  or _51556_ (_00084_, _00083_, _00079_);
  nor _51557_ (_00085_, _00056_, _29714_);
  or _51558_ (_00086_, _00085_, _00084_);
  and _51559_ (_00087_, _00086_, _43067_);
  or _51560_ (_00088_, _00087_, _00076_);
  and _51561_ (_39215_, _00088_, _41755_);
  nor _51562_ (_00089_, _00056_, _30404_);
  and _51563_ (_00090_, _43271_, _40294_);
  and _51564_ (_00091_, _43074_, _43114_);
  and _51565_ (_00092_, _36744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _51566_ (_00093_, _00092_, _00091_);
  or _51567_ (_00094_, _00093_, _00090_);
  or _51568_ (_00095_, _00094_, _00089_);
  nor _51569_ (_00096_, _43140_, _43138_);
  nor _51570_ (_00097_, _00096_, _43142_);
  nand _51571_ (_00098_, _00097_, _00067_);
  nand _51572_ (_00099_, _00098_, _43067_);
  or _51573_ (_00100_, _00099_, _00095_);
  not _51574_ (_00101_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _51575_ (_00102_, _43450_, _00101_);
  and _51576_ (_00103_, _43450_, _00101_);
  nor _51577_ (_00104_, _00103_, _00102_);
  or _51578_ (_00105_, _00104_, _43067_);
  and _51579_ (_00106_, _00105_, _41755_);
  and _51580_ (_39216_, _00106_, _00100_);
  nor _51581_ (_00107_, _00056_, _31213_);
  or _51582_ (_00108_, _43113_, _43111_);
  or _51583_ (_00109_, _00108_, _43143_);
  nand _51584_ (_00110_, _00108_, _43143_);
  and _51585_ (_00111_, _00110_, _43235_);
  nand _51586_ (_00112_, _00111_, _00109_);
  and _51587_ (_00113_, _43271_, _40336_);
  and _51588_ (_00114_, _43074_, _43107_);
  and _51589_ (_00115_, _36744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _51590_ (_00116_, _00115_, _00114_);
  nor _51591_ (_00117_, _00116_, _00113_);
  and _51592_ (_00118_, _00117_, _00112_);
  nand _51593_ (_00119_, _00118_, _43067_);
  or _51594_ (_00120_, _00119_, _00107_);
  and _51595_ (_00121_, _00102_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _51596_ (_00122_, _00102_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _51597_ (_00123_, _00122_, _00121_);
  or _51598_ (_00124_, _00123_, _43067_);
  and _51599_ (_00125_, _00124_, _41755_);
  and _51600_ (_39217_, _00125_, _00120_);
  nor _51601_ (_00126_, _00056_, _31997_);
  and _51602_ (_00127_, _43271_, _40465_);
  and _51603_ (_00128_, _43074_, _43101_);
  and _51604_ (_00129_, _36744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _51605_ (_00130_, _00129_, _00128_);
  or _51606_ (_00131_, _00130_, _00127_);
  or _51607_ (_00132_, _43148_, _43146_);
  and _51608_ (_00133_, _43235_, _43150_);
  and _51609_ (_00134_, _00133_, _00132_);
  nor _51610_ (_00135_, _00134_, _00131_);
  nand _51611_ (_00136_, _00135_, _43067_);
  or _51612_ (_00137_, _00136_, _00126_);
  and _51613_ (_00138_, _43435_, _43451_);
  nor _51614_ (_00139_, _00121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _51615_ (_00140_, _00139_, _00138_);
  or _51616_ (_00141_, _00140_, _43067_);
  and _51617_ (_00142_, _00141_, _41755_);
  and _51618_ (_39218_, _00142_, _00137_);
  nor _51619_ (_00143_, _00056_, _32814_);
  or _51620_ (_00144_, _43099_, _43098_);
  or _51621_ (_00145_, _00144_, _43151_);
  nand _51622_ (_00146_, _00144_, _43151_);
  and _51623_ (_00147_, _00146_, _43235_);
  nand _51624_ (_00148_, _00147_, _00145_);
  and _51625_ (_00149_, _43271_, _40271_);
  and _51626_ (_00150_, _43074_, _43093_);
  and _51627_ (_00151_, _36744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _51628_ (_00152_, _00151_, _00150_);
  nor _51629_ (_00153_, _00152_, _00149_);
  and _51630_ (_00154_, _00153_, _00148_);
  nand _51631_ (_00155_, _00154_, _43067_);
  or _51632_ (_00156_, _00155_, _00143_);
  and _51633_ (_00157_, _43436_, _43451_);
  nor _51634_ (_00158_, _00138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _51635_ (_00159_, _00158_, _00157_);
  or _51636_ (_00160_, _00159_, _43067_);
  and _51637_ (_00161_, _00160_, _41755_);
  and _51638_ (_39219_, _00161_, _00156_);
  nor _51639_ (_00162_, _00056_, _33533_);
  and _51640_ (_00163_, _43271_, _40421_);
  and _51641_ (_00164_, _43074_, _43085_);
  and _51642_ (_00165_, _36744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _51643_ (_00166_, _00165_, _00164_);
  or _51644_ (_00167_, _00166_, _00163_);
  nor _51645_ (_00168_, _43154_, _43092_);
  nor _51646_ (_00169_, _00168_, _43155_);
  and _51647_ (_00170_, _00169_, _00067_);
  nor _51648_ (_00171_, _00170_, _00167_);
  nand _51649_ (_00172_, _00171_, _43067_);
  or _51650_ (_00173_, _00172_, _00162_);
  and _51651_ (_00174_, _00157_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _51652_ (_00175_, _00157_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _51653_ (_00176_, _00175_, _00174_);
  or _51654_ (_00177_, _00176_, _43067_);
  and _51655_ (_00178_, _00177_, _41755_);
  and _51656_ (_39221_, _00178_, _00173_);
  or _51657_ (_00179_, _43083_, _43084_);
  nor _51658_ (_00180_, _00179_, _43157_);
  and _51659_ (_00181_, _00179_, _43157_);
  or _51660_ (_00182_, _00181_, _00180_);
  or _51661_ (_00183_, _00182_, _00081_);
  or _51662_ (_00184_, _00056_, _27841_);
  nand _51663_ (_00185_, _43271_, _40216_);
  nand _51664_ (_00186_, _43074_, _43069_);
  nand _51665_ (_00187_, _36744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _51666_ (_00188_, _00187_, _00186_);
  and _51667_ (_00189_, _00188_, _00185_);
  and _51668_ (_00190_, _00189_, _00184_);
  and _51669_ (_00191_, _00190_, _00183_);
  nand _51670_ (_00192_, _00191_, _43067_);
  and _51671_ (_00193_, _00174_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _51672_ (_00194_, _00174_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _51673_ (_00195_, _00194_, _00193_);
  or _51674_ (_00196_, _00195_, _43067_);
  and _51675_ (_00197_, _00196_, _41755_);
  and _51676_ (_39222_, _00197_, _00192_);
  and _51677_ (_00198_, _36744_, _29057_);
  nor _51678_ (_00199_, _43260_, _38560_);
  and _51679_ (_00200_, _43159_, _38487_);
  nor _51680_ (_00201_, _43159_, _38487_);
  nor _51681_ (_00202_, _00201_, _00200_);
  or _51682_ (_00203_, _00202_, _43169_);
  nand _51683_ (_00204_, _00202_, _43169_);
  and _51684_ (_00205_, _00204_, _43235_);
  and _51685_ (_00206_, _00205_, _00203_);
  and _51686_ (_00207_, _43074_, _40374_);
  and _51687_ (_00208_, _43271_, _42291_);
  or _51688_ (_00209_, _00208_, _00207_);
  and _51689_ (_00210_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _51690_ (_00211_, _00210_, _00209_);
  nand _51691_ (_00212_, _00211_, _43067_);
  or _51692_ (_00213_, _00212_, _00206_);
  or _51693_ (_00214_, _00213_, _00199_);
  or _51694_ (_00215_, _00214_, _00198_);
  and _51695_ (_00216_, _00193_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _51696_ (_00217_, _00193_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _51697_ (_00218_, _00217_, _00216_);
  or _51698_ (_00219_, _00218_, _43067_);
  and _51699_ (_00220_, _00219_, _41755_);
  and _51700_ (_39223_, _00220_, _00215_);
  and _51701_ (_00221_, _43159_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _51702_ (_00222_, _00221_, _43169_);
  and _51703_ (_00223_, _43170_, _43081_);
  nor _51704_ (_00224_, _00223_, _00222_);
  nand _51705_ (_00225_, _00224_, _38493_);
  or _51706_ (_00226_, _00224_, _38493_);
  and _51707_ (_00227_, _00226_, _43235_);
  and _51708_ (_00228_, _00227_, _00225_);
  nor _51709_ (_00229_, _43260_, _38589_);
  and _51710_ (_00230_, _43074_, _40552_);
  and _51711_ (_00231_, _43271_, _42286_);
  or _51712_ (_00232_, _00231_, _00230_);
  and _51713_ (_00233_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _51714_ (_00234_, _00233_, _00232_);
  nor _51715_ (_00235_, _00234_, _00229_);
  nand _51716_ (_00236_, _00235_, _43067_);
  or _51717_ (_00237_, _00236_, _00228_);
  nor _51718_ (_00238_, _37624_, _29714_);
  or _51719_ (_00239_, _00238_, _00237_);
  and _51720_ (_00240_, _43441_, _43451_);
  nor _51721_ (_00241_, _00216_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _51722_ (_00242_, _00241_, _00240_);
  or _51723_ (_00243_, _00242_, _43067_);
  and _51724_ (_00244_, _00243_, _41755_);
  and _51725_ (_39224_, _00244_, _00239_);
  not _51726_ (_00245_, _43067_);
  nor _51727_ (_00246_, _37624_, _30404_);
  nor _51728_ (_00247_, _43260_, _38617_);
  and _51729_ (_00248_, _43074_, _40294_);
  and _51730_ (_00249_, _43271_, _42301_);
  or _51731_ (_00250_, _00249_, _00248_);
  and _51732_ (_00251_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _51733_ (_00252_, _00251_, _00250_);
  or _51734_ (_00253_, _00252_, _00247_);
  and _51735_ (_00254_, _43171_, _43081_);
  and _51736_ (_00255_, _00222_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _51737_ (_00256_, _00255_, _00254_);
  nand _51738_ (_00257_, _00256_, _38498_);
  or _51739_ (_00258_, _00256_, _38498_);
  and _51740_ (_00259_, _00258_, _00257_);
  and _51741_ (_00260_, _00259_, _00067_);
  or _51742_ (_00261_, _00260_, _00253_);
  or _51743_ (_00262_, _00261_, _00246_);
  or _51744_ (_00263_, _00262_, _00245_);
  and _51745_ (_00264_, _00240_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _51746_ (_00265_, _00240_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _51747_ (_00266_, _00265_, _00264_);
  or _51748_ (_00267_, _00266_, _43067_);
  and _51749_ (_00268_, _00267_, _41755_);
  and _51750_ (_39225_, _00268_, _00263_);
  nor _51751_ (_00269_, _37624_, _31213_);
  nor _51752_ (_00270_, _43260_, _38646_);
  nor _51753_ (_00271_, _43316_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _51754_ (_00272_, _00271_, _43317_);
  and _51755_ (_00273_, _00272_, _43271_);
  and _51756_ (_00274_, _43074_, _40336_);
  or _51757_ (_00275_, _00274_, _00273_);
  and _51758_ (_00276_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _51759_ (_00277_, _00276_, _00275_);
  or _51760_ (_00278_, _00277_, _00270_);
  and _51761_ (_00279_, _43162_, _43169_);
  and _51762_ (_00280_, _43173_, _43081_);
  nor _51763_ (_00281_, _00280_, _00279_);
  nor _51764_ (_00282_, _00281_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _51765_ (_00283_, _00281_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _51766_ (_00284_, _00283_, _00282_);
  and _51767_ (_00285_, _00284_, _00067_);
  or _51768_ (_00286_, _00285_, _00278_);
  or _51769_ (_00287_, _00286_, _00269_);
  or _51770_ (_00288_, _00287_, _00245_);
  and _51771_ (_00289_, _00264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _51772_ (_00290_, _00264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _51773_ (_00291_, _00290_, _00289_);
  or _51774_ (_00292_, _00291_, _43067_);
  and _51775_ (_00293_, _00292_, _41755_);
  and _51776_ (_39226_, _00293_, _00288_);
  nor _51777_ (_00294_, _43317_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _51778_ (_00295_, _00294_, _43325_);
  nand _51779_ (_00296_, _00295_, _43271_);
  and _51780_ (_00297_, _43163_, _43169_);
  and _51781_ (_00298_, _43174_, _43081_);
  nor _51782_ (_00299_, _00298_, _00297_);
  nor _51783_ (_00300_, _00299_, _38504_);
  and _51784_ (_00301_, _00299_, _38504_);
  or _51785_ (_00302_, _00301_, _00081_);
  or _51786_ (_00303_, _00302_, _00300_);
  or _51787_ (_00304_, _37624_, _31997_);
  or _51788_ (_00305_, _43260_, _38675_);
  nand _51789_ (_00306_, _43074_, _40465_);
  nand _51790_ (_00307_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _51791_ (_00308_, _00307_, _00306_);
  and _51792_ (_00309_, _00308_, _00305_);
  and _51793_ (_00310_, _00309_, _00304_);
  and _51794_ (_00311_, _00310_, _00303_);
  and _51795_ (_00312_, _00311_, _00296_);
  nand _51796_ (_00313_, _00312_, _43067_);
  and _51797_ (_00314_, _00289_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _51798_ (_00315_, _00289_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _51799_ (_00316_, _00315_, _00314_);
  or _51800_ (_00317_, _00316_, _43067_);
  and _51801_ (_00318_, _00317_, _41755_);
  and _51802_ (_39227_, _00318_, _00313_);
  and _51803_ (_00319_, _36744_, _32825_);
  and _51804_ (_00320_, _00297_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _51805_ (_00321_, _00298_, _38504_);
  nor _51806_ (_00322_, _00321_, _00320_);
  nand _51807_ (_00323_, _00322_, _38479_);
  or _51808_ (_00324_, _00322_, _38479_);
  and _51809_ (_00325_, _00324_, _43235_);
  and _51810_ (_00326_, _00325_, _00323_);
  nor _51811_ (_00327_, _43260_, _38705_);
  nor _51812_ (_00328_, _43325_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _51813_ (_00329_, _00328_, _43332_);
  and _51814_ (_00330_, _00329_, _43271_);
  and _51815_ (_00331_, _43074_, _40271_);
  and _51816_ (_00332_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _51817_ (_00333_, _00332_, _00331_);
  or _51818_ (_00334_, _00333_, _00330_);
  nor _51819_ (_00335_, _00334_, _00327_);
  nand _51820_ (_00336_, _00335_, _43067_);
  or _51821_ (_00337_, _00336_, _00326_);
  or _51822_ (_00338_, _00337_, _00319_);
  or _51823_ (_00339_, _00314_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand _51824_ (_00340_, _00314_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _51825_ (_00341_, _00340_, _00339_);
  or _51826_ (_00342_, _00341_, _43067_);
  and _51827_ (_00343_, _00342_, _41755_);
  and _51828_ (_39228_, _00343_, _00338_);
  or _51829_ (_00344_, _43332_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _51830_ (_00345_, _00344_, _43333_);
  nand _51831_ (_00346_, _00345_, _43271_);
  or _51832_ (_00347_, _37624_, _33533_);
  or _51833_ (_00348_, _43260_, _38732_);
  nand _51834_ (_00349_, _43074_, _40421_);
  nand _51835_ (_00350_, _43386_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _51836_ (_00351_, _00350_, _00349_);
  and _51837_ (_00352_, _00351_, _00348_);
  and _51838_ (_00353_, _00352_, _00347_);
  nor _51839_ (_00354_, _43179_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _51840_ (_00355_, _43179_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _51841_ (_00356_, _00355_, _00081_);
  or _51842_ (_00357_, _00356_, _00354_);
  and _51843_ (_00358_, _00357_, _00353_);
  and _51844_ (_00359_, _00358_, _00346_);
  nand _51845_ (_00360_, _00359_, _43067_);
  or _51846_ (_00361_, _43453_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _51847_ (_00362_, _00361_, _43455_);
  or _51848_ (_00363_, _00362_, _43067_);
  and _51849_ (_00364_, _00363_, _41755_);
  and _51850_ (_39229_, _00364_, _00360_);
  and _51851_ (_00365_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _51852_ (_00366_, _43718_, _43715_);
  nor _51853_ (_00367_, _00366_, _43719_);
  or _51854_ (_00368_, _00367_, _43468_);
  or _51855_ (_00369_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _51856_ (_00370_, _00369_, _43762_);
  and _51857_ (_00371_, _00370_, _00368_);
  or _51858_ (_39230_, _00371_, _00365_);
  or _51859_ (_00372_, _43722_, _43719_);
  and _51860_ (_00373_, _00372_, _43723_);
  or _51861_ (_00374_, _00373_, _43468_);
  or _51862_ (_00375_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _51863_ (_00376_, _00375_, _43762_);
  and _51864_ (_00377_, _00376_, _00374_);
  and _51865_ (_00378_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _51866_ (_39232_, _00378_, _00377_);
  and _51867_ (_00379_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _51868_ (_00380_, _43728_, _43726_);
  nor _51869_ (_00381_, _00380_, _43730_);
  or _51870_ (_00382_, _00381_, _43468_);
  or _51871_ (_00383_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _51872_ (_00384_, _00383_, _43762_);
  and _51873_ (_00385_, _00384_, _00382_);
  or _51874_ (_39233_, _00385_, _00379_);
  and _51875_ (_00386_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _51876_ (_00387_, _43730_, _43581_);
  nor _51877_ (_00388_, _00387_, _43731_);
  or _51878_ (_00389_, _00388_, _43468_);
  or _51879_ (_00390_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _51880_ (_00391_, _00390_, _43762_);
  and _51881_ (_00392_, _00391_, _00389_);
  or _51882_ (_39234_, _00392_, _00386_);
  and _51883_ (_00393_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _51884_ (_00394_, _43735_, _43731_);
  nor _51885_ (_00395_, _00394_, _43736_);
  or _51886_ (_00396_, _00395_, _43468_);
  or _51887_ (_00397_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _51888_ (_00398_, _00397_, _43762_);
  and _51889_ (_00399_, _00398_, _00396_);
  or _51890_ (_39235_, _00399_, _00393_);
  nor _51891_ (_00400_, _43736_, _43574_);
  nor _51892_ (_00401_, _00400_, _43738_);
  or _51893_ (_00402_, _00401_, _43468_);
  or _51894_ (_00403_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _51895_ (_00404_, _00403_, _43762_);
  and _51896_ (_00405_, _00404_, _00402_);
  and _51897_ (_00406_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _51898_ (_39236_, _00406_, _00405_);
  nor _51899_ (_00407_, _43738_, _43569_);
  nor _51900_ (_00408_, _00407_, _43739_);
  or _51901_ (_00409_, _00408_, _43468_);
  or _51902_ (_00410_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _51903_ (_00411_, _00410_, _43762_);
  and _51904_ (_00412_, _00411_, _00409_);
  and _51905_ (_00413_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _51906_ (_39237_, _00413_, _00412_);
  and _51907_ (_00414_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _51908_ (_00415_, _43739_, _43563_);
  nor _51909_ (_00416_, _00415_, _43741_);
  or _51910_ (_00417_, _00416_, _43468_);
  or _51911_ (_00418_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _51912_ (_00419_, _00418_, _43762_);
  and _51913_ (_00420_, _00419_, _00417_);
  or _51914_ (_39238_, _00420_, _00414_);
  nor _51915_ (_00421_, _43743_, _43741_);
  nor _51916_ (_00422_, _00421_, _43744_);
  or _51917_ (_00423_, _00422_, _43468_);
  or _51918_ (_00424_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _51919_ (_00425_, _00424_, _43762_);
  and _51920_ (_00426_, _00425_, _00423_);
  and _51921_ (_00427_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _51922_ (_39239_, _00427_, _00426_);
  nor _51923_ (_00428_, _43744_, _43558_);
  nor _51924_ (_00429_, _00428_, _43746_);
  or _51925_ (_00430_, _00429_, _43468_);
  or _51926_ (_00431_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _51927_ (_00432_, _00431_, _43762_);
  and _51928_ (_00433_, _00432_, _00430_);
  and _51929_ (_00434_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or _51930_ (_39240_, _00434_, _00433_);
  nor _51931_ (_00435_, _43746_, _43549_);
  nor _51932_ (_00436_, _00435_, _43747_);
  or _51933_ (_00437_, _00436_, _43468_);
  or _51934_ (_00438_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _51935_ (_00439_, _00438_, _43762_);
  and _51936_ (_00440_, _00439_, _00437_);
  and _51937_ (_00441_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _51938_ (_39241_, _00441_, _00440_);
  nor _51939_ (_00442_, _43747_, _43546_);
  nor _51940_ (_00443_, _00442_, _43748_);
  or _51941_ (_00444_, _00443_, _43468_);
  or _51942_ (_00445_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _51943_ (_00446_, _00445_, _43762_);
  and _51944_ (_00447_, _00446_, _00444_);
  and _51945_ (_00448_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _51946_ (_39243_, _00448_, _00447_);
  nor _51947_ (_00449_, _43748_, _43539_);
  nor _51948_ (_00450_, _00449_, _43750_);
  or _51949_ (_00451_, _00450_, _43468_);
  or _51950_ (_00452_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _51951_ (_00453_, _00452_, _43762_);
  and _51952_ (_00454_, _00453_, _00451_);
  and _51953_ (_00455_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _51954_ (_39244_, _00455_, _00454_);
  nor _51955_ (_00456_, _43750_, _43535_);
  nor _51956_ (_00457_, _00456_, _43751_);
  or _51957_ (_00458_, _00457_, _43468_);
  or _51958_ (_00459_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _51959_ (_00460_, _00459_, _43762_);
  and _51960_ (_00461_, _00460_, _00458_);
  and _51961_ (_00462_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _51962_ (_39245_, _00462_, _00461_);
  and _51963_ (_00463_, _43463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _51964_ (_00464_, _43751_, _43527_);
  nor _51965_ (_00465_, _00464_, _43752_);
  or _51966_ (_00466_, _00465_, _43468_);
  or _51967_ (_00467_, _43467_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _51968_ (_00468_, _00467_, _43762_);
  and _51969_ (_00469_, _00468_, _00466_);
  or _51970_ (_39246_, _00469_, _00463_);
  and _51971_ (_00470_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _51972_ (_00471_, _00470_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _51973_ (_39247_, _00471_, _41755_);
  and _51974_ (_00472_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _51975_ (_00473_, _00472_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _51976_ (_39248_, _00473_, _41755_);
  and _51977_ (_00474_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _51978_ (_00475_, _00474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _51979_ (_39249_, _00475_, _41755_);
  and _51980_ (_00476_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _51981_ (_00477_, _00476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _51982_ (_39250_, _00477_, _41755_);
  and _51983_ (_00478_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _51984_ (_00479_, _00478_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _51985_ (_39251_, _00479_, _41755_);
  and _51986_ (_00480_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _51987_ (_00481_, _00480_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _51988_ (_39252_, _00481_, _41755_);
  and _51989_ (_00482_, _43776_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _51990_ (_00483_, _00482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _51991_ (_39254_, _00483_, _41755_);
  nor _51992_ (_00484_, _43714_, _40199_);
  nand _51993_ (_00485_, _00484_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _51994_ (_00486_, _00484_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _51995_ (_00487_, _00486_, _43762_);
  and _51996_ (_39255_, _00487_, _00485_);
  or _51997_ (_00488_, _43791_, _43789_);
  and _51998_ (_00489_, _00488_, _43793_);
  or _51999_ (_00490_, _00489_, _40199_);
  or _52000_ (_00491_, _33793_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _52001_ (_00492_, _00491_, _43762_);
  and _52002_ (_39256_, _00492_, _00490_);
  and _52003_ (_00493_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _52004_ (_00494_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _52005_ (_00495_, _00494_, _38883_);
  or _52006_ (_39272_, _00495_, _00493_);
  and _52007_ (_00496_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _52008_ (_00497_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _52009_ (_00498_, _00497_, _38883_);
  or _52010_ (_39273_, _00498_, _00496_);
  and _52011_ (_00499_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _52012_ (_00500_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _52013_ (_00501_, _00500_, _38883_);
  or _52014_ (_39274_, _00501_, _00499_);
  and _52015_ (_00502_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _52016_ (_00503_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _52017_ (_00504_, _00503_, _38883_);
  or _52018_ (_39275_, _00504_, _00502_);
  and _52019_ (_00505_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _52020_ (_00506_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _52021_ (_00507_, _00506_, _38883_);
  or _52022_ (_39276_, _00507_, _00505_);
  and _52023_ (_00508_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _52024_ (_00509_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _52025_ (_00510_, _00509_, _38883_);
  or _52026_ (_39277_, _00510_, _00508_);
  and _52027_ (_00511_, _43815_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _52028_ (_00512_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _52029_ (_00513_, _00512_, _38883_);
  or _52030_ (_39278_, _00513_, _00511_);
  and _52031_ (_39279_, _43823_, _41755_);
  nor _52032_ (_39280_, _43833_, rst);
  and _52033_ (_39281_, _43829_, _41755_);
  and _52034_ (_00514_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _52035_ (_00515_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or _52036_ (_00516_, _00515_, _00514_);
  and _52037_ (_39282_, _00516_, _41755_);
  and _52038_ (_00517_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _52039_ (_00518_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _52040_ (_00519_, _00518_, _00517_);
  and _52041_ (_39283_, _00519_, _41755_);
  and _52042_ (_00520_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _52043_ (_00521_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or _52044_ (_00522_, _00521_, _00520_);
  and _52045_ (_39284_, _00522_, _41755_);
  and _52046_ (_00523_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _52047_ (_00524_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or _52048_ (_00525_, _00524_, _00523_);
  and _52049_ (_39286_, _00525_, _41755_);
  and _52050_ (_00526_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _52051_ (_00527_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or _52052_ (_00528_, _00527_, _00526_);
  and _52053_ (_39287_, _00528_, _41755_);
  and _52054_ (_00529_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _52055_ (_00530_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or _52056_ (_00531_, _00530_, _00529_);
  and _52057_ (_39288_, _00531_, _41755_);
  and _52058_ (_00532_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _52059_ (_00533_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or _52060_ (_00534_, _00533_, _00532_);
  and _52061_ (_39289_, _00534_, _41755_);
  and _52062_ (_00535_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _52063_ (_00536_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or _52064_ (_00537_, _00536_, _00535_);
  and _52065_ (_39290_, _00537_, _41755_);
  and _52066_ (_00538_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _52067_ (_00539_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _52068_ (_00540_, _00539_, _00538_);
  and _52069_ (_39291_, _00540_, _41755_);
  and _52070_ (_00541_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _52071_ (_00542_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _52072_ (_00543_, _00542_, _00541_);
  and _52073_ (_39292_, _00543_, _41755_);
  and _52074_ (_00544_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _52075_ (_00545_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _52076_ (_00546_, _00545_, _00544_);
  and _52077_ (_39293_, _00546_, _41755_);
  and _52078_ (_00547_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _52079_ (_00548_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _52080_ (_00549_, _00548_, _00547_);
  and _52081_ (_39294_, _00549_, _41755_);
  and _52082_ (_00550_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _52083_ (_00551_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _52084_ (_00552_, _00551_, _00550_);
  and _52085_ (_39295_, _00552_, _41755_);
  and _52086_ (_00553_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _52087_ (_00554_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _52088_ (_00555_, _00554_, _00553_);
  and _52089_ (_39297_, _00555_, _41755_);
  and _52090_ (_00556_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _52091_ (_00557_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _52092_ (_00558_, _00557_, _00556_);
  and _52093_ (_39298_, _00558_, _41755_);
  and _52094_ (_00559_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _52095_ (_00560_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _52096_ (_00561_, _00560_, _00559_);
  and _52097_ (_39299_, _00561_, _41755_);
  and _52098_ (_00562_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _52099_ (_00563_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _52100_ (_00564_, _00563_, _00562_);
  and _52101_ (_39300_, _00564_, _41755_);
  and _52102_ (_00565_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _52103_ (_00566_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _52104_ (_00567_, _00566_, _00565_);
  and _52105_ (_39301_, _00567_, _41755_);
  and _52106_ (_00568_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _52107_ (_00569_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _52108_ (_00570_, _00569_, _00568_);
  and _52109_ (_39302_, _00570_, _41755_);
  and _52110_ (_00571_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _52111_ (_00572_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _52112_ (_00573_, _00572_, _00571_);
  and _52113_ (_39303_, _00573_, _41755_);
  and _52114_ (_00574_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _52115_ (_00575_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _52116_ (_00576_, _00575_, _00574_);
  and _52117_ (_39304_, _00576_, _41755_);
  and _52118_ (_00577_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _52119_ (_00578_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _52120_ (_00579_, _00578_, _00577_);
  and _52121_ (_39305_, _00579_, _41755_);
  and _52122_ (_00580_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _52123_ (_00581_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _52124_ (_00582_, _00581_, _00580_);
  and _52125_ (_39306_, _00582_, _41755_);
  and _52126_ (_00583_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _52127_ (_00584_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _52128_ (_00585_, _00584_, _00583_);
  and _52129_ (_39308_, _00585_, _41755_);
  and _52130_ (_00586_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _52131_ (_00587_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _52132_ (_00588_, _00587_, _00586_);
  and _52133_ (_39309_, _00588_, _41755_);
  and _52134_ (_00589_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _52135_ (_00590_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _52136_ (_00591_, _00590_, _00589_);
  and _52137_ (_39310_, _00591_, _41755_);
  and _52138_ (_00592_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _52139_ (_00593_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _52140_ (_00594_, _00593_, _00592_);
  and _52141_ (_39311_, _00594_, _41755_);
  and _52142_ (_00595_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _52143_ (_00596_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _52144_ (_00597_, _00596_, _00595_);
  and _52145_ (_39312_, _00597_, _41755_);
  and _52146_ (_00598_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _52147_ (_00599_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _52148_ (_00600_, _00599_, _00598_);
  and _52149_ (_39313_, _00600_, _41755_);
  and _52150_ (_00601_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _52151_ (_00602_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _52152_ (_00603_, _00602_, _00601_);
  and _52153_ (_39314_, _00603_, _41755_);
  and _52154_ (_00604_, _43837_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _52155_ (_00605_, _43839_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _52156_ (_00606_, _00605_, _00604_);
  and _52157_ (_39315_, _00606_, _41755_);
  and _52158_ (_00607_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52159_ (_00608_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _52160_ (_00609_, _00608_, _00607_);
  and _52161_ (_39316_, _00609_, _41755_);
  and _52162_ (_00610_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52163_ (_00611_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _52164_ (_00612_, _00611_, _00610_);
  and _52165_ (_39317_, _00612_, _41755_);
  and _52166_ (_00613_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52167_ (_00614_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _52168_ (_00615_, _00614_, _00613_);
  and _52169_ (_39319_, _00615_, _41755_);
  and _52170_ (_00616_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52171_ (_00617_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _52172_ (_00618_, _00617_, _00616_);
  and _52173_ (_39320_, _00618_, _41755_);
  and _52174_ (_00619_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52175_ (_00620_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _52176_ (_00621_, _00620_, _00619_);
  and _52177_ (_39321_, _00621_, _41755_);
  and _52178_ (_00622_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52179_ (_00623_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _52180_ (_00624_, _00623_, _00622_);
  and _52181_ (_39322_, _00624_, _41755_);
  and _52182_ (_00625_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52183_ (_00626_, _43847_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _52184_ (_00627_, _00626_, _00625_);
  and _52185_ (_39323_, _00627_, _41755_);
  and _52186_ (_00628_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52187_ (_00629_, _40385_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52188_ (_00630_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _52189_ (_00631_, _00630_, _43846_);
  and _52190_ (_00632_, _00631_, _00629_);
  or _52191_ (_00633_, _00632_, _00628_);
  and _52192_ (_39324_, _00633_, _41755_);
  and _52193_ (_00634_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52194_ (_00635_, _40508_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52195_ (_00636_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _52196_ (_00637_, _00636_, _43846_);
  and _52197_ (_00638_, _00637_, _00635_);
  or _52198_ (_00639_, _00638_, _00634_);
  and _52199_ (_39325_, _00639_, _41755_);
  and _52200_ (_00640_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52201_ (_00641_, _40309_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52202_ (_00642_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _52203_ (_00643_, _00642_, _43846_);
  and _52204_ (_00644_, _00643_, _00641_);
  or _52205_ (_00645_, _00644_, _00640_);
  and _52206_ (_39326_, _00645_, _41755_);
  and _52207_ (_00646_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52208_ (_00647_, _40348_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52209_ (_00648_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _52210_ (_00649_, _00648_, _43846_);
  and _52211_ (_00650_, _00649_, _00647_);
  or _52212_ (_00651_, _00650_, _00646_);
  and _52213_ (_39327_, _00651_, _41755_);
  and _52214_ (_00652_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52215_ (_00653_, _40482_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52216_ (_00654_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _52217_ (_00655_, _00654_, _43846_);
  and _52218_ (_00656_, _00655_, _00653_);
  or _52219_ (_00657_, _00656_, _00652_);
  and _52220_ (_39328_, _00657_, _41755_);
  and _52221_ (_00658_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52222_ (_00659_, _40246_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52223_ (_00660_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _52224_ (_00661_, _00660_, _43846_);
  and _52225_ (_00662_, _00661_, _00659_);
  or _52226_ (_00663_, _00662_, _00658_);
  and _52227_ (_39330_, _00663_, _41755_);
  and _52228_ (_00664_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52229_ (_00665_, _40434_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52230_ (_00666_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _52231_ (_00667_, _00666_, _43846_);
  and _52232_ (_00668_, _00667_, _00665_);
  or _52233_ (_00669_, _00668_, _00664_);
  and _52234_ (_39331_, _00669_, _41755_);
  and _52235_ (_00670_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _52236_ (_00671_, _40195_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _52237_ (_00672_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _52238_ (_00673_, _00672_, _43846_);
  and _52239_ (_00674_, _00673_, _00671_);
  or _52240_ (_00675_, _00674_, _00670_);
  and _52241_ (_39332_, _00675_, _41755_);
  and _52242_ (_00676_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _52243_ (_00677_, _00676_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52244_ (_00678_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _43846_);
  and _52245_ (_00679_, _00678_, _41755_);
  and _52246_ (_39333_, _00679_, _00677_);
  and _52247_ (_00680_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _52248_ (_00681_, _00680_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52249_ (_00682_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _43846_);
  and _52250_ (_00683_, _00682_, _41755_);
  and _52251_ (_39334_, _00683_, _00681_);
  and _52252_ (_00684_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _52253_ (_00685_, _00684_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52254_ (_00686_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _43846_);
  and _52255_ (_00687_, _00686_, _41755_);
  and _52256_ (_39335_, _00687_, _00685_);
  and _52257_ (_00688_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _52258_ (_00689_, _00688_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52259_ (_00690_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _43846_);
  and _52260_ (_00691_, _00690_, _41755_);
  and _52261_ (_39336_, _00691_, _00689_);
  and _52262_ (_00692_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _52263_ (_00693_, _00692_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52264_ (_00694_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _43846_);
  and _52265_ (_00695_, _00694_, _41755_);
  and _52266_ (_39337_, _00695_, _00693_);
  and _52267_ (_00696_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _52268_ (_00697_, _00696_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52269_ (_00698_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _43846_);
  and _52270_ (_00699_, _00698_, _41755_);
  and _52271_ (_39338_, _00699_, _00697_);
  and _52272_ (_00700_, _43853_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _52273_ (_00701_, _00700_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52274_ (_00702_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _43846_);
  and _52275_ (_00703_, _00702_, _41755_);
  and _52276_ (_39339_, _00703_, _00701_);
  nand _52277_ (_00704_, _43860_, _29046_);
  or _52278_ (_00705_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _52279_ (_00706_, _00705_, _41755_);
  and _52280_ (_39341_, _00706_, _00704_);
  nand _52281_ (_00707_, _43860_, _29714_);
  or _52282_ (_00708_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _52283_ (_00709_, _00708_, _41755_);
  and _52284_ (_39342_, _00709_, _00707_);
  nand _52285_ (_00710_, _43860_, _30404_);
  or _52286_ (_00711_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _52287_ (_00712_, _00711_, _41755_);
  and _52288_ (_39343_, _00712_, _00710_);
  nand _52289_ (_00713_, _43860_, _31213_);
  or _52290_ (_00714_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _52291_ (_00715_, _00714_, _41755_);
  and _52292_ (_39344_, _00715_, _00713_);
  nand _52293_ (_00716_, _43860_, _31997_);
  or _52294_ (_00717_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _52295_ (_00718_, _00717_, _41755_);
  and _52296_ (_39345_, _00718_, _00716_);
  nand _52297_ (_00719_, _43860_, _32814_);
  or _52298_ (_00720_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _52299_ (_00721_, _00720_, _41755_);
  and _52300_ (_39346_, _00721_, _00719_);
  nand _52301_ (_00722_, _43860_, _33533_);
  or _52302_ (_00723_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _52303_ (_00724_, _00723_, _41755_);
  and _52304_ (_39347_, _00724_, _00722_);
  nand _52305_ (_00725_, _43860_, _27841_);
  or _52306_ (_00726_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _52307_ (_00727_, _00726_, _41755_);
  and _52308_ (_39348_, _00727_, _00725_);
  nand _52309_ (_00728_, _43860_, _38560_);
  or _52310_ (_00729_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _52311_ (_00730_, _00729_, _41755_);
  and _52312_ (_39349_, _00730_, _00728_);
  nand _52313_ (_00731_, _43860_, _38589_);
  or _52314_ (_00732_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _52315_ (_00733_, _00732_, _41755_);
  and _52316_ (_39350_, _00733_, _00731_);
  nand _52317_ (_00734_, _43860_, _38617_);
  or _52318_ (_00735_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _52319_ (_00736_, _00735_, _41755_);
  and _52320_ (_39352_, _00736_, _00734_);
  nand _52321_ (_00737_, _43860_, _38646_);
  or _52322_ (_00738_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _52323_ (_00739_, _00738_, _41755_);
  and _52324_ (_39353_, _00739_, _00737_);
  nand _52325_ (_00740_, _43860_, _38675_);
  or _52326_ (_00741_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _52327_ (_00742_, _00741_, _41755_);
  and _52328_ (_39354_, _00742_, _00740_);
  nand _52329_ (_00743_, _43860_, _38705_);
  or _52330_ (_00744_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _52331_ (_00745_, _00744_, _41755_);
  and _52332_ (_39355_, _00745_, _00743_);
  nand _52333_ (_00746_, _43860_, _38732_);
  or _52334_ (_00747_, _43860_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _52335_ (_00748_, _00747_, _41755_);
  and _52336_ (_39356_, _00748_, _00746_);
  nor _52337_ (_39563_, _40232_, rst);
  nor _52338_ (_00749_, _40439_, _40220_);
  nor _52339_ (_00750_, _40358_, _40492_);
  and _52340_ (_00751_, _00750_, _40274_);
  and _52341_ (_00752_, _00751_, _00749_);
  not _52342_ (_00753_, _40313_);
  nor _52343_ (_00754_, _39035_, _39019_);
  and _52344_ (_00755_, _39035_, _39019_);
  nor _52345_ (_00756_, _00755_, _00754_);
  and _52346_ (_00757_, _39008_, _38996_);
  nor _52347_ (_00758_, _39008_, _38996_);
  or _52348_ (_00759_, _00758_, _00757_);
  nor _52349_ (_00760_, _00759_, _00756_);
  and _52350_ (_00761_, _00759_, _00756_);
  nor _52351_ (_00762_, _00761_, _00760_);
  nor _52352_ (_00763_, _39057_, _39046_);
  and _52353_ (_00764_, _39057_, _39046_);
  nor _52354_ (_00765_, _00764_, _00763_);
  not _52355_ (_00766_, _38985_);
  nor _52356_ (_00767_, _39068_, _00766_);
  and _52357_ (_00768_, _39068_, _00766_);
  nor _52358_ (_00769_, _00768_, _00767_);
  nor _52359_ (_00770_, _00769_, _00765_);
  and _52360_ (_00771_, _00769_, _00765_);
  or _52361_ (_00772_, _00771_, _00770_);
  or _52362_ (_00773_, _00772_, _00762_);
  nand _52363_ (_00774_, _00772_, _00762_);
  and _52364_ (_00775_, _00774_, _00773_);
  or _52365_ (_00776_, _00775_, _00753_);
  and _52366_ (_00777_, _40393_, _40558_);
  or _52367_ (_00778_, _40313_, _38901_);
  and _52368_ (_00779_, _00778_, _00777_);
  and _52369_ (_00780_, _00779_, _00776_);
  nor _52370_ (_00781_, _40393_, _40558_);
  and _52371_ (_00782_, _00781_, _00753_);
  and _52372_ (_00783_, _00782_, _38805_);
  not _52373_ (_00784_, _40393_);
  and _52374_ (_00785_, _00784_, _40558_);
  or _52375_ (_00786_, _00753_, _38813_);
  or _52376_ (_00787_, _40313_, _38908_);
  and _52377_ (_00788_, _00787_, _00786_);
  and _52378_ (_00789_, _00788_, _00785_);
  and _52379_ (_00790_, _00781_, _40313_);
  and _52380_ (_00791_, _00790_, _38858_);
  or _52381_ (_00792_, _00791_, _00789_);
  or _52382_ (_00793_, _00792_, _00783_);
  or _52383_ (_00794_, _00753_, _38850_);
  nor _52384_ (_00795_, _00784_, _40558_);
  or _52385_ (_00796_, _40313_, _38926_);
  and _52386_ (_00797_, _00796_, _00795_);
  and _52387_ (_00798_, _00797_, _00794_);
  or _52388_ (_00799_, _00798_, _00793_);
  or _52389_ (_00800_, _00799_, _00780_);
  and _52390_ (_00801_, _00800_, _00752_);
  nor _52391_ (_00802_, _42482_, _37497_);
  and _52392_ (_00803_, _36295_, _36262_);
  nor _52393_ (_00804_, _00803_, _36590_);
  and _52394_ (_00805_, _00804_, _00802_);
  and _52395_ (_00806_, _36306_, _36459_);
  or _52396_ (_00807_, _00806_, _37027_);
  or _52397_ (_00808_, _00807_, _37398_);
  nor _52398_ (_00809_, _00808_, _42485_);
  and _52399_ (_00810_, _00809_, _00805_);
  and _52400_ (_00811_, _42784_, _42417_);
  and _52401_ (_00812_, _00811_, _00810_);
  and _52402_ (_00813_, _00812_, _37387_);
  nor _52403_ (_00814_, _00813_, _33750_);
  and _52404_ (_00815_, _42967_, p0in_reg[0]);
  and _52405_ (_00816_, _42963_, p0_in[0]);
  or _52406_ (_00817_, _00816_, _00815_);
  or _52407_ (_00818_, _00817_, _00814_);
  nand _52408_ (_00819_, _00814_, _39133_);
  and _52409_ (_00820_, _00819_, _00818_);
  and _52410_ (_00821_, _00820_, _00777_);
  or _52411_ (_00822_, _00821_, _00753_);
  and _52412_ (_00823_, _42967_, p0in_reg[3]);
  and _52413_ (_00824_, _42963_, p0_in[3]);
  or _52414_ (_00825_, _00824_, _00823_);
  or _52415_ (_00826_, _00825_, _00814_);
  nand _52416_ (_00827_, _00814_, _39365_);
  and _52417_ (_00828_, _00827_, _00826_);
  and _52418_ (_00829_, _00828_, _00781_);
  and _52419_ (_00830_, _42967_, p0in_reg[2]);
  and _52420_ (_00831_, _42963_, p0_in[2]);
  or _52421_ (_00832_, _00831_, _00830_);
  or _52422_ (_00833_, _00832_, _00814_);
  not _52423_ (_00834_, _00814_);
  or _52424_ (_00835_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _52425_ (_00836_, _00835_, _00833_);
  and _52426_ (_00837_, _00836_, _00795_);
  and _52427_ (_00838_, _42967_, p0in_reg[1]);
  and _52428_ (_00839_, _42963_, p0_in[1]);
  or _52429_ (_00840_, _00839_, _00838_);
  or _52430_ (_00841_, _00840_, _00814_);
  or _52431_ (_00842_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _52432_ (_00843_, _00842_, _00841_);
  and _52433_ (_00844_, _00843_, _00785_);
  or _52434_ (_00845_, _00844_, _00837_);
  or _52435_ (_00846_, _00845_, _00829_);
  or _52436_ (_00847_, _00846_, _00822_);
  and _52437_ (_00848_, _40439_, _40274_);
  not _52438_ (_00849_, _40220_);
  and _52439_ (_00850_, _40492_, _00849_);
  and _52440_ (_00851_, _00850_, _00848_);
  and _52441_ (_00852_, _00851_, _40357_);
  and _52442_ (_00853_, _42967_, p0in_reg[4]);
  and _52443_ (_00854_, _42963_, p0_in[4]);
  or _52444_ (_00855_, _00854_, _00853_);
  or _52445_ (_00856_, _00855_, _00814_);
  or _52446_ (_00857_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _52447_ (_00858_, _00857_, _00856_);
  and _52448_ (_00859_, _00858_, _00777_);
  or _52449_ (_00860_, _00859_, _40313_);
  and _52450_ (_00861_, _42967_, p0in_reg[7]);
  and _52451_ (_00862_, _42963_, p0_in[7]);
  or _52452_ (_00864_, _00862_, _00861_);
  or _52453_ (_00865_, _00864_, _00814_);
  or _52454_ (_00866_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _52455_ (_00867_, _00866_, _00865_);
  and _52456_ (_00868_, _00867_, _00781_);
  and _52457_ (_00869_, _42967_, p0in_reg[6]);
  and _52458_ (_00870_, _42963_, p0_in[6]);
  or _52459_ (_00871_, _00870_, _00869_);
  or _52460_ (_00872_, _00871_, _00814_);
  or _52461_ (_00873_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _52462_ (_00874_, _00873_, _00872_);
  and _52463_ (_00875_, _00874_, _00795_);
  and _52464_ (_00876_, _42967_, p0in_reg[5]);
  and _52465_ (_00877_, _42963_, p0_in[5]);
  or _52466_ (_00878_, _00877_, _00876_);
  or _52467_ (_00879_, _00878_, _00814_);
  or _52468_ (_00880_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _52469_ (_00881_, _00880_, _00879_);
  and _52470_ (_00882_, _00881_, _00785_);
  or _52471_ (_00883_, _00882_, _00875_);
  or _52472_ (_00884_, _00883_, _00868_);
  or _52473_ (_00885_, _00884_, _00860_);
  and _52474_ (_00886_, _00885_, _00852_);
  and _52475_ (_00887_, _00886_, _00847_);
  and _52476_ (_00888_, _42967_, p2in_reg[0]);
  and _52477_ (_00889_, _42963_, p2_in[0]);
  or _52478_ (_00890_, _00889_, _00888_);
  or _52479_ (_00891_, _00890_, _00814_);
  or _52480_ (_00892_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _52481_ (_00893_, _00892_, _00891_);
  and _52482_ (_00895_, _00893_, _00777_);
  or _52483_ (_00896_, _00895_, _00753_);
  and _52484_ (_00897_, _42967_, p2in_reg[3]);
  and _52485_ (_00898_, _42963_, p2_in[3]);
  or _52486_ (_00899_, _00898_, _00897_);
  or _52487_ (_00900_, _00899_, _00814_);
  or _52488_ (_00901_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _52489_ (_00902_, _00901_, _00900_);
  and _52490_ (_00903_, _00902_, _00781_);
  and _52491_ (_00904_, _42967_, p2in_reg[1]);
  and _52492_ (_00905_, _42963_, p2_in[1]);
  or _52493_ (_00906_, _00905_, _00904_);
  or _52494_ (_00907_, _00906_, _00814_);
  or _52495_ (_00908_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _52496_ (_00909_, _00908_, _00907_);
  and _52497_ (_00910_, _00909_, _00785_);
  and _52498_ (_00911_, _42967_, p2in_reg[2]);
  and _52499_ (_00912_, _42963_, p2_in[2]);
  or _52500_ (_00913_, _00912_, _00911_);
  or _52501_ (_00914_, _00913_, _00814_);
  or _52502_ (_00916_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _52503_ (_00917_, _00916_, _00914_);
  and _52504_ (_00918_, _00917_, _00795_);
  or _52505_ (_00919_, _00918_, _00910_);
  or _52506_ (_00920_, _00919_, _00903_);
  or _52507_ (_00921_, _00920_, _00896_);
  and _52508_ (_00922_, _00850_, _40357_);
  and _52509_ (_00923_, _40439_, _40275_);
  and _52510_ (_00924_, _00923_, _00922_);
  and _52511_ (_00925_, _42967_, p2in_reg[4]);
  and _52512_ (_00926_, _42963_, p2_in[4]);
  or _52513_ (_00927_, _00926_, _00925_);
  or _52514_ (_00928_, _00927_, _00814_);
  or _52515_ (_00929_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _52516_ (_00930_, _00929_, _00928_);
  and _52517_ (_00931_, _00930_, _00777_);
  or _52518_ (_00932_, _00931_, _40313_);
  and _52519_ (_00933_, _42967_, p2in_reg[7]);
  and _52520_ (_00934_, _42963_, p2_in[7]);
  or _52521_ (_00935_, _00934_, _00933_);
  or _52522_ (_00936_, _00935_, _00814_);
  or _52523_ (_00937_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _52524_ (_00938_, _00937_, _00936_);
  and _52525_ (_00939_, _00938_, _00781_);
  and _52526_ (_00940_, _42967_, p2in_reg[5]);
  and _52527_ (_00941_, _42963_, p2_in[5]);
  or _52528_ (_00942_, _00941_, _00940_);
  or _52529_ (_00943_, _00942_, _00814_);
  or _52530_ (_00944_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _52531_ (_00945_, _00944_, _00943_);
  and _52532_ (_00946_, _00945_, _00785_);
  and _52533_ (_00947_, _42967_, p2in_reg[6]);
  and _52534_ (_00948_, _42963_, p2_in[6]);
  or _52535_ (_00949_, _00948_, _00947_);
  or _52536_ (_00950_, _00949_, _00814_);
  or _52537_ (_00951_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _52538_ (_00952_, _00951_, _00950_);
  and _52539_ (_00953_, _00952_, _00795_);
  or _52540_ (_00954_, _00953_, _00946_);
  or _52541_ (_00955_, _00954_, _00939_);
  or _52542_ (_00956_, _00955_, _00932_);
  and _52543_ (_00957_, _00956_, _00924_);
  and _52544_ (_00958_, _00957_, _00921_);
  or _52545_ (_00959_, _00958_, _00887_);
  and _52546_ (_00960_, _42967_, p1in_reg[4]);
  and _52547_ (_00961_, _42963_, p1_in[4]);
  or _52548_ (_00962_, _00961_, _00960_);
  or _52549_ (_00963_, _00962_, _00814_);
  or _52550_ (_00964_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _52551_ (_00965_, _00964_, _00963_);
  and _52552_ (_00966_, _00965_, _00777_);
  or _52553_ (_00967_, _00966_, _40313_);
  and _52554_ (_00968_, _42967_, p1in_reg[7]);
  and _52555_ (_00969_, _42963_, p1_in[7]);
  or _52556_ (_00970_, _00969_, _00968_);
  or _52557_ (_00971_, _00970_, _00814_);
  or _52558_ (_00972_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _52559_ (_00973_, _00972_, _00971_);
  and _52560_ (_00974_, _00973_, _00781_);
  and _52561_ (_00975_, _42967_, p1in_reg[6]);
  and _52562_ (_00976_, _42963_, p1_in[6]);
  or _52563_ (_00977_, _00976_, _00975_);
  or _52564_ (_00978_, _00977_, _00814_);
  or _52565_ (_00979_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _52566_ (_00980_, _00979_, _00978_);
  and _52567_ (_00981_, _00980_, _00795_);
  and _52568_ (_00982_, _42967_, p1in_reg[5]);
  and _52569_ (_00983_, _42963_, p1_in[5]);
  or _52570_ (_00984_, _00983_, _00982_);
  or _52571_ (_00985_, _00984_, _00814_);
  or _52572_ (_00986_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _52573_ (_00987_, _00986_, _00985_);
  and _52574_ (_00988_, _00987_, _00785_);
  or _52575_ (_00989_, _00988_, _00981_);
  or _52576_ (_00990_, _00989_, _00974_);
  or _52577_ (_00991_, _00990_, _00967_);
  nor _52578_ (_00992_, _40492_, _40275_);
  and _52579_ (_00993_, _40439_, _00849_);
  and _52580_ (_00994_, _00993_, _00992_);
  and _52581_ (_00995_, _00994_, _40357_);
  and _52582_ (_00996_, _42967_, p1in_reg[0]);
  and _52583_ (_00997_, _42963_, p1_in[0]);
  or _52584_ (_00998_, _00997_, _00996_);
  or _52585_ (_00999_, _00998_, _00814_);
  or _52586_ (_01000_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _52587_ (_01001_, _01000_, _00999_);
  and _52588_ (_01002_, _01001_, _00777_);
  or _52589_ (_01003_, _01002_, _00753_);
  and _52590_ (_01004_, _42967_, p1in_reg[3]);
  and _52591_ (_01005_, _42963_, p1_in[3]);
  or _52592_ (_01006_, _01005_, _01004_);
  or _52593_ (_01007_, _01006_, _00814_);
  or _52594_ (_01008_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _52595_ (_01009_, _01008_, _01007_);
  and _52596_ (_01010_, _01009_, _00781_);
  and _52597_ (_01011_, _42967_, p1in_reg[2]);
  and _52598_ (_01012_, _42963_, p1_in[2]);
  or _52599_ (_01013_, _01012_, _01011_);
  or _52600_ (_01014_, _01013_, _00814_);
  or _52601_ (_01015_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _52602_ (_01016_, _01015_, _01014_);
  and _52603_ (_01017_, _01016_, _00795_);
  and _52604_ (_01018_, _42967_, p1in_reg[1]);
  and _52605_ (_01019_, _42963_, p1_in[1]);
  or _52606_ (_01020_, _01019_, _01018_);
  or _52607_ (_01021_, _01020_, _00814_);
  or _52608_ (_01022_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _52609_ (_01023_, _01022_, _01021_);
  and _52610_ (_01024_, _01023_, _00785_);
  or _52611_ (_01025_, _01024_, _01017_);
  or _52612_ (_01026_, _01025_, _01010_);
  or _52613_ (_01027_, _01026_, _01003_);
  and _52614_ (_01028_, _01027_, _00995_);
  and _52615_ (_01029_, _01028_, _00991_);
  and _52616_ (_01030_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _52617_ (_01031_, _01030_, _00753_);
  and _52618_ (_01032_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _52619_ (_01033_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _52620_ (_01034_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _52621_ (_01035_, _01034_, _01033_);
  or _52622_ (_01036_, _01035_, _01032_);
  or _52623_ (_01037_, _01036_, _01031_);
  and _52624_ (_01038_, _40357_, _40492_);
  and _52625_ (_01039_, _00749_, _40275_);
  and _52626_ (_01040_, _01039_, _01038_);
  and _52627_ (_01041_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _52628_ (_01042_, _01041_, _40313_);
  and _52629_ (_01043_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _52630_ (_01044_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _52631_ (_01045_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _52632_ (_01046_, _01045_, _01044_);
  or _52633_ (_01047_, _01046_, _01043_);
  or _52634_ (_01048_, _01047_, _01042_);
  and _52635_ (_01049_, _01048_, _01040_);
  and _52636_ (_01050_, _01049_, _01037_);
  or _52637_ (_01051_, _01050_, _01029_);
  and _52638_ (_01052_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _52639_ (_01053_, _01052_, _00753_);
  and _52640_ (_01054_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _52641_ (_01055_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _52642_ (_01056_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _52643_ (_01057_, _01056_, _01055_);
  or _52644_ (_01058_, _01057_, _01054_);
  or _52645_ (_01059_, _01058_, _01053_);
  and _52646_ (_01060_, _00851_, _40358_);
  and _52647_ (_01061_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or _52648_ (_01062_, _01061_, _40313_);
  and _52649_ (_01063_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _52650_ (_01064_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _52651_ (_01065_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _52652_ (_01066_, _01065_, _01064_);
  or _52653_ (_01067_, _01066_, _01063_);
  or _52654_ (_01068_, _01067_, _01062_);
  and _52655_ (_01069_, _01068_, _01060_);
  and _52656_ (_01070_, _01069_, _01059_);
  and _52657_ (_01071_, _42967_, p3in_reg[0]);
  and _52658_ (_01072_, _42963_, p3_in[0]);
  or _52659_ (_01073_, _01072_, _01071_);
  or _52660_ (_01074_, _01073_, _00814_);
  or _52661_ (_01075_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _52662_ (_01076_, _01075_, _01074_);
  and _52663_ (_01077_, _01076_, _00777_);
  or _52664_ (_01078_, _01077_, _00753_);
  and _52665_ (_01079_, _42967_, p3in_reg[3]);
  and _52666_ (_01080_, _42963_, p3_in[3]);
  or _52667_ (_01081_, _01080_, _01079_);
  or _52668_ (_01082_, _01081_, _00814_);
  or _52669_ (_01083_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _52670_ (_01084_, _01083_, _01082_);
  and _52671_ (_01085_, _01084_, _00781_);
  and _52672_ (_01086_, _42967_, p3in_reg[1]);
  and _52673_ (_01087_, _42963_, p3_in[1]);
  or _52674_ (_01088_, _01087_, _01086_);
  or _52675_ (_01089_, _01088_, _00814_);
  or _52676_ (_01090_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _52677_ (_01091_, _01090_, _01089_);
  and _52678_ (_01092_, _01091_, _00785_);
  and _52679_ (_01093_, _42967_, p3in_reg[2]);
  and _52680_ (_01094_, _42963_, p3_in[2]);
  or _52681_ (_01095_, _01094_, _01093_);
  or _52682_ (_01096_, _01095_, _00814_);
  or _52683_ (_01097_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _52684_ (_01098_, _01097_, _01096_);
  and _52685_ (_01099_, _01098_, _00795_);
  or _52686_ (_01100_, _01099_, _01092_);
  or _52687_ (_01101_, _01100_, _01085_);
  or _52688_ (_01102_, _01101_, _01078_);
  nor _52689_ (_01103_, _40492_, _40274_);
  and _52690_ (_01104_, _01103_, _00993_);
  and _52691_ (_01105_, _01104_, _40357_);
  and _52692_ (_01106_, _42967_, p3in_reg[4]);
  and _52693_ (_01107_, _42963_, p3_in[4]);
  or _52694_ (_01108_, _01107_, _01106_);
  or _52695_ (_01109_, _01108_, _00814_);
  or _52696_ (_01110_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _52697_ (_01111_, _01110_, _01109_);
  and _52698_ (_01112_, _01111_, _00777_);
  or _52699_ (_01113_, _01112_, _40313_);
  and _52700_ (_01114_, _42967_, p3in_reg[7]);
  and _52701_ (_01115_, _42963_, p3_in[7]);
  or _52702_ (_01116_, _01115_, _01114_);
  or _52703_ (_01117_, _01116_, _00814_);
  or _52704_ (_01118_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _52705_ (_01119_, _01118_, _01117_);
  and _52706_ (_01120_, _01119_, _00781_);
  and _52707_ (_01121_, _42967_, p3in_reg[5]);
  and _52708_ (_01122_, _42963_, p3_in[5]);
  or _52709_ (_01123_, _01122_, _01121_);
  or _52710_ (_01124_, _01123_, _00814_);
  or _52711_ (_01125_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _52712_ (_01126_, _01125_, _01124_);
  and _52713_ (_01127_, _01126_, _00785_);
  and _52714_ (_01128_, _42967_, p3in_reg[6]);
  and _52715_ (_01129_, _42963_, p3_in[6]);
  or _52716_ (_01130_, _01129_, _01128_);
  or _52717_ (_01131_, _01130_, _00814_);
  or _52718_ (_01132_, _00834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _52719_ (_01133_, _01132_, _01131_);
  and _52720_ (_01134_, _01133_, _00795_);
  or _52721_ (_01135_, _01134_, _01127_);
  or _52722_ (_01136_, _01135_, _01120_);
  or _52723_ (_01137_, _01136_, _01113_);
  and _52724_ (_01138_, _01137_, _01105_);
  and _52725_ (_01139_, _01138_, _01102_);
  or _52726_ (_01140_, _01139_, _01070_);
  or _52727_ (_01141_, _01140_, _01051_);
  or _52728_ (_01142_, _01141_, _00959_);
  nor _52729_ (_01143_, _01105_, _00995_);
  nor _52730_ (_01144_, _00924_, _00852_);
  and _52731_ (_01145_, _01144_, _01143_);
  and _52732_ (_01146_, _00994_, _40358_);
  and _52733_ (_01147_, _00850_, _40358_);
  and _52734_ (_01148_, _01147_, _00923_);
  and _52735_ (_01149_, _01104_, _40358_);
  and _52736_ (_01150_, _01039_, _00750_);
  or _52737_ (_01151_, _01040_, _00752_);
  or _52738_ (_01152_, _01151_, _01150_);
  or _52739_ (_01153_, _01152_, _01149_);
  or _52740_ (_01154_, _01153_, _01148_);
  or _52741_ (_01155_, _01154_, _01146_);
  nor _52742_ (_01156_, _01155_, _01060_);
  and _52743_ (_01157_, _01156_, _01145_);
  nand _52744_ (_01158_, _43063_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or _52745_ (_01159_, _01158_, _01157_);
  and _52746_ (_01160_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _52747_ (_01161_, _01160_, _00753_);
  and _52748_ (_01162_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _52749_ (_01163_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _52750_ (_01164_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _52751_ (_01165_, _01164_, _01163_);
  or _52752_ (_01166_, _01165_, _01162_);
  or _52753_ (_01167_, _01166_, _01161_);
  and _52754_ (_01168_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _52755_ (_01169_, _01168_, _40313_);
  and _52756_ (_01170_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _52757_ (_01171_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _52758_ (_01172_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _52759_ (_01173_, _01172_, _01171_);
  or _52760_ (_01174_, _01173_, _01170_);
  or _52761_ (_01175_, _01174_, _01169_);
  and _52762_ (_01176_, _01175_, _01149_);
  and _52763_ (_01177_, _01176_, _01167_);
  and _52764_ (_01178_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _52765_ (_01179_, _01178_, _00753_);
  and _52766_ (_01180_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _52767_ (_01181_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _52768_ (_01182_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _52769_ (_01183_, _01182_, _01181_);
  or _52770_ (_01184_, _01183_, _01180_);
  or _52771_ (_01185_, _01184_, _01179_);
  and _52772_ (_01186_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _52773_ (_01187_, _01186_, _40313_);
  and _52774_ (_01188_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _52775_ (_01189_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _52776_ (_01190_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _52777_ (_01191_, _01190_, _01189_);
  or _52778_ (_01192_, _01191_, _01188_);
  or _52779_ (_01193_, _01192_, _01187_);
  and _52780_ (_01194_, _01193_, _01150_);
  and _52781_ (_01195_, _01194_, _01185_);
  or _52782_ (_01196_, _01195_, _01177_);
  and _52783_ (_01197_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _52784_ (_01198_, _01197_, _00753_);
  and _52785_ (_01199_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _52786_ (_01200_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _52787_ (_01201_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _52788_ (_01202_, _01201_, _01200_);
  or _52789_ (_01203_, _01202_, _01199_);
  or _52790_ (_01204_, _01203_, _01198_);
  and _52791_ (_01205_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _52792_ (_01206_, _01205_, _40313_);
  and _52793_ (_01207_, _00781_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _52794_ (_01208_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _52795_ (_01209_, _00785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _52796_ (_01210_, _01209_, _01208_);
  or _52797_ (_01211_, _01210_, _01207_);
  or _52798_ (_01212_, _01211_, _01206_);
  and _52799_ (_01213_, _01212_, _01148_);
  and _52800_ (_01214_, _01213_, _01204_);
  nor _52801_ (_01215_, _01214_, _01196_);
  nand _52802_ (_01216_, _01215_, _01159_);
  or _52803_ (_01217_, _01216_, _01142_);
  or _52804_ (_01218_, _01217_, _00801_);
  and _52805_ (_01219_, _01040_, _38931_);
  nor _52806_ (_01220_, _01159_, _29134_);
  nor _52807_ (_01221_, _01220_, _01219_);
  and _52808_ (_01222_, _01221_, _01218_);
  or _52809_ (_01223_, _00753_, _38996_);
  or _52810_ (_01224_, _40313_, _39046_);
  and _52811_ (_01225_, _01224_, _00777_);
  and _52812_ (_01226_, _01225_, _01223_);
  and _52813_ (_01227_, _40313_, _39019_);
  and _52814_ (_01228_, _00753_, _39068_);
  or _52815_ (_01229_, _01228_, _01227_);
  and _52816_ (_01230_, _01229_, _00795_);
  or _52817_ (_01231_, _40313_, _39057_);
  or _52818_ (_01232_, _00753_, _39008_);
  and _52819_ (_01233_, _01232_, _00785_);
  and _52820_ (_01234_, _01233_, _01231_);
  and _52821_ (_01235_, _00782_, _38985_);
  not _52822_ (_01236_, _39035_);
  and _52823_ (_01237_, _00790_, _01236_);
  or _52824_ (_01238_, _01237_, _01235_);
  or _52825_ (_01239_, _01238_, _01234_);
  or _52826_ (_01240_, _01239_, _01230_);
  or _52827_ (_01241_, _01240_, _01226_);
  and _52828_ (_01242_, _01241_, _01219_);
  nor _52829_ (_01243_, _01145_, _00814_);
  not _52830_ (_01244_, _01243_);
  and _52831_ (_01245_, _42989_, _38770_);
  and _52832_ (_01246_, _01245_, _01244_);
  not _52833_ (_01247_, _01246_);
  nor _52834_ (_01248_, _01247_, _01157_);
  or _52835_ (_01249_, _01248_, _01242_);
  or _52836_ (_01250_, _01249_, _01222_);
  or _52837_ (_01251_, _40313_, _40432_);
  nand _52838_ (_01252_, _40313_, _38348_);
  and _52839_ (_01253_, _01252_, _00795_);
  and _52840_ (_01254_, _01253_, _01251_);
  or _52841_ (_01255_, _40313_, _40472_);
  nand _52842_ (_01256_, _40313_, _38364_);
  and _52843_ (_01257_, _01256_, _00777_);
  and _52844_ (_01258_, _01257_, _01255_);
  or _52845_ (_01259_, _01258_, _01254_);
  not _52846_ (_01260_, _00782_);
  nor _52847_ (_01261_, _01260_, _38386_);
  and _52848_ (_01262_, _00790_, _40346_);
  or _52849_ (_01263_, _40313_, _40236_);
  nand _52850_ (_01264_, _40313_, _38355_);
  and _52851_ (_01265_, _01264_, _01263_);
  and _52852_ (_01266_, _01265_, _00785_);
  or _52853_ (_01267_, _01266_, _01262_);
  or _52854_ (_01268_, _01267_, _01261_);
  nor _52855_ (_01269_, _01268_, _01259_);
  nand _52856_ (_01270_, _01269_, _01248_);
  and _52857_ (_01271_, _01270_, _41755_);
  and _52858_ (_39594_, _01271_, _01250_);
  and _52859_ (_01272_, _00777_, _40313_);
  and _52860_ (_01273_, _01272_, _01040_);
  and _52861_ (_01274_, _01273_, _38928_);
  and _52862_ (_01275_, _01272_, _00752_);
  and _52863_ (_01276_, _01275_, _38788_);
  and _52864_ (_01277_, _00852_, _00790_);
  and _52865_ (_01278_, _01277_, _38437_);
  or _52866_ (_01279_, _01278_, _01276_);
  nor _52867_ (_01280_, _01279_, _01274_);
  nor _52868_ (_01281_, _01280_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _52869_ (_01282_, _01281_);
  and _52870_ (_01283_, _01272_, _01219_);
  and _52871_ (_01284_, _01260_, _38760_);
  and _52872_ (_01285_, _01284_, _42989_);
  nor _52873_ (_01286_, _01285_, _01283_);
  and _52874_ (_01287_, _01286_, _43066_);
  and _52875_ (_01288_, _01287_, _01282_);
  and _52876_ (_01289_, _40357_, _40313_);
  and _52877_ (_01290_, _01289_, _00851_);
  and _52878_ (_01291_, _01290_, _00795_);
  and _52879_ (_01292_, _01291_, _38437_);
  or _52880_ (_01293_, _01292_, rst);
  nor _52881_ (_39595_, _01293_, _01288_);
  nand _52882_ (_01294_, _01292_, _27841_);
  or _52883_ (_01295_, _01288_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _52884_ (_01296_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _52885_ (_01297_, _01272_, _01149_);
  and _52886_ (_01298_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _52887_ (_01299_, _01298_, _01296_);
  and _52888_ (_01300_, _40358_, _40313_);
  and _52889_ (_01301_, _01300_, _00777_);
  and _52890_ (_01302_, _01301_, _00851_);
  and _52891_ (_01303_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _52892_ (_01304_, _00923_, _00850_);
  and _52893_ (_01305_, _01301_, _01304_);
  and _52894_ (_01306_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _52895_ (_01307_, _01306_, _01303_);
  or _52896_ (_01308_, _01307_, _01299_);
  and _52897_ (_01309_, _01272_, _01150_);
  and _52898_ (_01310_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _52899_ (_01311_, _01289_, _00781_);
  and _52900_ (_01312_, _01311_, _00851_);
  and _52901_ (_01313_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _52902_ (_01314_, _01313_, _01310_);
  and _52903_ (_01315_, _01289_, _00785_);
  and _52904_ (_01316_, _01315_, _00851_);
  and _52905_ (_01317_, _01316_, _38388_);
  and _52906_ (_01318_, _01289_, _00777_);
  and _52907_ (_01319_, _01318_, _01104_);
  and _52908_ (_01320_, _01319_, _01119_);
  or _52909_ (_01321_, _01320_, _01317_);
  or _52910_ (_01322_, _01321_, _01314_);
  or _52911_ (_01323_, _01322_, _01308_);
  and _52912_ (_01324_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _52913_ (_01325_, _01318_, _00994_);
  and _52914_ (_01326_, _01325_, _00973_);
  and _52915_ (_01327_, _01318_, _01304_);
  and _52916_ (_01328_, _01327_, _00938_);
  or _52917_ (_01329_, _01328_, _01326_);
  and _52918_ (_01330_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _52919_ (_01331_, _01318_, _00851_);
  and _52920_ (_01332_, _01331_, _00867_);
  or _52921_ (_01333_, _01332_, _01330_);
  or _52922_ (_01334_, _01333_, _01329_);
  or _52923_ (_01335_, _01334_, _01324_);
  nor _52924_ (_01336_, _01335_, _01323_);
  nand _52925_ (_01337_, _01336_, _01288_);
  and _52926_ (_01338_, _01337_, _01295_);
  or _52927_ (_01339_, _01338_, _01292_);
  and _52928_ (_01340_, _01339_, _41755_);
  and _52929_ (_39596_, _01340_, _01294_);
  and _52930_ (_01341_, _01275_, _00775_);
  and _52931_ (_01342_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _52932_ (_01343_, _01272_, _00995_);
  and _52933_ (_01344_, _01343_, _01001_);
  or _52934_ (_01345_, _01344_, _01342_);
  and _52935_ (_01346_, _01272_, _00852_);
  and _52936_ (_01347_, _01346_, _00820_);
  and _52937_ (_01348_, _01272_, _01060_);
  and _52938_ (_01349_, _01348_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _52939_ (_01350_, _01349_, _01347_);
  or _52940_ (_01351_, _01350_, _01345_);
  and _52941_ (_01352_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _52942_ (_01353_, _01277_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _52943_ (_01354_, _01353_, _01352_);
  and _52944_ (_01355_, _01272_, _00924_);
  and _52945_ (_01356_, _01355_, _00893_);
  and _52946_ (_01357_, _01290_, _00785_);
  and _52947_ (_01358_, _01357_, _40389_);
  or _52948_ (_01359_, _01358_, _01356_);
  or _52949_ (_01360_, _01359_, _01354_);
  and _52950_ (_01361_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _52951_ (_01362_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _52952_ (_01363_, _01362_, _01361_);
  and _52953_ (_01364_, _01272_, _01148_);
  and _52954_ (_01365_, _01364_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _52955_ (_01366_, _01272_, _01105_);
  and _52956_ (_01367_, _01366_, _01076_);
  or _52957_ (_01368_, _01367_, _01365_);
  or _52958_ (_01369_, _01368_, _01363_);
  or _52959_ (_01370_, _01369_, _01360_);
  nor _52960_ (_01371_, _01370_, _01351_);
  nand _52961_ (_01372_, _01371_, _01288_);
  or _52962_ (_01373_, _01372_, _01341_);
  or _52963_ (_01374_, _01288_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _52964_ (_01375_, _01374_, _01373_);
  or _52965_ (_01376_, _01375_, _01292_);
  nand _52966_ (_01377_, _01292_, _29046_);
  and _52967_ (_01378_, _01377_, _41755_);
  and _52968_ (_39659_, _01378_, _01376_);
  not _52969_ (_01379_, _01292_);
  and _52970_ (_01380_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _52971_ (_01381_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or _52972_ (_01382_, _01381_, _01380_);
  and _52973_ (_01383_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _52974_ (_01384_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _52975_ (_01385_, _01384_, _01383_);
  or _52976_ (_01386_, _01385_, _01382_);
  and _52977_ (_01387_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _52978_ (_01388_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _52979_ (_01389_, _01388_, _01387_);
  and _52980_ (_01390_, _01316_, _40496_);
  and _52981_ (_01391_, _01319_, _01091_);
  or _52982_ (_01392_, _01391_, _01390_);
  or _52983_ (_01393_, _01392_, _01389_);
  or _52984_ (_01394_, _01393_, _01386_);
  and _52985_ (_01395_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _52986_ (_01396_, _01325_, _01023_);
  and _52987_ (_01397_, _01327_, _00909_);
  or _52988_ (_01398_, _01397_, _01396_);
  and _52989_ (_01399_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _52990_ (_01400_, _01331_, _00843_);
  or _52991_ (_01401_, _01400_, _01399_);
  or _52992_ (_01402_, _01401_, _01398_);
  or _52993_ (_01403_, _01402_, _01395_);
  or _52994_ (_01404_, _01403_, _01394_);
  and _52995_ (_01405_, _01404_, _01288_);
  nor _52996_ (_01406_, _01288_, _17195_);
  or _52997_ (_01408_, _01406_, _01405_);
  and _52998_ (_01410_, _01408_, _01379_);
  nor _52999_ (_01412_, _01379_, _29714_);
  or _53000_ (_01414_, _01412_, _01410_);
  and _53001_ (_39660_, _01414_, _41755_);
  and _53002_ (_01417_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _53003_ (_01419_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _53004_ (_01420_, _01419_, _01417_);
  and _53005_ (_01421_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _53006_ (_01422_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _53007_ (_01423_, _01422_, _01421_);
  or _53008_ (_01424_, _01423_, _01420_);
  and _53009_ (_01425_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _53010_ (_01427_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _53011_ (_01428_, _01427_, _01425_);
  and _53012_ (_01430_, _01316_, _40297_);
  and _53013_ (_01431_, _01319_, _01098_);
  or _53014_ (_01432_, _01431_, _01430_);
  or _53015_ (_01434_, _01432_, _01428_);
  or _53016_ (_01435_, _01434_, _01424_);
  and _53017_ (_01436_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _53018_ (_01438_, _01325_, _01016_);
  and _53019_ (_01439_, _01327_, _00917_);
  or _53020_ (_01440_, _01439_, _01438_);
  and _53021_ (_01442_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _53022_ (_01443_, _01331_, _00836_);
  or _53023_ (_01444_, _01443_, _01442_);
  or _53024_ (_01446_, _01444_, _01440_);
  or _53025_ (_01447_, _01446_, _01436_);
  or _53026_ (_01448_, _01447_, _01435_);
  and _53027_ (_01450_, _01448_, _01288_);
  nor _53028_ (_01451_, _01288_, _15846_);
  or _53029_ (_01452_, _01451_, _01450_);
  and _53030_ (_01454_, _01452_, _01379_);
  nor _53031_ (_01455_, _01379_, _30404_);
  or _53032_ (_01456_, _01455_, _01454_);
  and _53033_ (_39661_, _01456_, _41755_);
  and _53034_ (_01458_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _53035_ (_01459_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _53036_ (_01460_, _01459_, _01458_);
  and _53037_ (_01461_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _53038_ (_01462_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _53039_ (_01463_, _01462_, _01461_);
  or _53040_ (_01464_, _01463_, _01460_);
  and _53041_ (_01465_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _53042_ (_01466_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _53043_ (_01467_, _01466_, _01465_);
  and _53044_ (_01468_, _01316_, _40352_);
  and _53045_ (_01469_, _01319_, _01084_);
  or _53046_ (_01470_, _01469_, _01468_);
  or _53047_ (_01471_, _01470_, _01467_);
  or _53048_ (_01472_, _01471_, _01464_);
  and _53049_ (_01473_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _53050_ (_01474_, _01325_, _01009_);
  and _53051_ (_01475_, _01327_, _00902_);
  or _53052_ (_01476_, _01475_, _01474_);
  and _53053_ (_01477_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _53054_ (_01479_, _01331_, _00828_);
  or _53055_ (_01480_, _01479_, _01477_);
  or _53056_ (_01482_, _01480_, _01476_);
  or _53057_ (_01483_, _01482_, _01473_);
  or _53058_ (_01484_, _01483_, _01472_);
  and _53059_ (_01486_, _01484_, _01288_);
  nor _53060_ (_01487_, _01288_, _16878_);
  or _53061_ (_01488_, _01487_, _01486_);
  and _53062_ (_01490_, _01488_, _01379_);
  nor _53063_ (_01491_, _01379_, _31213_);
  or _53064_ (_01492_, _01491_, _01490_);
  and _53065_ (_39662_, _01492_, _41755_);
  and _53066_ (_01494_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _53067_ (_01495_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or _53068_ (_01497_, _01495_, _01494_);
  and _53069_ (_01498_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _53070_ (_01499_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _53071_ (_01501_, _01499_, _01498_);
  or _53072_ (_01502_, _01501_, _01497_);
  and _53073_ (_01503_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _53074_ (_01505_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _53075_ (_01506_, _01505_, _01503_);
  and _53076_ (_01507_, _01316_, _40486_);
  and _53077_ (_01509_, _01319_, _01111_);
  or _53078_ (_01510_, _01509_, _01507_);
  or _53079_ (_01511_, _01510_, _01506_);
  or _53080_ (_01512_, _01511_, _01502_);
  and _53081_ (_01513_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _53082_ (_01514_, _01325_, _00965_);
  and _53083_ (_01515_, _01327_, _00930_);
  or _53084_ (_01516_, _01515_, _01514_);
  and _53085_ (_01517_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _53086_ (_01518_, _01331_, _00858_);
  or _53087_ (_01519_, _01518_, _01517_);
  or _53088_ (_01520_, _01519_, _01516_);
  or _53089_ (_01521_, _01520_, _01513_);
  or _53090_ (_01522_, _01521_, _01512_);
  and _53091_ (_01523_, _01522_, _01288_);
  nor _53092_ (_01524_, _01288_, _16044_);
  or _53093_ (_01525_, _01524_, _01523_);
  and _53094_ (_01526_, _01525_, _01379_);
  nor _53095_ (_01527_, _01379_, _31997_);
  or _53096_ (_01528_, _01527_, _01526_);
  and _53097_ (_39663_, _01528_, _41755_);
  and _53098_ (_01530_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _53099_ (_01531_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or _53100_ (_01533_, _01531_, _01530_);
  and _53101_ (_01534_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _53102_ (_01535_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _53103_ (_01537_, _01535_, _01534_);
  or _53104_ (_01538_, _01537_, _01533_);
  and _53105_ (_01539_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _53106_ (_01541_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _53107_ (_01542_, _01541_, _01539_);
  and _53108_ (_01543_, _01316_, _40254_);
  and _53109_ (_01545_, _01319_, _01126_);
  or _53110_ (_01546_, _01545_, _01543_);
  or _53111_ (_01547_, _01546_, _01542_);
  or _53112_ (_01549_, _01547_, _01538_);
  and _53113_ (_01550_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _53114_ (_01551_, _01325_, _00987_);
  and _53115_ (_01553_, _01327_, _00945_);
  or _53116_ (_01554_, _01553_, _01551_);
  and _53117_ (_01555_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _53118_ (_01557_, _01331_, _00881_);
  or _53119_ (_01558_, _01557_, _01555_);
  or _53120_ (_01559_, _01558_, _01554_);
  or _53121_ (_01561_, _01559_, _01550_);
  or _53122_ (_01562_, _01561_, _01549_);
  and _53123_ (_01563_, _01562_, _01288_);
  nor _53124_ (_01564_, _01288_, _17032_);
  or _53125_ (_01565_, _01564_, _01563_);
  and _53126_ (_01566_, _01565_, _01379_);
  nor _53127_ (_01567_, _01379_, _32814_);
  or _53128_ (_01568_, _01567_, _01566_);
  and _53129_ (_39664_, _01568_, _41755_);
  and _53130_ (_01569_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _53131_ (_01570_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or _53132_ (_01571_, _01570_, _01569_);
  and _53133_ (_01572_, _01302_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _53134_ (_01573_, _01305_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or _53135_ (_01574_, _01573_, _01572_);
  or _53136_ (_01575_, _01574_, _01571_);
  and _53137_ (_01576_, _01309_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _53138_ (_01577_, _01312_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _53139_ (_01578_, _01577_, _01576_);
  and _53140_ (_01579_, _01316_, _40404_);
  and _53141_ (_01580_, _01319_, _01133_);
  or _53142_ (_01582_, _01580_, _01579_);
  or _53143_ (_01583_, _01582_, _01578_);
  or _53144_ (_01585_, _01583_, _01575_);
  and _53145_ (_01586_, _01273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _53146_ (_01587_, _01325_, _00980_);
  and _53147_ (_01589_, _01327_, _00952_);
  or _53148_ (_01590_, _01589_, _01587_);
  and _53149_ (_01591_, _01275_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _53150_ (_01593_, _01331_, _00874_);
  or _53151_ (_01594_, _01593_, _01591_);
  or _53152_ (_01595_, _01594_, _01590_);
  or _53153_ (_01597_, _01595_, _01586_);
  or _53154_ (_01598_, _01597_, _01585_);
  and _53155_ (_01599_, _01598_, _01288_);
  nor _53156_ (_01601_, _01288_, _16384_);
  or _53157_ (_01602_, _01601_, _01599_);
  and _53158_ (_01603_, _01602_, _01379_);
  nor _53159_ (_01605_, _01379_, _33533_);
  or _53160_ (_01606_, _01605_, _01603_);
  and _53161_ (_39665_, _01606_, _41755_);
  and _53162_ (_39709_, _40598_, _41755_);
  and _53163_ (_39710_, _40777_, _41755_);
  nor _53164_ (_39712_, _40313_, rst);
  and _53165_ (_39728_, _40795_, _41755_);
  and _53166_ (_39729_, _40808_, _41755_);
  and _53167_ (_39730_, _40821_, _41755_);
  and _53168_ (_39731_, _40829_, _41755_);
  and _53169_ (_39732_, _40840_, _41755_);
  and _53170_ (_39733_, _40851_, _41755_);
  and _53171_ (_39734_, _40862_, _41755_);
  nor _53172_ (_39735_, _40393_, rst);
  nor _53173_ (_39736_, _40558_, rst);
  not _53174_ (_01609_, _41953_);
  nor _53175_ (_01610_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _53176_ (_01611_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53177_ (_01612_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01611_);
  nor _53178_ (_01613_, _01612_, _01610_);
  nor _53179_ (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53180_ (_01615_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01611_);
  nor _53181_ (_01616_, _01615_, _01614_);
  nor _53182_ (_01617_, _01616_, _01613_);
  not _53183_ (_01618_, _01617_);
  nor _53184_ (_01619_, _00104_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53185_ (_01621_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01611_);
  nor _53186_ (_01622_, _01621_, _01619_);
  and _53187_ (_01624_, _01622_, _01618_);
  nor _53188_ (_01625_, _01622_, _01618_);
  nor _53189_ (_01626_, _01625_, _01624_);
  nor _53190_ (_01628_, _00123_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _53191_ (_01629_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01611_);
  nor _53192_ (_01630_, _01629_, _01628_);
  not _53193_ (_01632_, _01630_);
  and _53194_ (_01633_, _01632_, _01624_);
  nor _53195_ (_01634_, _01632_, _01624_);
  nor _53196_ (_01636_, _01634_, _01633_);
  nor _53197_ (_01637_, _01636_, _01626_);
  not _53198_ (_01638_, _01613_);
  nor _53199_ (_01640_, _01616_, _01638_);
  and _53200_ (_01641_, _01640_, _01637_);
  and _53201_ (_01642_, _01641_, _01609_);
  not _53202_ (_01644_, _41994_);
  and _53203_ (_01645_, _01616_, _01638_);
  and _53204_ (_01646_, _01645_, _01637_);
  and _53205_ (_01648_, _01646_, _01644_);
  not _53206_ (_01649_, _41692_);
  and _53207_ (_01650_, _01616_, _01613_);
  not _53208_ (_01652_, _01626_);
  and _53209_ (_01653_, _01636_, _01652_);
  and _53210_ (_01654_, _01653_, _01650_);
  and _53211_ (_01655_, _01654_, _01649_);
  or _53212_ (_01656_, _01655_, _01648_);
  or _53213_ (_01657_, _01656_, _01642_);
  not _53214_ (_01658_, _41830_);
  and _53215_ (_01659_, _01632_, _01626_);
  and _53216_ (_01660_, _01659_, _01645_);
  and _53217_ (_01661_, _01660_, _01658_);
  not _53218_ (_01662_, _42240_);
  and _53219_ (_01663_, _01622_, _01617_);
  and _53220_ (_01664_, _01630_, _01663_);
  and _53221_ (_01665_, _01664_, _01662_);
  not _53222_ (_01666_, _42076_);
  and _53223_ (_01667_, _01630_, _01625_);
  and _53224_ (_01668_, _01667_, _01666_);
  or _53225_ (_01669_, _01668_, _01665_);
  not _53226_ (_01670_, _41912_);
  and _53227_ (_01671_, _01632_, _01663_);
  and _53228_ (_01672_, _01671_, _01670_);
  not _53229_ (_01674_, _41740_);
  and _53230_ (_01675_, _01632_, _01625_);
  and _53231_ (_01677_, _01675_, _01674_);
  or _53232_ (_01678_, _01677_, _01672_);
  or _53233_ (_01679_, _01678_, _01669_);
  or _53234_ (_01681_, _01679_, _01661_);
  not _53235_ (_01682_, _41871_);
  and _53236_ (_01683_, _01659_, _01650_);
  and _53237_ (_01685_, _01683_, _01682_);
  not _53238_ (_01686_, _41789_);
  and _53239_ (_01687_, _01659_, _01640_);
  and _53240_ (_01689_, _01687_, _01686_);
  or _53241_ (_01690_, _01689_, _01685_);
  or _53242_ (_01691_, _01690_, _01681_);
  not _53243_ (_01693_, _42035_);
  and _53244_ (_01694_, _01650_, _01637_);
  and _53245_ (_01695_, _01694_, _01693_);
  not _53246_ (_01697_, _42199_);
  and _53247_ (_01698_, _01650_, _01634_);
  and _53248_ (_01699_, _01698_, _01697_);
  not _53249_ (_01701_, _42158_);
  and _53250_ (_01702_, _01645_, _01634_);
  and _53251_ (_01703_, _01702_, _01701_);
  not _53252_ (_01705_, _42117_);
  and _53253_ (_01706_, _01640_, _01634_);
  and _53254_ (_01707_, _01706_, _01705_);
  or _53255_ (_01708_, _01707_, _01703_);
  or _53256_ (_01709_, _01708_, _01699_);
  or _53257_ (_01710_, _01709_, _01695_);
  not _53258_ (_01711_, _41610_);
  and _53259_ (_01712_, _01653_, _01640_);
  and _53260_ (_01713_, _01712_, _01711_);
  not _53261_ (_01714_, _41651_);
  and _53262_ (_01715_, _01653_, _01645_);
  and _53263_ (_01716_, _01715_, _01714_);
  or _53264_ (_01717_, _01716_, _01713_);
  or _53265_ (_01718_, _01717_, _01710_);
  or _53266_ (_01719_, _01718_, _01691_);
  or _53267_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01719_, _01657_);
  and _53268_ (_01720_, _01715_, _01662_);
  and _53269_ (_01721_, _01712_, _01697_);
  and _53270_ (_01722_, _01694_, _01609_);
  or _53271_ (_01723_, _01722_, _01721_);
  or _53272_ (_01724_, _01723_, _01720_);
  and _53273_ (_01726_, _01660_, _01674_);
  and _53274_ (_01727_, _01667_, _01644_);
  and _53275_ (_01729_, _01671_, _01658_);
  or _53276_ (_01730_, _01729_, _01727_);
  and _53277_ (_01731_, _01664_, _01701_);
  and _53278_ (_01733_, _01675_, _01714_);
  or _53279_ (_01734_, _01733_, _01731_);
  or _53280_ (_01735_, _01734_, _01730_);
  or _53281_ (_01737_, _01735_, _01726_);
  and _53282_ (_01738_, _01687_, _01649_);
  and _53283_ (_01739_, _01683_, _01686_);
  or _53284_ (_01741_, _01739_, _01738_);
  or _53285_ (_01742_, _01741_, _01737_);
  and _53286_ (_01743_, _01646_, _01670_);
  and _53287_ (_01745_, _01702_, _01666_);
  and _53288_ (_01746_, _01698_, _01705_);
  and _53289_ (_01747_, _01706_, _01693_);
  or _53290_ (_01749_, _01747_, _01746_);
  or _53291_ (_01750_, _01749_, _01745_);
  or _53292_ (_01751_, _01750_, _01743_);
  and _53293_ (_01753_, _01654_, _01711_);
  and _53294_ (_01754_, _01641_, _01682_);
  or _53295_ (_01755_, _01754_, _01753_);
  or _53296_ (_01757_, _01755_, _01751_);
  or _53297_ (_01758_, _01757_, _01742_);
  or _53298_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01758_, _01724_);
  and _53299_ (_01759_, _01698_, _01701_);
  and _53300_ (_01760_, _01706_, _01666_);
  and _53301_ (_01761_, _01702_, _01705_);
  or _53302_ (_01762_, _01761_, _01760_);
  or _53303_ (_01763_, _01762_, _01759_);
  and _53304_ (_01764_, _01712_, _01662_);
  and _53305_ (_01765_, _01646_, _01609_);
  or _53306_ (_01766_, _01765_, _01764_);
  or _53307_ (_01767_, _01766_, _01763_);
  and _53308_ (_01768_, _01687_, _01674_);
  and _53309_ (_01769_, _01671_, _01682_);
  and _53310_ (_01770_, _01683_, _01658_);
  or _53311_ (_01771_, _01770_, _01769_);
  or _53312_ (_01772_, _01771_, _01768_);
  and _53313_ (_01773_, _01654_, _01714_);
  and _53314_ (_01774_, _01660_, _01686_);
  or _53315_ (_01775_, _01774_, _01773_);
  or _53316_ (_01776_, _01775_, _01772_);
  or _53317_ (_01778_, _01776_, _01767_);
  and _53318_ (_01779_, _01641_, _01670_);
  and _53319_ (_01781_, _01694_, _01644_);
  and _53320_ (_01782_, _01667_, _01693_);
  or _53321_ (_01783_, _01782_, _01781_);
  or _53322_ (_01785_, _01783_, _01779_);
  and _53323_ (_01786_, _01664_, _01697_);
  and _53324_ (_01787_, _01675_, _01649_);
  and _53325_ (_01789_, _01715_, _01711_);
  or _53326_ (_01790_, _01789_, _01787_);
  or _53327_ (_01791_, _01790_, _01786_);
  or _53328_ (_01793_, _01791_, _01785_);
  or _53329_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01793_, _01778_);
  and _53330_ (_01794_, _01646_, _01682_);
  and _53331_ (_01796_, _01641_, _01658_);
  and _53332_ (_01797_, _01712_, _01701_);
  or _53333_ (_01798_, _01797_, _01796_);
  or _53334_ (_01800_, _01798_, _01794_);
  and _53335_ (_01801_, _01660_, _01649_);
  and _53336_ (_01802_, _01687_, _01714_);
  or _53337_ (_01804_, _01802_, _01801_);
  and _53338_ (_01805_, _01683_, _01674_);
  and _53339_ (_01806_, _01671_, _01686_);
  and _53340_ (_01808_, _01667_, _01609_);
  or _53341_ (_01809_, _01808_, _01806_);
  and _53342_ (_01810_, _01675_, _01711_);
  and _53343_ (_01811_, _01664_, _01705_);
  or _53344_ (_01812_, _01811_, _01810_);
  or _53345_ (_01813_, _01812_, _01809_);
  or _53346_ (_01814_, _01813_, _01805_);
  or _53347_ (_01815_, _01814_, _01804_);
  and _53348_ (_01816_, _01715_, _01697_);
  and _53349_ (_01817_, _01702_, _01693_);
  and _53350_ (_01818_, _01706_, _01644_);
  or _53351_ (_01819_, _01818_, _01817_);
  and _53352_ (_01820_, _01698_, _01666_);
  or _53353_ (_01821_, _01820_, _01819_);
  or _53354_ (_01822_, _01821_, _01816_);
  and _53355_ (_01823_, _01654_, _01662_);
  and _53356_ (_01824_, _01694_, _01670_);
  or _53357_ (_01825_, _01824_, _01823_);
  or _53358_ (_01826_, _01825_, _01822_);
  or _53359_ (_01827_, _01826_, _01815_);
  or _53360_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01827_, _01800_);
  not _53361_ (_01829_, _42081_);
  and _53362_ (_01830_, _01702_, _01829_);
  not _53363_ (_01832_, _42122_);
  and _53364_ (_01833_, _01698_, _01832_);
  or _53365_ (_01834_, _01833_, _01830_);
  not _53366_ (_01836_, _42204_);
  and _53367_ (_01837_, _01712_, _01836_);
  or _53368_ (_01838_, _01837_, _01834_);
  not _53369_ (_01840_, _41958_);
  and _53370_ (_01841_, _01694_, _01840_);
  not _53371_ (_01842_, _42245_);
  and _53372_ (_01844_, _01715_, _01842_);
  or _53373_ (_01845_, _01844_, _01841_);
  or _53374_ (_01846_, _01845_, _01838_);
  not _53375_ (_01848_, _41835_);
  and _53376_ (_01849_, _01671_, _01848_);
  not _53377_ (_01850_, _41749_);
  and _53378_ (_01852_, _01660_, _01850_);
  not _53379_ (_01853_, _41794_);
  and _53380_ (_01854_, _01683_, _01853_);
  or _53381_ (_01856_, _01854_, _01852_);
  or _53382_ (_01857_, _01856_, _01849_);
  not _53383_ (_01858_, _41656_);
  and _53384_ (_01860_, _01675_, _01858_);
  not _53385_ (_01861_, _41876_);
  and _53386_ (_01862_, _01641_, _01861_);
  or _53387_ (_01863_, _01862_, _01860_);
  or _53388_ (_01864_, _01863_, _01857_);
  or _53389_ (_01865_, _01864_, _01846_);
  not _53390_ (_01866_, _42163_);
  and _53391_ (_01867_, _01664_, _01866_);
  not _53392_ (_01868_, _41615_);
  and _53393_ (_01869_, _01654_, _01868_);
  not _53394_ (_01870_, _41697_);
  and _53395_ (_01871_, _01687_, _01870_);
  or _53396_ (_01872_, _01871_, _01869_);
  not _53397_ (_01873_, _41917_);
  and _53398_ (_01874_, _01646_, _01873_);
  not _53399_ (_01875_, _41999_);
  and _53400_ (_01876_, _01667_, _01875_);
  not _53401_ (_01877_, _42040_);
  and _53402_ (_01878_, _01706_, _01877_);
  or _53403_ (_01879_, _01878_, _01876_);
  or _53404_ (_01880_, _01879_, _01874_);
  or _53405_ (_01882_, _01880_, _01872_);
  or _53406_ (_01883_, _01882_, _01867_);
  or _53407_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01883_, _01865_);
  not _53408_ (_01885_, _42209_);
  and _53409_ (_01886_, _01712_, _01885_);
  not _53410_ (_01888_, _42250_);
  and _53411_ (_01889_, _01715_, _01888_);
  not _53412_ (_01890_, _41620_);
  and _53413_ (_01892_, _01654_, _01890_);
  or _53414_ (_01893_, _01892_, _01889_);
  or _53415_ (_01894_, _01893_, _01886_);
  not _53416_ (_01896_, _41758_);
  and _53417_ (_01897_, _01660_, _01896_);
  not _53418_ (_01898_, _41799_);
  and _53419_ (_01900_, _01683_, _01898_);
  or _53420_ (_01901_, _01900_, _01897_);
  not _53421_ (_01902_, _41706_);
  and _53422_ (_01904_, _01687_, _01902_);
  not _53423_ (_01905_, _41840_);
  and _53424_ (_01906_, _01671_, _01905_);
  not _53425_ (_01908_, _41661_);
  and _53426_ (_01909_, _01675_, _01908_);
  or _53427_ (_01910_, _01909_, _01906_);
  not _53428_ (_01912_, _42004_);
  and _53429_ (_01913_, _01667_, _01912_);
  not _53430_ (_01914_, _42168_);
  and _53431_ (_01915_, _01664_, _01914_);
  or _53432_ (_01916_, _01915_, _01913_);
  or _53433_ (_01917_, _01916_, _01910_);
  or _53434_ (_01918_, _01917_, _01904_);
  or _53435_ (_01919_, _01918_, _01901_);
  not _53436_ (_01920_, _41922_);
  and _53437_ (_01921_, _01646_, _01920_);
  not _53438_ (_01922_, _41963_);
  and _53439_ (_01923_, _01694_, _01922_);
  or _53440_ (_01924_, _01923_, _01921_);
  not _53441_ (_01925_, _41881_);
  and _53442_ (_01926_, _01641_, _01925_);
  not _53443_ (_01927_, _42127_);
  and _53444_ (_01928_, _01698_, _01927_);
  not _53445_ (_01929_, _42045_);
  and _53446_ (_01930_, _01706_, _01929_);
  not _53447_ (_01931_, _42086_);
  and _53448_ (_01932_, _01702_, _01931_);
  or _53449_ (_01934_, _01932_, _01930_);
  or _53450_ (_01935_, _01934_, _01928_);
  or _53451_ (_01937_, _01935_, _01926_);
  or _53452_ (_01938_, _01937_, _01924_);
  or _53453_ (_01939_, _01938_, _01919_);
  or _53454_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01939_, _01894_);
  not _53455_ (_01941_, _42214_);
  and _53456_ (_01942_, _01712_, _01941_);
  not _53457_ (_01944_, _42132_);
  and _53458_ (_01945_, _01698_, _01944_);
  not _53459_ (_01946_, _42091_);
  and _53460_ (_01948_, _01702_, _01946_);
  or _53461_ (_01949_, _01948_, _01945_);
  or _53462_ (_01950_, _01949_, _01942_);
  not _53463_ (_01952_, _42255_);
  and _53464_ (_01953_, _01715_, _01952_);
  not _53465_ (_01954_, _41968_);
  and _53466_ (_01956_, _01694_, _01954_);
  or _53467_ (_01957_, _01956_, _01953_);
  or _53468_ (_01958_, _01957_, _01950_);
  not _53469_ (_01960_, _41804_);
  and _53470_ (_01961_, _01683_, _01960_);
  not _53471_ (_01962_, _41763_);
  and _53472_ (_01964_, _01660_, _01962_);
  or _53473_ (_01965_, _01964_, _01961_);
  not _53474_ (_01966_, _41845_);
  and _53475_ (_01967_, _01671_, _01966_);
  or _53476_ (_01968_, _01967_, _01965_);
  not _53477_ (_01969_, _41666_);
  and _53478_ (_01970_, _01675_, _01969_);
  not _53479_ (_01971_, _41886_);
  and _53480_ (_01972_, _01641_, _01971_);
  or _53481_ (_01973_, _01972_, _01970_);
  or _53482_ (_01974_, _01973_, _01968_);
  or _53483_ (_01975_, _01974_, _01958_);
  not _53484_ (_01976_, _42173_);
  and _53485_ (_01977_, _01664_, _01976_);
  not _53486_ (_01978_, _41714_);
  and _53487_ (_01979_, _01687_, _01978_);
  not _53488_ (_01980_, _41625_);
  and _53489_ (_01981_, _01654_, _01980_);
  or _53490_ (_01982_, _01981_, _01979_);
  not _53491_ (_01983_, _41927_);
  and _53492_ (_01984_, _01646_, _01983_);
  not _53493_ (_01986_, _42009_);
  and _53494_ (_01987_, _01667_, _01986_);
  not _53495_ (_01989_, _42050_);
  and _53496_ (_01990_, _01706_, _01989_);
  or _53497_ (_01991_, _01990_, _01987_);
  or _53498_ (_01993_, _01991_, _01984_);
  or _53499_ (_01994_, _01993_, _01982_);
  or _53500_ (_01995_, _01994_, _01977_);
  or _53501_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01995_, _01975_);
  not _53502_ (_01997_, _41932_);
  and _53503_ (_01998_, _01646_, _01997_);
  not _53504_ (_02000_, _42260_);
  and _53505_ (_02001_, _01715_, _02000_);
  not _53506_ (_02002_, _41630_);
  and _53507_ (_02004_, _01654_, _02002_);
  or _53508_ (_02005_, _02004_, _02001_);
  or _53509_ (_02006_, _02005_, _01998_);
  not _53510_ (_02008_, _41809_);
  and _53511_ (_02009_, _01683_, _02008_);
  not _53512_ (_02010_, _41850_);
  and _53513_ (_02012_, _01671_, _02010_);
  not _53514_ (_02013_, _41671_);
  and _53515_ (_02014_, _01675_, _02013_);
  or _53516_ (_02016_, _02014_, _02012_);
  not _53517_ (_02017_, _42014_);
  and _53518_ (_02018_, _01667_, _02017_);
  not _53519_ (_02019_, _42178_);
  and _53520_ (_02020_, _01664_, _02019_);
  or _53521_ (_02021_, _02020_, _02018_);
  or _53522_ (_02022_, _02021_, _02016_);
  or _53523_ (_02023_, _02022_, _02009_);
  not _53524_ (_02024_, _41768_);
  and _53525_ (_02025_, _01660_, _02024_);
  not _53526_ (_02026_, _41719_);
  and _53527_ (_02027_, _01687_, _02026_);
  or _53528_ (_02028_, _02027_, _02025_);
  or _53529_ (_02029_, _02028_, _02023_);
  not _53530_ (_02030_, _41973_);
  and _53531_ (_02031_, _01694_, _02030_);
  not _53532_ (_02032_, _42096_);
  and _53533_ (_02033_, _01702_, _02032_);
  not _53534_ (_02034_, _42055_);
  and _53535_ (_02035_, _01706_, _02034_);
  not _53536_ (_02036_, _42137_);
  and _53537_ (_02038_, _01698_, _02036_);
  or _53538_ (_02039_, _02038_, _02035_);
  or _53539_ (_02041_, _02039_, _02033_);
  or _53540_ (_02042_, _02041_, _02031_);
  not _53541_ (_02043_, _42219_);
  and _53542_ (_02045_, _01712_, _02043_);
  not _53543_ (_02046_, _41891_);
  and _53544_ (_02047_, _01641_, _02046_);
  or _53545_ (_02049_, _02047_, _02045_);
  or _53546_ (_02050_, _02049_, _02042_);
  or _53547_ (_02051_, _02050_, _02029_);
  or _53548_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _02051_, _02006_);
  not _53549_ (_02053_, _42101_);
  and _53550_ (_02054_, _01702_, _02053_);
  not _53551_ (_02056_, _42142_);
  and _53552_ (_02057_, _01698_, _02056_);
  or _53553_ (_02058_, _02057_, _02054_);
  not _53554_ (_02060_, _42224_);
  and _53555_ (_02061_, _01712_, _02060_);
  or _53556_ (_02062_, _02061_, _02058_);
  not _53557_ (_02064_, _41978_);
  and _53558_ (_02065_, _01694_, _02064_);
  not _53559_ (_02066_, _42265_);
  and _53560_ (_02068_, _01715_, _02066_);
  or _53561_ (_02069_, _02068_, _02065_);
  or _53562_ (_02070_, _02069_, _02062_);
  not _53563_ (_02071_, _41855_);
  and _53564_ (_02072_, _01671_, _02071_);
  not _53565_ (_02073_, _41773_);
  and _53566_ (_02074_, _01660_, _02073_);
  not _53567_ (_02075_, _41814_);
  and _53568_ (_02076_, _01683_, _02075_);
  or _53569_ (_02077_, _02076_, _02074_);
  or _53570_ (_02078_, _02077_, _02072_);
  not _53571_ (_02079_, _41676_);
  and _53572_ (_02080_, _01675_, _02079_);
  not _53573_ (_02081_, _41896_);
  and _53574_ (_02082_, _01641_, _02081_);
  or _53575_ (_02083_, _02082_, _02080_);
  or _53576_ (_02084_, _02083_, _02078_);
  or _53577_ (_02085_, _02084_, _02070_);
  not _53578_ (_02086_, _42183_);
  and _53579_ (_02087_, _01664_, _02086_);
  not _53580_ (_02088_, _41635_);
  and _53581_ (_02090_, _01654_, _02088_);
  not _53582_ (_02091_, _41724_);
  and _53583_ (_02093_, _01687_, _02091_);
  or _53584_ (_02094_, _02093_, _02090_);
  not _53585_ (_02095_, _41937_);
  and _53586_ (_02097_, _01646_, _02095_);
  not _53587_ (_02098_, _42019_);
  and _53588_ (_02099_, _01667_, _02098_);
  not _53589_ (_02101_, _42060_);
  and _53590_ (_02102_, _01706_, _02101_);
  or _53591_ (_02103_, _02102_, _02099_);
  or _53592_ (_02105_, _02103_, _02097_);
  or _53593_ (_02106_, _02105_, _02094_);
  or _53594_ (_02107_, _02106_, _02087_);
  or _53595_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _02107_, _02085_);
  not _53596_ (_02109_, _42229_);
  and _53597_ (_02110_, _01712_, _02109_);
  not _53598_ (_02112_, _42147_);
  and _53599_ (_02113_, _01698_, _02112_);
  not _53600_ (_02114_, _42106_);
  and _53601_ (_02116_, _01702_, _02114_);
  or _53602_ (_02117_, _02116_, _02113_);
  or _53603_ (_02118_, _02117_, _02110_);
  not _53604_ (_02120_, _42270_);
  and _53605_ (_02121_, _01715_, _02120_);
  not _53606_ (_02122_, _41983_);
  and _53607_ (_02123_, _01694_, _02122_);
  or _53608_ (_02124_, _02123_, _02121_);
  or _53609_ (_02125_, _02124_, _02118_);
  not _53610_ (_02126_, _41819_);
  and _53611_ (_02127_, _01683_, _02126_);
  not _53612_ (_02128_, _41778_);
  and _53613_ (_02129_, _01660_, _02128_);
  or _53614_ (_02130_, _02129_, _02127_);
  not _53615_ (_02131_, _41860_);
  and _53616_ (_02132_, _01671_, _02131_);
  or _53617_ (_02133_, _02132_, _02130_);
  not _53618_ (_02134_, _41681_);
  and _53619_ (_02135_, _01675_, _02134_);
  not _53620_ (_02136_, _41901_);
  and _53621_ (_02137_, _01641_, _02136_);
  or _53622_ (_02138_, _02137_, _02135_);
  or _53623_ (_02139_, _02138_, _02133_);
  or _53624_ (_02140_, _02139_, _02125_);
  not _53625_ (_02142_, _42188_);
  and _53626_ (_02143_, _01664_, _02142_);
  not _53627_ (_02145_, _41729_);
  and _53628_ (_02146_, _01687_, _02145_);
  not _53629_ (_02147_, _41640_);
  and _53630_ (_02149_, _01654_, _02147_);
  or _53631_ (_02150_, _02149_, _02146_);
  not _53632_ (_02151_, _41942_);
  and _53633_ (_02153_, _01646_, _02151_);
  not _53634_ (_02154_, _42024_);
  and _53635_ (_02155_, _01667_, _02154_);
  not _53636_ (_02157_, _42065_);
  and _53637_ (_02158_, _01706_, _02157_);
  or _53638_ (_02159_, _02158_, _02155_);
  or _53639_ (_02161_, _02159_, _02153_);
  or _53640_ (_02162_, _02161_, _02150_);
  or _53641_ (_02163_, _02162_, _02143_);
  or _53642_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _02163_, _02140_);
  not _53643_ (_02165_, _42111_);
  and _53644_ (_02166_, _01702_, _02165_);
  not _53645_ (_02168_, _42152_);
  and _53646_ (_02169_, _01698_, _02168_);
  or _53647_ (_02170_, _02169_, _02166_);
  not _53648_ (_02172_, _42234_);
  and _53649_ (_02173_, _01712_, _02172_);
  or _53650_ (_02174_, _02173_, _02170_);
  not _53651_ (_02175_, _41947_);
  and _53652_ (_02176_, _01646_, _02175_);
  not _53653_ (_02177_, _42275_);
  and _53654_ (_02178_, _01715_, _02177_);
  or _53655_ (_02179_, _02178_, _02176_);
  or _53656_ (_02180_, _02179_, _02174_);
  not _53657_ (_02181_, _41865_);
  and _53658_ (_02182_, _01671_, _02181_);
  not _53659_ (_02183_, _41783_);
  and _53660_ (_02184_, _01660_, _02183_);
  not _53661_ (_02185_, _41824_);
  and _53662_ (_02186_, _01683_, _02185_);
  or _53663_ (_02187_, _02186_, _02184_);
  or _53664_ (_02188_, _02187_, _02182_);
  not _53665_ (_02189_, _41686_);
  and _53666_ (_02190_, _01675_, _02189_);
  not _53667_ (_02191_, _41906_);
  and _53668_ (_02192_, _01641_, _02191_);
  or _53669_ (_02194_, _02192_, _02190_);
  or _53670_ (_02195_, _02194_, _02188_);
  or _53671_ (_02197_, _02195_, _02180_);
  not _53672_ (_02198_, _42193_);
  and _53673_ (_02199_, _01664_, _02198_);
  not _53674_ (_02201_, _41645_);
  and _53675_ (_02202_, _01654_, _02201_);
  not _53676_ (_02203_, _41734_);
  and _53677_ (_02205_, _01687_, _02203_);
  or _53678_ (_02206_, _02205_, _02202_);
  not _53679_ (_02207_, _41988_);
  and _53680_ (_02209_, _01694_, _02207_);
  not _53681_ (_02210_, _42029_);
  and _53682_ (_02211_, _01667_, _02210_);
  not _53683_ (_02213_, _42070_);
  and _53684_ (_02214_, _01706_, _02213_);
  or _53685_ (_02215_, _02214_, _02211_);
  or _53686_ (_02217_, _02215_, _02209_);
  or _53687_ (_02218_, _02217_, _02206_);
  or _53688_ (_02219_, _02218_, _02199_);
  or _53689_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _02219_, _02197_);
  and _53690_ (_02221_, _01646_, _01875_);
  and _53691_ (_02222_, _01694_, _01877_);
  and _53692_ (_02224_, _01641_, _01840_);
  or _53693_ (_02225_, _02224_, _02222_);
  or _53694_ (_02226_, _02225_, _02221_);
  and _53695_ (_02227_, _01660_, _01848_);
  and _53696_ (_02228_, _01683_, _01861_);
  or _53697_ (_02229_, _02228_, _02227_);
  and _53698_ (_02230_, _01687_, _01853_);
  and _53699_ (_02231_, _01671_, _01873_);
  and _53700_ (_02232_, _01675_, _01850_);
  or _53701_ (_02233_, _02232_, _02231_);
  and _53702_ (_02234_, _01664_, _01842_);
  and _53703_ (_02235_, _01667_, _01829_);
  or _53704_ (_02236_, _02235_, _02234_);
  or _53705_ (_02237_, _02236_, _02233_);
  or _53706_ (_02238_, _02237_, _02230_);
  or _53707_ (_02239_, _02238_, _02229_);
  and _53708_ (_02240_, _01706_, _01832_);
  and _53709_ (_02241_, _01702_, _01866_);
  and _53710_ (_02242_, _01698_, _01836_);
  or _53711_ (_02243_, _02242_, _02241_);
  or _53712_ (_02244_, _02243_, _02240_);
  and _53713_ (_02245_, _01654_, _01870_);
  or _53714_ (_02246_, _02245_, _02244_);
  and _53715_ (_02247_, _01712_, _01868_);
  and _53716_ (_02248_, _01715_, _01858_);
  or _53717_ (_02249_, _02248_, _02247_);
  or _53718_ (_02250_, _02249_, _02246_);
  or _53719_ (_02251_, _02250_, _02239_);
  or _53720_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _02251_, _02226_);
  and _53721_ (_02252_, _01694_, _01929_);
  and _53722_ (_02253_, _01646_, _01912_);
  or _53723_ (_02254_, _02253_, _02252_);
  and _53724_ (_02255_, _01641_, _01922_);
  and _53725_ (_02256_, _01671_, _01920_);
  or _53726_ (_02257_, _02256_, _02255_);
  or _53727_ (_02258_, _02257_, _02254_);
  and _53728_ (_02259_, _01683_, _01925_);
  and _53729_ (_02260_, _01660_, _01905_);
  or _53730_ (_02261_, _02260_, _02259_);
  and _53731_ (_02262_, _01687_, _01898_);
  or _53732_ (_02263_, _02262_, _02261_);
  and _53733_ (_02264_, _01675_, _01896_);
  and _53734_ (_02265_, _01715_, _01908_);
  or _53735_ (_02266_, _02265_, _02264_);
  or _53736_ (_02267_, _02266_, _02263_);
  or _53737_ (_02268_, _02267_, _02258_);
  and _53738_ (_02269_, _01698_, _01885_);
  and _53739_ (_02270_, _01702_, _01914_);
  or _53740_ (_02271_, _02270_, _02269_);
  and _53741_ (_02272_, _01667_, _01931_);
  and _53742_ (_02273_, _01706_, _01927_);
  or _53743_ (_02274_, _02273_, _02272_);
  or _53744_ (_02275_, _02274_, _02271_);
  and _53745_ (_02276_, _01664_, _01888_);
  and _53746_ (_02277_, _01654_, _01902_);
  and _53747_ (_02278_, _01712_, _01890_);
  or _53748_ (_02279_, _02278_, _02277_);
  or _53749_ (_02280_, _02279_, _02276_);
  or _53750_ (_02281_, _02280_, _02275_);
  or _53751_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _02281_, _02268_);
  and _53752_ (_02282_, _01641_, _01954_);
  and _53753_ (_02283_, _01694_, _01989_);
  and _53754_ (_02284_, _01646_, _01986_);
  or _53755_ (_02285_, _02284_, _02283_);
  or _53756_ (_02286_, _02285_, _02282_);
  and _53757_ (_02287_, _01683_, _01971_);
  and _53758_ (_02288_, _01660_, _01966_);
  or _53759_ (_02289_, _02288_, _02287_);
  and _53760_ (_02290_, _01687_, _01960_);
  and _53761_ (_02291_, _01671_, _01983_);
  and _53762_ (_02292_, _01675_, _01962_);
  or _53763_ (_02293_, _02292_, _02291_);
  and _53764_ (_02294_, _01664_, _01952_);
  and _53765_ (_02295_, _01667_, _01946_);
  or _53766_ (_02296_, _02295_, _02294_);
  or _53767_ (_02297_, _02296_, _02293_);
  or _53768_ (_02298_, _02297_, _02290_);
  or _53769_ (_02299_, _02298_, _02289_);
  and _53770_ (_02300_, _01654_, _01978_);
  and _53771_ (_02301_, _01698_, _01941_);
  and _53772_ (_02302_, _01702_, _01976_);
  or _53773_ (_02303_, _02302_, _02301_);
  and _53774_ (_02304_, _01706_, _01944_);
  or _53775_ (_02305_, _02304_, _02303_);
  or _53776_ (_02306_, _02305_, _02300_);
  and _53777_ (_02307_, _01712_, _01980_);
  and _53778_ (_02308_, _01715_, _01969_);
  or _53779_ (_02309_, _02308_, _02307_);
  or _53780_ (_02310_, _02309_, _02306_);
  or _53781_ (_02311_, _02310_, _02299_);
  or _53782_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _02311_, _02286_);
  and _53783_ (_02312_, _01641_, _02030_);
  and _53784_ (_02313_, _01694_, _02034_);
  and _53785_ (_02314_, _01646_, _02017_);
  or _53786_ (_02315_, _02314_, _02313_);
  or _53787_ (_02316_, _02315_, _02312_);
  and _53788_ (_02317_, _01683_, _02046_);
  and _53789_ (_02318_, _01671_, _01997_);
  and _53790_ (_02319_, _01675_, _02024_);
  or _53791_ (_02320_, _02319_, _02318_);
  and _53792_ (_02321_, _01664_, _02000_);
  and _53793_ (_02322_, _01667_, _02032_);
  or _53794_ (_02323_, _02322_, _02321_);
  or _53795_ (_02324_, _02323_, _02320_);
  or _53796_ (_02325_, _02324_, _02317_);
  and _53797_ (_02326_, _01660_, _02010_);
  and _53798_ (_02327_, _01687_, _02008_);
  or _53799_ (_02328_, _02327_, _02326_);
  or _53800_ (_02329_, _02328_, _02325_);
  and _53801_ (_02330_, _01654_, _02026_);
  and _53802_ (_02331_, _01698_, _02043_);
  and _53803_ (_02332_, _01702_, _02019_);
  or _53804_ (_02333_, _02332_, _02331_);
  and _53805_ (_02334_, _01706_, _02036_);
  or _53806_ (_02335_, _02334_, _02333_);
  or _53807_ (_02336_, _02335_, _02330_);
  and _53808_ (_02337_, _01712_, _02002_);
  and _53809_ (_02338_, _01715_, _02013_);
  or _53810_ (_02339_, _02338_, _02337_);
  or _53811_ (_02340_, _02339_, _02336_);
  or _53812_ (_02341_, _02340_, _02329_);
  or _53813_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _02341_, _02316_);
  and _53814_ (_02342_, _01646_, _02098_);
  and _53815_ (_02343_, _01694_, _02101_);
  and _53816_ (_02344_, _01641_, _02064_);
  or _53817_ (_02345_, _02344_, _02343_);
  or _53818_ (_02346_, _02345_, _02342_);
  and _53819_ (_02347_, _01683_, _02081_);
  and _53820_ (_02348_, _01660_, _02071_);
  or _53821_ (_02349_, _02348_, _02347_);
  and _53822_ (_02350_, _01687_, _02075_);
  and _53823_ (_02351_, _01671_, _02095_);
  and _53824_ (_02352_, _01675_, _02073_);
  or _53825_ (_02353_, _02352_, _02351_);
  and _53826_ (_02354_, _01664_, _02066_);
  and _53827_ (_02355_, _01667_, _02053_);
  or _53828_ (_02356_, _02355_, _02354_);
  or _53829_ (_02357_, _02356_, _02353_);
  or _53830_ (_02358_, _02357_, _02350_);
  or _53831_ (_02359_, _02358_, _02349_);
  and _53832_ (_02360_, _01654_, _02091_);
  and _53833_ (_02361_, _01702_, _02086_);
  and _53834_ (_02362_, _01698_, _02060_);
  and _53835_ (_02363_, _01706_, _02056_);
  or _53836_ (_02364_, _02363_, _02362_);
  or _53837_ (_02365_, _02364_, _02361_);
  or _53838_ (_02366_, _02365_, _02360_);
  and _53839_ (_02367_, _01712_, _02088_);
  and _53840_ (_02368_, _01715_, _02079_);
  or _53841_ (_02369_, _02368_, _02367_);
  or _53842_ (_02370_, _02369_, _02366_);
  or _53843_ (_02371_, _02370_, _02359_);
  or _53844_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _02371_, _02346_);
  and _53845_ (_02372_, _01641_, _02122_);
  and _53846_ (_02373_, _01654_, _02145_);
  and _53847_ (_02374_, _01646_, _02154_);
  or _53848_ (_02375_, _02374_, _02373_);
  or _53849_ (_02376_, _02375_, _02372_);
  and _53850_ (_02377_, _01683_, _02136_);
  and _53851_ (_02378_, _01675_, _02128_);
  and _53852_ (_02379_, _01671_, _02151_);
  or _53853_ (_02380_, _02379_, _02378_);
  and _53854_ (_02381_, _01664_, _02120_);
  and _53855_ (_02382_, _01667_, _02114_);
  or _53856_ (_02383_, _02382_, _02381_);
  or _53857_ (_02384_, _02383_, _02380_);
  or _53858_ (_02385_, _02384_, _02377_);
  and _53859_ (_02386_, _01660_, _02131_);
  and _53860_ (_02387_, _01687_, _02126_);
  or _53861_ (_02388_, _02387_, _02386_);
  or _53862_ (_02389_, _02388_, _02385_);
  and _53863_ (_02390_, _01694_, _02157_);
  and _53864_ (_02391_, _01698_, _02109_);
  and _53865_ (_02392_, _01702_, _02142_);
  and _53866_ (_02393_, _01706_, _02112_);
  or _53867_ (_02394_, _02393_, _02392_);
  or _53868_ (_02395_, _02394_, _02391_);
  or _53869_ (_02396_, _02395_, _02390_);
  and _53870_ (_02397_, _01712_, _02147_);
  and _53871_ (_02398_, _01715_, _02134_);
  or _53872_ (_02399_, _02398_, _02397_);
  or _53873_ (_02400_, _02399_, _02396_);
  or _53874_ (_02401_, _02400_, _02389_);
  or _53875_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _02401_, _02376_);
  and _53876_ (_02402_, _01641_, _02207_);
  and _53877_ (_02403_, _01694_, _02213_);
  and _53878_ (_02404_, _01646_, _02210_);
  or _53879_ (_02405_, _02404_, _02403_);
  or _53880_ (_02406_, _02405_, _02402_);
  and _53881_ (_02407_, _01683_, _02191_);
  and _53882_ (_02408_, _01660_, _02181_);
  or _53883_ (_02409_, _02408_, _02407_);
  and _53884_ (_02410_, _01687_, _02185_);
  and _53885_ (_02411_, _01671_, _02175_);
  and _53886_ (_02412_, _01675_, _02183_);
  or _53887_ (_02413_, _02412_, _02411_);
  and _53888_ (_02414_, _01664_, _02177_);
  and _53889_ (_02415_, _01667_, _02165_);
  or _53890_ (_02416_, _02415_, _02414_);
  or _53891_ (_02417_, _02416_, _02413_);
  or _53892_ (_02418_, _02417_, _02410_);
  or _53893_ (_02419_, _02418_, _02409_);
  and _53894_ (_02420_, _01654_, _02203_);
  and _53895_ (_02421_, _01698_, _02172_);
  and _53896_ (_02422_, _01702_, _02198_);
  or _53897_ (_02423_, _02422_, _02421_);
  and _53898_ (_02424_, _01706_, _02168_);
  or _53899_ (_02425_, _02424_, _02423_);
  or _53900_ (_02426_, _02425_, _02420_);
  and _53901_ (_02427_, _01712_, _02201_);
  and _53902_ (_02428_, _01715_, _02189_);
  or _53903_ (_02429_, _02428_, _02427_);
  or _53904_ (_02430_, _02429_, _02426_);
  or _53905_ (_02431_, _02430_, _02419_);
  or _53906_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _02431_, _02406_);
  and _53907_ (_02432_, _01715_, _01836_);
  and _53908_ (_02433_, _01694_, _01873_);
  and _53909_ (_02434_, _01641_, _01848_);
  or _53910_ (_02435_, _02434_, _02433_);
  or _53911_ (_02436_, _02435_, _02432_);
  and _53912_ (_02437_, _01660_, _01870_);
  and _53913_ (_02438_, _01664_, _01832_);
  and _53914_ (_02439_, _01671_, _01853_);
  or _53915_ (_02440_, _02439_, _02438_);
  and _53916_ (_02441_, _01667_, _01840_);
  and _53917_ (_02442_, _01675_, _01868_);
  or _53918_ (_02443_, _02442_, _02441_);
  or _53919_ (_02444_, _02443_, _02440_);
  or _53920_ (_02445_, _02444_, _02437_);
  and _53921_ (_02446_, _01687_, _01858_);
  and _53922_ (_02447_, _01683_, _01850_);
  or _53923_ (_02448_, _02447_, _02446_);
  or _53924_ (_02449_, _02448_, _02445_);
  and _53925_ (_02450_, _01646_, _01861_);
  and _53926_ (_02451_, _01706_, _01875_);
  and _53927_ (_02452_, _01698_, _01829_);
  and _53928_ (_02453_, _01702_, _01877_);
  or _53929_ (_02454_, _02453_, _02452_);
  or _53930_ (_02455_, _02454_, _02451_);
  or _53931_ (_02456_, _02455_, _02450_);
  and _53932_ (_02457_, _01654_, _01842_);
  and _53933_ (_02458_, _01712_, _01866_);
  or _53934_ (_02459_, _02458_, _02457_);
  or _53935_ (_02460_, _02459_, _02456_);
  or _53936_ (_02461_, _02460_, _02449_);
  or _53937_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02461_, _02436_);
  and _53938_ (_02462_, _01694_, _01920_);
  and _53939_ (_02463_, _01712_, _01914_);
  and _53940_ (_02464_, _01641_, _01905_);
  or _53941_ (_02466_, _02464_, _02463_);
  or _53942_ (_02467_, _02466_, _02462_);
  and _53943_ (_02468_, _01660_, _01902_);
  and _53944_ (_02469_, _01664_, _01927_);
  and _53945_ (_02470_, _01671_, _01898_);
  or _53946_ (_02471_, _02470_, _02469_);
  and _53947_ (_02472_, _01667_, _01922_);
  and _53948_ (_02473_, _01675_, _01890_);
  or _53949_ (_02474_, _02473_, _02472_);
  or _53950_ (_02475_, _02474_, _02471_);
  or _53951_ (_02476_, _02475_, _02468_);
  and _53952_ (_02477_, _01687_, _01908_);
  and _53953_ (_02478_, _01683_, _01896_);
  or _53954_ (_02479_, _02478_, _02477_);
  or _53955_ (_02480_, _02479_, _02476_);
  and _53956_ (_02481_, _01654_, _01888_);
  and _53957_ (_02482_, _01715_, _01885_);
  or _53958_ (_02483_, _02482_, _02481_);
  and _53959_ (_02484_, _01646_, _01925_);
  and _53960_ (_02485_, _01702_, _01929_);
  and _53961_ (_02486_, _01698_, _01931_);
  and _53962_ (_02487_, _01706_, _01912_);
  or _53963_ (_02488_, _02487_, _02486_);
  or _53964_ (_02489_, _02488_, _02485_);
  or _53965_ (_02490_, _02489_, _02484_);
  or _53966_ (_02491_, _02490_, _02483_);
  or _53967_ (_02492_, _02491_, _02480_);
  or _53968_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02492_, _02467_);
  and _53969_ (_02493_, _01654_, _01952_);
  and _53970_ (_02494_, _01715_, _01941_);
  and _53971_ (_02495_, _01641_, _01966_);
  or _53972_ (_02496_, _02495_, _02494_);
  or _53973_ (_02497_, _02496_, _02493_);
  and _53974_ (_02498_, _01660_, _01978_);
  and _53975_ (_02499_, _01687_, _01969_);
  or _53976_ (_02500_, _02499_, _02498_);
  and _53977_ (_02501_, _01683_, _01962_);
  and _53978_ (_02502_, _01667_, _01954_);
  and _53979_ (_02503_, _01671_, _01960_);
  or _53980_ (_02504_, _02503_, _02502_);
  and _53981_ (_02505_, _01664_, _01944_);
  and _53982_ (_02506_, _01675_, _01980_);
  or _53983_ (_02507_, _02506_, _02505_);
  or _53984_ (_02508_, _02507_, _02504_);
  or _53985_ (_02509_, _02508_, _02501_);
  or _53986_ (_02510_, _02509_, _02500_);
  and _53987_ (_02511_, _01712_, _01976_);
  and _53988_ (_02512_, _01698_, _01946_);
  and _53989_ (_02513_, _01702_, _01989_);
  and _53990_ (_02514_, _01706_, _01986_);
  or _53991_ (_02515_, _02514_, _02513_);
  or _53992_ (_02516_, _02515_, _02512_);
  or _53993_ (_02517_, _02516_, _02511_);
  and _53994_ (_02518_, _01694_, _01983_);
  and _53995_ (_02519_, _01646_, _01971_);
  or _53996_ (_02520_, _02519_, _02518_);
  or _53997_ (_02521_, _02520_, _02517_);
  or _53998_ (_02522_, _02521_, _02510_);
  or _53999_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02522_, _02497_);
  and _54000_ (_02523_, _01694_, _01997_);
  and _54001_ (_02524_, _01654_, _02000_);
  and _54002_ (_02525_, _01712_, _02019_);
  or _54003_ (_02526_, _02525_, _02524_);
  or _54004_ (_02527_, _02526_, _02523_);
  and _54005_ (_02528_, _01687_, _02013_);
  and _54006_ (_02529_, _01675_, _02002_);
  and _54007_ (_02530_, _01671_, _02008_);
  or _54008_ (_02531_, _02530_, _02529_);
  and _54009_ (_02532_, _01667_, _02030_);
  and _54010_ (_02533_, _01664_, _02036_);
  or _54011_ (_02534_, _02533_, _02532_);
  or _54012_ (_02535_, _02534_, _02531_);
  or _54013_ (_02536_, _02535_, _02528_);
  and _54014_ (_02537_, _01660_, _02026_);
  and _54015_ (_02538_, _01683_, _02024_);
  or _54016_ (_02539_, _02538_, _02537_);
  or _54017_ (_02540_, _02539_, _02536_);
  and _54018_ (_02541_, _01641_, _02010_);
  and _54019_ (_02542_, _01646_, _02046_);
  or _54020_ (_02543_, _02542_, _02541_);
  and _54021_ (_02544_, _01715_, _02043_);
  and _54022_ (_02545_, _01702_, _02034_);
  and _54023_ (_02546_, _01706_, _02017_);
  and _54024_ (_02547_, _01698_, _02032_);
  or _54025_ (_02548_, _02547_, _02546_);
  or _54026_ (_02549_, _02548_, _02545_);
  or _54027_ (_02550_, _02549_, _02544_);
  or _54028_ (_02551_, _02550_, _02543_);
  or _54029_ (_02552_, _02551_, _02540_);
  or _54030_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02552_, _02527_);
  and _54031_ (_02553_, _01641_, _02071_);
  and _54032_ (_02554_, _01646_, _02081_);
  and _54033_ (_02555_, _01694_, _02095_);
  or _54034_ (_02556_, _02555_, _02554_);
  or _54035_ (_02557_, _02556_, _02553_);
  and _54036_ (_02558_, _01687_, _02079_);
  and _54037_ (_02559_, _01660_, _02091_);
  or _54038_ (_02560_, _02559_, _02558_);
  and _54039_ (_02561_, _01683_, _02073_);
  and _54040_ (_02562_, _01675_, _02088_);
  and _54041_ (_02563_, _01671_, _02075_);
  or _54042_ (_02564_, _02563_, _02562_);
  and _54043_ (_02565_, _01667_, _02064_);
  and _54044_ (_02566_, _01664_, _02056_);
  or _54045_ (_02567_, _02566_, _02565_);
  or _54046_ (_02568_, _02567_, _02564_);
  or _54047_ (_02569_, _02568_, _02561_);
  or _54048_ (_02570_, _02569_, _02560_);
  and _54049_ (_02571_, _01715_, _02060_);
  and _54050_ (_02572_, _01712_, _02086_);
  or _54051_ (_02573_, _02572_, _02571_);
  and _54052_ (_02574_, _01654_, _02066_);
  and _54053_ (_02575_, _01706_, _02098_);
  and _54054_ (_02576_, _01702_, _02101_);
  and _54055_ (_02577_, _01698_, _02053_);
  or _54056_ (_02578_, _02577_, _02576_);
  or _54057_ (_02579_, _02578_, _02575_);
  or _54058_ (_02580_, _02579_, _02574_);
  or _54059_ (_02581_, _02580_, _02573_);
  or _54060_ (_02582_, _02581_, _02570_);
  or _54061_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02582_, _02557_);
  and _54062_ (_02583_, _01654_, _02120_);
  and _54063_ (_02584_, _01646_, _02136_);
  and _54064_ (_02585_, _01715_, _02109_);
  or _54065_ (_02586_, _02585_, _02584_);
  or _54066_ (_02587_, _02586_, _02583_);
  and _54067_ (_02588_, _01660_, _02145_);
  and _54068_ (_02589_, _01675_, _02147_);
  and _54069_ (_02590_, _01671_, _02126_);
  or _54070_ (_02591_, _02590_, _02589_);
  and _54071_ (_02592_, _01667_, _02122_);
  and _54072_ (_02593_, _01664_, _02112_);
  or _54073_ (_02594_, _02593_, _02592_);
  or _54074_ (_02595_, _02594_, _02591_);
  or _54075_ (_02596_, _02595_, _02588_);
  and _54076_ (_02597_, _01687_, _02134_);
  and _54077_ (_02598_, _01683_, _02128_);
  or _54078_ (_02599_, _02598_, _02597_);
  or _54079_ (_02600_, _02599_, _02596_);
  and _54080_ (_02601_, _01712_, _02142_);
  and _54081_ (_02602_, _01702_, _02157_);
  and _54082_ (_02603_, _01706_, _02154_);
  and _54083_ (_02604_, _01698_, _02114_);
  or _54084_ (_02605_, _02604_, _02603_);
  or _54085_ (_02606_, _02605_, _02602_);
  or _54086_ (_02607_, _02606_, _02601_);
  and _54087_ (_02608_, _01641_, _02131_);
  and _54088_ (_02609_, _01694_, _02151_);
  or _54089_ (_02610_, _02609_, _02608_);
  or _54090_ (_02611_, _02610_, _02607_);
  or _54091_ (_02612_, _02611_, _02600_);
  or _54092_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02612_, _02587_);
  and _54093_ (_02613_, _01654_, _02177_);
  and _54094_ (_02614_, _01646_, _02191_);
  and _54095_ (_02615_, _01715_, _02172_);
  or _54096_ (_02616_, _02615_, _02614_);
  or _54097_ (_02617_, _02616_, _02613_);
  and _54098_ (_02618_, _01660_, _02203_);
  and _54099_ (_02619_, _01675_, _02201_);
  and _54100_ (_02620_, _01671_, _02185_);
  or _54101_ (_02621_, _02620_, _02619_);
  and _54102_ (_02622_, _01667_, _02207_);
  and _54103_ (_02623_, _01664_, _02168_);
  or _54104_ (_02624_, _02623_, _02622_);
  or _54105_ (_02625_, _02624_, _02621_);
  or _54106_ (_02626_, _02625_, _02618_);
  and _54107_ (_02627_, _01687_, _02189_);
  and _54108_ (_02628_, _01683_, _02183_);
  or _54109_ (_02629_, _02628_, _02627_);
  or _54110_ (_02630_, _02629_, _02626_);
  and _54111_ (_02631_, _01712_, _02198_);
  and _54112_ (_02632_, _01702_, _02213_);
  and _54113_ (_02633_, _01706_, _02210_);
  and _54114_ (_02634_, _01698_, _02165_);
  or _54115_ (_02635_, _02634_, _02633_);
  or _54116_ (_02636_, _02635_, _02632_);
  or _54117_ (_02637_, _02636_, _02631_);
  and _54118_ (_02638_, _01641_, _02181_);
  and _54119_ (_02639_, _01694_, _02175_);
  or _54120_ (_02640_, _02639_, _02638_);
  or _54121_ (_02641_, _02640_, _02637_);
  or _54122_ (_02642_, _02641_, _02630_);
  or _54123_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02642_, _02617_);
  and _54124_ (_02643_, _01712_, _01842_);
  and _54125_ (_02644_, _01694_, _01875_);
  and _54126_ (_02645_, _01646_, _01840_);
  or _54127_ (_02646_, _02645_, _02644_);
  or _54128_ (_02647_, _02646_, _02643_);
  and _54129_ (_02648_, _01687_, _01850_);
  and _54130_ (_02649_, _01667_, _01877_);
  and _54131_ (_02650_, _01671_, _01861_);
  or _54132_ (_02651_, _02650_, _02649_);
  and _54133_ (_02652_, _01664_, _01836_);
  and _54134_ (_02653_, _01675_, _01870_);
  or _54135_ (_02654_, _02653_, _02652_);
  or _54136_ (_02655_, _02654_, _02651_);
  or _54137_ (_02656_, _02655_, _02648_);
  and _54138_ (_02657_, _01683_, _01848_);
  and _54139_ (_02658_, _01660_, _01853_);
  or _54140_ (_02659_, _02658_, _02657_);
  or _54141_ (_02661_, _02659_, _02656_);
  and _54142_ (_02662_, _01715_, _01868_);
  and _54143_ (_02663_, _01698_, _01866_);
  and _54144_ (_02664_, _01706_, _01829_);
  and _54145_ (_02665_, _01702_, _01832_);
  or _54146_ (_02666_, _02665_, _02664_);
  or _54147_ (_02667_, _02666_, _02663_);
  or _54148_ (_02668_, _02667_, _02662_);
  and _54149_ (_02669_, _01641_, _01873_);
  and _54150_ (_02670_, _01654_, _01858_);
  or _54151_ (_02671_, _02670_, _02669_);
  or _54152_ (_02672_, _02671_, _02668_);
  or _54153_ (_02673_, _02672_, _02661_);
  or _54154_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _02673_, _02647_);
  and _54155_ (_02674_, _01712_, _01888_);
  and _54156_ (_02675_, _01694_, _01912_);
  and _54157_ (_02676_, _01646_, _01922_);
  or _54158_ (_02677_, _02676_, _02675_);
  or _54159_ (_02678_, _02677_, _02674_);
  and _54160_ (_02679_, _01687_, _01896_);
  and _54161_ (_02680_, _01667_, _01929_);
  and _54162_ (_02681_, _01671_, _01925_);
  or _54163_ (_02682_, _02681_, _02680_);
  and _54164_ (_02683_, _01664_, _01885_);
  and _54165_ (_02684_, _01675_, _01902_);
  or _54166_ (_02685_, _02684_, _02683_);
  or _54167_ (_02686_, _02685_, _02682_);
  or _54168_ (_02687_, _02686_, _02679_);
  and _54169_ (_02688_, _01683_, _01905_);
  and _54170_ (_02689_, _01660_, _01898_);
  or _54171_ (_02690_, _02689_, _02688_);
  or _54172_ (_02691_, _02690_, _02687_);
  and _54173_ (_02692_, _01715_, _01890_);
  and _54174_ (_02693_, _01698_, _01914_);
  and _54175_ (_02694_, _01706_, _01931_);
  and _54176_ (_02695_, _01702_, _01927_);
  or _54177_ (_02696_, _02695_, _02694_);
  or _54178_ (_02697_, _02696_, _02693_);
  or _54179_ (_02698_, _02697_, _02692_);
  and _54180_ (_02699_, _01641_, _01920_);
  and _54181_ (_02700_, _01654_, _01908_);
  or _54182_ (_02701_, _02700_, _02699_);
  or _54183_ (_02702_, _02701_, _02698_);
  or _54184_ (_02703_, _02702_, _02691_);
  or _54185_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02703_, _02678_);
  and _54186_ (_02704_, _01712_, _01952_);
  and _54187_ (_02705_, _01694_, _01986_);
  and _54188_ (_02706_, _01646_, _01954_);
  or _54189_ (_02707_, _02706_, _02705_);
  or _54190_ (_02708_, _02707_, _02704_);
  and _54191_ (_02709_, _01660_, _01960_);
  and _54192_ (_02710_, _01667_, _01989_);
  and _54193_ (_02711_, _01671_, _01971_);
  or _54194_ (_02712_, _02711_, _02710_);
  and _54195_ (_02713_, _01664_, _01941_);
  and _54196_ (_02714_, _01675_, _01978_);
  or _54197_ (_02715_, _02714_, _02713_);
  or _54198_ (_02716_, _02715_, _02712_);
  or _54199_ (_02717_, _02716_, _02709_);
  and _54200_ (_02718_, _01683_, _01966_);
  and _54201_ (_02719_, _01687_, _01962_);
  or _54202_ (_02720_, _02719_, _02718_);
  or _54203_ (_02721_, _02720_, _02717_);
  and _54204_ (_02722_, _01715_, _01980_);
  and _54205_ (_02723_, _01698_, _01976_);
  and _54206_ (_02724_, _01706_, _01946_);
  and _54207_ (_02725_, _01702_, _01944_);
  or _54208_ (_02726_, _02725_, _02724_);
  or _54209_ (_02727_, _02726_, _02723_);
  or _54210_ (_02728_, _02727_, _02722_);
  and _54211_ (_02729_, _01641_, _01983_);
  and _54212_ (_02730_, _01654_, _01969_);
  or _54213_ (_02731_, _02730_, _02729_);
  or _54214_ (_02732_, _02731_, _02728_);
  or _54215_ (_02733_, _02732_, _02721_);
  or _54216_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02733_, _02708_);
  and _54217_ (_02734_, _01646_, _02030_);
  and _54218_ (_02735_, _01694_, _02017_);
  and _54219_ (_02736_, _01641_, _01997_);
  or _54220_ (_02737_, _02736_, _02735_);
  or _54221_ (_02738_, _02737_, _02734_);
  and _54222_ (_02739_, _01687_, _02024_);
  and _54223_ (_02740_, _01667_, _02034_);
  and _54224_ (_02741_, _01671_, _02046_);
  or _54225_ (_02742_, _02741_, _02740_);
  and _54226_ (_02743_, _01664_, _02043_);
  and _54227_ (_02744_, _01675_, _02026_);
  or _54228_ (_02745_, _02744_, _02743_);
  or _54229_ (_02746_, _02745_, _02742_);
  or _54230_ (_02747_, _02746_, _02739_);
  and _54231_ (_02748_, _01683_, _02010_);
  and _54232_ (_02749_, _01660_, _02008_);
  or _54233_ (_02750_, _02749_, _02748_);
  or _54234_ (_02751_, _02750_, _02747_);
  and _54235_ (_02752_, _01712_, _02000_);
  and _54236_ (_02753_, _01698_, _02019_);
  and _54237_ (_02754_, _01706_, _02032_);
  and _54238_ (_02755_, _01702_, _02036_);
  or _54239_ (_02756_, _02755_, _02754_);
  or _54240_ (_02757_, _02756_, _02753_);
  or _54241_ (_02758_, _02757_, _02752_);
  and _54242_ (_02759_, _01715_, _02002_);
  and _54243_ (_02760_, _01654_, _02013_);
  or _54244_ (_02761_, _02760_, _02759_);
  or _54245_ (_02762_, _02761_, _02758_);
  or _54246_ (_02763_, _02762_, _02751_);
  or _54247_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02763_, _02738_);
  and _54248_ (_02764_, _01646_, _02064_);
  and _54249_ (_02765_, _01694_, _02098_);
  and _54250_ (_02766_, _01641_, _02095_);
  or _54251_ (_02767_, _02766_, _02765_);
  or _54252_ (_02768_, _02767_, _02764_);
  and _54253_ (_02769_, _01660_, _02075_);
  and _54254_ (_02770_, _01667_, _02101_);
  and _54255_ (_02771_, _01671_, _02081_);
  or _54256_ (_02772_, _02771_, _02770_);
  and _54257_ (_02773_, _01664_, _02060_);
  and _54258_ (_02774_, _01675_, _02091_);
  or _54259_ (_02775_, _02774_, _02773_);
  or _54260_ (_02776_, _02775_, _02772_);
  or _54261_ (_02777_, _02776_, _02769_);
  and _54262_ (_02778_, _01683_, _02071_);
  and _54263_ (_02779_, _01687_, _02073_);
  or _54264_ (_02780_, _02779_, _02778_);
  or _54265_ (_02781_, _02780_, _02777_);
  and _54266_ (_02782_, _01712_, _02066_);
  and _54267_ (_02783_, _01698_, _02086_);
  and _54268_ (_02784_, _01706_, _02053_);
  and _54269_ (_02785_, _01702_, _02056_);
  or _54270_ (_02786_, _02785_, _02784_);
  or _54271_ (_02787_, _02786_, _02783_);
  or _54272_ (_02788_, _02787_, _02782_);
  and _54273_ (_02789_, _01715_, _02088_);
  and _54274_ (_02790_, _01654_, _02079_);
  or _54275_ (_02791_, _02790_, _02789_);
  or _54276_ (_02792_, _02791_, _02788_);
  or _54277_ (_02793_, _02792_, _02781_);
  or _54278_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02793_, _02768_);
  and _54279_ (_02794_, _01694_, _02154_);
  and _54280_ (_02795_, _01715_, _02147_);
  and _54281_ (_02796_, _01646_, _02122_);
  or _54282_ (_02797_, _02796_, _02795_);
  or _54283_ (_02798_, _02797_, _02794_);
  and _54284_ (_02799_, _01660_, _02126_);
  and _54285_ (_02800_, _01671_, _02136_);
  and _54286_ (_02801_, _01675_, _02145_);
  or _54287_ (_02802_, _02801_, _02800_);
  and _54288_ (_02803_, _01667_, _02157_);
  and _54289_ (_02804_, _01664_, _02109_);
  or _54290_ (_02805_, _02804_, _02803_);
  or _54291_ (_02806_, _02805_, _02802_);
  or _54292_ (_02807_, _02806_, _02799_);
  and _54293_ (_02808_, _01683_, _02131_);
  and _54294_ (_02809_, _01687_, _02128_);
  or _54295_ (_02810_, _02809_, _02808_);
  or _54296_ (_02811_, _02810_, _02807_);
  and _54297_ (_02812_, _01641_, _02151_);
  and _54298_ (_02813_, _01698_, _02142_);
  and _54299_ (_02814_, _01702_, _02112_);
  and _54300_ (_02815_, _01706_, _02114_);
  or _54301_ (_02816_, _02815_, _02814_);
  or _54302_ (_02817_, _02816_, _02813_);
  or _54303_ (_02818_, _02817_, _02812_);
  and _54304_ (_02819_, _01712_, _02120_);
  and _54305_ (_02820_, _01654_, _02134_);
  or _54306_ (_02821_, _02820_, _02819_);
  or _54307_ (_02822_, _02821_, _02818_);
  or _54308_ (_02823_, _02822_, _02811_);
  or _54309_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02823_, _02798_);
  and _54310_ (_02824_, _01712_, _02177_);
  and _54311_ (_02825_, _01694_, _02210_);
  and _54312_ (_02826_, _01641_, _02175_);
  or _54313_ (_02827_, _02826_, _02825_);
  or _54314_ (_02828_, _02827_, _02824_);
  and _54315_ (_02829_, _01687_, _02183_);
  and _54316_ (_02830_, _01667_, _02213_);
  and _54317_ (_02831_, _01671_, _02191_);
  or _54318_ (_02832_, _02831_, _02830_);
  and _54319_ (_02833_, _01664_, _02172_);
  and _54320_ (_02834_, _01675_, _02203_);
  or _54321_ (_02835_, _02834_, _02833_);
  or _54322_ (_02836_, _02835_, _02832_);
  or _54323_ (_02837_, _02836_, _02829_);
  and _54324_ (_02838_, _01683_, _02181_);
  and _54325_ (_02839_, _01660_, _02185_);
  or _54326_ (_02840_, _02839_, _02838_);
  or _54327_ (_02841_, _02840_, _02837_);
  and _54328_ (_02842_, _01715_, _02201_);
  and _54329_ (_02843_, _01698_, _02198_);
  and _54330_ (_02844_, _01706_, _02165_);
  and _54331_ (_02845_, _01702_, _02168_);
  or _54332_ (_02846_, _02845_, _02844_);
  or _54333_ (_02847_, _02846_, _02843_);
  or _54334_ (_02848_, _02847_, _02842_);
  and _54335_ (_02849_, _01646_, _02207_);
  and _54336_ (_02850_, _01654_, _02189_);
  or _54337_ (_02851_, _02850_, _02849_);
  or _54338_ (_02852_, _02851_, _02848_);
  or _54339_ (_02853_, _02852_, _02841_);
  or _54340_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02853_, _02828_);
  nand _54341_ (_02855_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not _54342_ (_02856_, \oc8051_golden_model_1.PC [3]);
  or _54343_ (_02857_, \oc8051_golden_model_1.PC [2], _02856_);
  or _54344_ (_02858_, _02857_, _02855_);
  or _54345_ (_02859_, _02858_, _42111_);
  not _54346_ (_02860_, \oc8051_golden_model_1.PC [1]);
  or _54347_ (_02861_, _02860_, \oc8051_golden_model_1.PC [0]);
  or _54348_ (_02862_, _02861_, _02857_);
  or _54349_ (_02863_, _02862_, _42070_);
  and _54350_ (_02864_, _02863_, _02859_);
  not _54351_ (_02865_, \oc8051_golden_model_1.PC [2]);
  or _54352_ (_02866_, _02865_, \oc8051_golden_model_1.PC [3]);
  or _54353_ (_02867_, _02866_, _02855_);
  or _54354_ (_02868_, _02867_, _41947_);
  or _54355_ (_02869_, _02866_, _02861_);
  or _54356_ (_02870_, _02869_, _41906_);
  and _54357_ (_02871_, _02870_, _02868_);
  and _54358_ (_02872_, _02871_, _02864_);
  nand _54359_ (_02873_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _54360_ (_02874_, _02873_, _02855_);
  or _54361_ (_02875_, _02874_, _42275_);
  or _54362_ (_02876_, _02873_, _02861_);
  or _54363_ (_02877_, _02876_, _42234_);
  and _54364_ (_02878_, _02877_, _02875_);
  or _54365_ (_02879_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _54366_ (_02880_, _02879_, _02855_);
  or _54367_ (_02881_, _02880_, _41783_);
  or _54368_ (_02882_, _02879_, _02861_);
  or _54369_ (_02883_, _02882_, _41734_);
  and _54370_ (_02884_, _02883_, _02881_);
  and _54371_ (_02885_, _02884_, _02878_);
  and _54372_ (_02886_, _02885_, _02872_);
  not _54373_ (_02887_, \oc8051_golden_model_1.PC [0]);
  or _54374_ (_02888_, \oc8051_golden_model_1.PC [1], _02887_);
  or _54375_ (_02889_, _02888_, _02873_);
  or _54376_ (_02890_, _02889_, _42193_);
  or _54377_ (_02891_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or _54378_ (_02892_, _02891_, _02873_);
  or _54379_ (_02893_, _02892_, _42152_);
  and _54380_ (_02894_, _02893_, _02890_);
  or _54381_ (_02895_, _02879_, _02891_);
  or _54382_ (_02896_, _02895_, _41645_);
  or _54383_ (_02897_, _02879_, _02888_);
  or _54384_ (_02898_, _02897_, _41686_);
  and _54385_ (_02899_, _02898_, _02896_);
  and _54386_ (_02900_, _02899_, _02894_);
  or _54387_ (_02901_, _02888_, _02857_);
  or _54388_ (_02902_, _02901_, _42029_);
  or _54389_ (_02903_, _02891_, _02857_);
  or _54390_ (_02904_, _02903_, _41988_);
  and _54391_ (_02905_, _02904_, _02902_);
  or _54392_ (_02906_, _02888_, _02866_);
  or _54393_ (_02907_, _02906_, _41865_);
  or _54394_ (_02908_, _02891_, _02866_);
  or _54395_ (_02909_, _02908_, _41824_);
  and _54396_ (_02910_, _02909_, _02907_);
  and _54397_ (_02911_, _02910_, _02905_);
  and _54398_ (_02912_, _02911_, _02900_);
  and _54399_ (_02913_, _02912_, _02886_);
  or _54400_ (_02914_, _02858_, _42076_);
  or _54401_ (_02915_, _02862_, _42035_);
  and _54402_ (_02916_, _02915_, _02914_);
  or _54403_ (_02917_, _02867_, _41912_);
  or _54404_ (_02918_, _02869_, _41871_);
  and _54405_ (_02919_, _02918_, _02917_);
  and _54406_ (_02920_, _02919_, _02916_);
  or _54407_ (_02921_, _02874_, _42240_);
  or _54408_ (_02922_, _02876_, _42199_);
  and _54409_ (_02923_, _02922_, _02921_);
  or _54410_ (_02924_, _02880_, _41740_);
  or _54411_ (_02925_, _02882_, _41692_);
  and _54412_ (_02926_, _02925_, _02924_);
  and _54413_ (_02927_, _02926_, _02923_);
  and _54414_ (_02928_, _02927_, _02920_);
  or _54415_ (_02929_, _02889_, _42158_);
  or _54416_ (_02930_, _02892_, _42117_);
  and _54417_ (_02931_, _02930_, _02929_);
  or _54418_ (_02932_, _02895_, _41610_);
  or _54419_ (_02933_, _02897_, _41651_);
  and _54420_ (_02934_, _02933_, _02932_);
  and _54421_ (_02935_, _02934_, _02931_);
  or _54422_ (_02936_, _02901_, _41994_);
  or _54423_ (_02937_, _02903_, _41953_);
  and _54424_ (_02938_, _02937_, _02936_);
  or _54425_ (_02939_, _02906_, _41830_);
  or _54426_ (_02940_, _02908_, _41789_);
  and _54427_ (_02941_, _02940_, _02939_);
  and _54428_ (_02942_, _02941_, _02938_);
  and _54429_ (_02943_, _02942_, _02935_);
  and _54430_ (_02944_, _02943_, _02928_);
  and _54431_ (_02945_, _02944_, _02913_);
  or _54432_ (_02946_, _02858_, _42101_);
  or _54433_ (_02947_, _02862_, _42060_);
  and _54434_ (_02948_, _02947_, _02946_);
  or _54435_ (_02949_, _02867_, _41937_);
  or _54436_ (_02950_, _02869_, _41896_);
  and _54437_ (_02951_, _02950_, _02949_);
  and _54438_ (_02952_, _02951_, _02948_);
  or _54439_ (_02953_, _02874_, _42265_);
  or _54440_ (_02954_, _02876_, _42224_);
  and _54441_ (_02955_, _02954_, _02953_);
  or _54442_ (_02956_, _02880_, _41773_);
  or _54443_ (_02957_, _02882_, _41724_);
  and _54444_ (_02958_, _02957_, _02956_);
  and _54445_ (_02959_, _02958_, _02955_);
  and _54446_ (_02960_, _02959_, _02952_);
  or _54447_ (_02961_, _02889_, _42183_);
  or _54448_ (_02962_, _02892_, _42142_);
  and _54449_ (_02963_, _02962_, _02961_);
  or _54450_ (_02964_, _02895_, _41635_);
  or _54451_ (_02965_, _02897_, _41676_);
  and _54452_ (_02966_, _02965_, _02964_);
  and _54453_ (_02967_, _02966_, _02963_);
  or _54454_ (_02968_, _02901_, _42019_);
  or _54455_ (_02969_, _02903_, _41978_);
  and _54456_ (_02970_, _02969_, _02968_);
  or _54457_ (_02971_, _02906_, _41855_);
  or _54458_ (_02972_, _02908_, _41814_);
  and _54459_ (_02973_, _02972_, _02971_);
  and _54460_ (_02974_, _02973_, _02970_);
  and _54461_ (_02975_, _02974_, _02967_);
  and _54462_ (_02976_, _02975_, _02960_);
  or _54463_ (_02977_, _02858_, _42106_);
  or _54464_ (_02978_, _02862_, _42065_);
  and _54465_ (_02979_, _02978_, _02977_);
  or _54466_ (_02980_, _02867_, _41942_);
  or _54467_ (_02981_, _02869_, _41901_);
  and _54468_ (_02982_, _02981_, _02980_);
  and _54469_ (_02983_, _02982_, _02979_);
  or _54470_ (_02984_, _02874_, _42270_);
  or _54471_ (_02985_, _02876_, _42229_);
  and _54472_ (_02986_, _02985_, _02984_);
  or _54473_ (_02987_, _02880_, _41778_);
  or _54474_ (_02988_, _02882_, _41729_);
  and _54475_ (_02989_, _02988_, _02987_);
  and _54476_ (_02990_, _02989_, _02986_);
  and _54477_ (_02991_, _02990_, _02983_);
  or _54478_ (_02992_, _02889_, _42188_);
  or _54479_ (_02993_, _02892_, _42147_);
  and _54480_ (_02994_, _02993_, _02992_);
  or _54481_ (_02995_, _02895_, _41640_);
  or _54482_ (_02996_, _02897_, _41681_);
  and _54483_ (_02997_, _02996_, _02995_);
  and _54484_ (_02998_, _02997_, _02994_);
  or _54485_ (_02999_, _02901_, _42024_);
  or _54486_ (_03000_, _02903_, _41983_);
  and _54487_ (_03001_, _03000_, _02999_);
  or _54488_ (_03002_, _02906_, _41860_);
  or _54489_ (_03003_, _02908_, _41819_);
  and _54490_ (_03004_, _03003_, _03002_);
  and _54491_ (_03005_, _03004_, _03001_);
  and _54492_ (_03006_, _03005_, _02998_);
  nand _54493_ (_03007_, _03006_, _02991_);
  or _54494_ (_03008_, _03007_, _02976_);
  not _54495_ (_03009_, _03008_);
  and _54496_ (_03010_, _03009_, _02945_);
  or _54497_ (_03011_, _02858_, _42081_);
  or _54498_ (_03012_, _02862_, _42040_);
  and _54499_ (_03013_, _03012_, _03011_);
  or _54500_ (_03014_, _02867_, _41917_);
  or _54501_ (_03016_, _02869_, _41876_);
  and _54502_ (_03017_, _03016_, _03014_);
  and _54503_ (_03018_, _03017_, _03013_);
  or _54504_ (_03019_, _02874_, _42245_);
  or _54505_ (_03020_, _02876_, _42204_);
  and _54506_ (_03021_, _03020_, _03019_);
  or _54507_ (_03022_, _02880_, _41749_);
  or _54508_ (_03023_, _02882_, _41697_);
  and _54509_ (_03024_, _03023_, _03022_);
  and _54510_ (_03025_, _03024_, _03021_);
  and _54511_ (_03027_, _03025_, _03018_);
  or _54512_ (_03028_, _02889_, _42163_);
  or _54513_ (_03029_, _02892_, _42122_);
  and _54514_ (_03030_, _03029_, _03028_);
  or _54515_ (_03031_, _02895_, _41615_);
  or _54516_ (_03032_, _02897_, _41656_);
  and _54517_ (_03033_, _03032_, _03031_);
  and _54518_ (_03034_, _03033_, _03030_);
  or _54519_ (_03035_, _02901_, _41999_);
  or _54520_ (_03036_, _02903_, _41958_);
  and _54521_ (_03037_, _03036_, _03035_);
  or _54522_ (_03038_, _02906_, _41835_);
  or _54523_ (_03039_, _02908_, _41794_);
  and _54524_ (_03040_, _03039_, _03038_);
  and _54525_ (_03041_, _03040_, _03037_);
  and _54526_ (_03042_, _03041_, _03034_);
  and _54527_ (_03043_, _03042_, _03027_);
  or _54528_ (_03044_, _02858_, _42086_);
  or _54529_ (_03045_, _02862_, _42045_);
  and _54530_ (_03046_, _03045_, _03044_);
  or _54531_ (_03048_, _02867_, _41922_);
  or _54532_ (_03049_, _02869_, _41881_);
  and _54533_ (_03050_, _03049_, _03048_);
  and _54534_ (_03051_, _03050_, _03046_);
  or _54535_ (_03052_, _02874_, _42250_);
  or _54536_ (_03053_, _02876_, _42209_);
  and _54537_ (_03054_, _03053_, _03052_);
  or _54538_ (_03055_, _02880_, _41758_);
  or _54539_ (_03056_, _02882_, _41706_);
  and _54540_ (_03057_, _03056_, _03055_);
  and _54541_ (_03059_, _03057_, _03054_);
  and _54542_ (_03060_, _03059_, _03051_);
  or _54543_ (_03061_, _02889_, _42168_);
  or _54544_ (_03062_, _02892_, _42127_);
  and _54545_ (_03063_, _03062_, _03061_);
  or _54546_ (_03064_, _02895_, _41620_);
  or _54547_ (_03065_, _02897_, _41661_);
  and _54548_ (_03066_, _03065_, _03064_);
  and _54549_ (_03067_, _03066_, _03063_);
  or _54550_ (_03068_, _02901_, _42004_);
  or _54551_ (_03070_, _02903_, _41963_);
  and _54552_ (_03071_, _03070_, _03068_);
  or _54553_ (_03072_, _02906_, _41840_);
  or _54554_ (_03073_, _02908_, _41799_);
  and _54555_ (_03074_, _03073_, _03072_);
  and _54556_ (_03075_, _03074_, _03071_);
  and _54557_ (_03076_, _03075_, _03067_);
  nand _54558_ (_03077_, _03076_, _03060_);
  not _54559_ (_03078_, _03077_);
  and _54560_ (_03079_, _03078_, _03043_);
  or _54561_ (_03080_, _02858_, _42091_);
  or _54562_ (_03081_, _02862_, _42050_);
  and _54563_ (_03082_, _03081_, _03080_);
  or _54564_ (_03083_, _02867_, _41927_);
  or _54565_ (_03084_, _02869_, _41886_);
  and _54566_ (_03085_, _03084_, _03083_);
  and _54567_ (_03086_, _03085_, _03082_);
  or _54568_ (_03087_, _02874_, _42255_);
  or _54569_ (_03088_, _02876_, _42214_);
  and _54570_ (_03089_, _03088_, _03087_);
  or _54571_ (_03091_, _02880_, _41763_);
  or _54572_ (_03092_, _02882_, _41714_);
  and _54573_ (_03093_, _03092_, _03091_);
  and _54574_ (_03094_, _03093_, _03089_);
  and _54575_ (_03095_, _03094_, _03086_);
  or _54576_ (_03096_, _02889_, _42173_);
  or _54577_ (_03097_, _02892_, _42132_);
  and _54578_ (_03098_, _03097_, _03096_);
  or _54579_ (_03099_, _02895_, _41625_);
  or _54580_ (_03100_, _02897_, _41666_);
  and _54581_ (_03102_, _03100_, _03099_);
  and _54582_ (_03103_, _03102_, _03098_);
  or _54583_ (_03104_, _02901_, _42009_);
  or _54584_ (_03105_, _02903_, _41968_);
  and _54585_ (_03106_, _03105_, _03104_);
  or _54586_ (_03107_, _02906_, _41845_);
  or _54587_ (_03108_, _02908_, _41804_);
  and _54588_ (_03109_, _03108_, _03107_);
  and _54589_ (_03110_, _03109_, _03106_);
  and _54590_ (_03111_, _03110_, _03103_);
  nand _54591_ (_03113_, _03111_, _03095_);
  or _54592_ (_03114_, _02858_, _42096_);
  or _54593_ (_03115_, _02862_, _42055_);
  and _54594_ (_03116_, _03115_, _03114_);
  or _54595_ (_03117_, _02867_, _41932_);
  or _54596_ (_03118_, _02869_, _41891_);
  and _54597_ (_03119_, _03118_, _03117_);
  and _54598_ (_03120_, _03119_, _03116_);
  or _54599_ (_03121_, _02874_, _42260_);
  or _54600_ (_03122_, _02876_, _42219_);
  and _54601_ (_03124_, _03122_, _03121_);
  or _54602_ (_03125_, _02880_, _41768_);
  or _54603_ (_03126_, _02882_, _41719_);
  and _54604_ (_03127_, _03126_, _03125_);
  and _54605_ (_03128_, _03127_, _03124_);
  and _54606_ (_03129_, _03128_, _03120_);
  or _54607_ (_03130_, _02889_, _42178_);
  or _54608_ (_03131_, _02892_, _42137_);
  and _54609_ (_03132_, _03131_, _03130_);
  or _54610_ (_03133_, _02895_, _41630_);
  or _54611_ (_03135_, _02897_, _41671_);
  and _54612_ (_03136_, _03135_, _03133_);
  and _54613_ (_03137_, _03136_, _03132_);
  or _54614_ (_03138_, _02901_, _42014_);
  or _54615_ (_03139_, _02903_, _41973_);
  and _54616_ (_03140_, _03139_, _03138_);
  or _54617_ (_03141_, _02906_, _41850_);
  or _54618_ (_03142_, _02908_, _41809_);
  and _54619_ (_03143_, _03142_, _03141_);
  and _54620_ (_03144_, _03143_, _03140_);
  and _54621_ (_03146_, _03144_, _03137_);
  nand _54622_ (_03147_, _03146_, _03129_);
  or _54623_ (_03148_, _03147_, _03113_);
  not _54624_ (_03149_, _03148_);
  and _54625_ (_03150_, _03149_, _03079_);
  and _54626_ (_03151_, _03150_, _03010_);
  not _54627_ (_03152_, _03151_);
  and _54628_ (_03153_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _54629_ (_03154_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _54630_ (_03155_, _03154_, _03153_);
  or _54631_ (_03157_, _03077_, _03043_);
  or _54632_ (_03158_, _03157_, _03148_);
  not _54633_ (_03159_, _03158_);
  and _54634_ (_03160_, _03159_, _03010_);
  not _54635_ (_03161_, _03160_);
  nand _54636_ (_03162_, _02975_, _02960_);
  or _54637_ (_03163_, _03007_, _03162_);
  not _54638_ (_03164_, _03163_);
  and _54639_ (_03165_, _03164_, _02945_);
  and _54640_ (_03166_, _03165_, _03159_);
  and _54641_ (_03168_, _03006_, _02991_);
  or _54642_ (_03169_, _03168_, _03162_);
  not _54643_ (_03170_, _03169_);
  and _54644_ (_03171_, _03170_, _02945_);
  and _54645_ (_03172_, _03171_, _03159_);
  nor _54646_ (_03173_, _03172_, _03166_);
  and _54647_ (_03174_, _03173_, _03161_);
  or _54648_ (_03175_, _03168_, _02976_);
  not _54649_ (_03176_, _03175_);
  and _54650_ (_03177_, _03176_, _02945_);
  and _54651_ (_03179_, _03177_, _03159_);
  nand _54652_ (_03180_, _02912_, _02886_);
  and _54653_ (_03181_, _02944_, _03180_);
  and _54654_ (_03182_, _03181_, _03164_);
  and _54655_ (_03183_, _03182_, _03159_);
  nor _54656_ (_03184_, _03183_, _03179_);
  or _54657_ (_03185_, _02944_, _03180_);
  nor _54658_ (_03186_, _03185_, _03163_);
  and _54659_ (_03187_, _03186_, _03159_);
  and _54660_ (_03188_, _03181_, _03176_);
  and _54661_ (_03189_, _03188_, _03159_);
  nor _54662_ (_03190_, _03189_, _03187_);
  and _54663_ (_03191_, _03181_, _03009_);
  and _54664_ (_03192_, _03191_, _03159_);
  and _54665_ (_03193_, _03181_, _03170_);
  and _54666_ (_03194_, _03193_, _03159_);
  nor _54667_ (_03195_, _03194_, _03192_);
  and _54668_ (_03196_, _03195_, _03190_);
  and _54669_ (_03197_, _03196_, _03184_);
  and _54670_ (_03198_, _03197_, _03174_);
  or _54671_ (_03199_, _03175_, _03185_);
  or _54672_ (_03200_, _03199_, _03158_);
  or _54673_ (_03201_, _02944_, _02913_);
  or _54674_ (_03202_, _03201_, _03008_);
  or _54675_ (_03203_, _03202_, _03158_);
  and _54676_ (_03204_, _03203_, _03200_);
  or _54677_ (_03205_, _03201_, _03163_);
  or _54678_ (_03206_, _03205_, _03158_);
  or _54679_ (_03207_, _03201_, _03169_);
  or _54680_ (_03208_, _03207_, _03158_);
  and _54681_ (_03209_, _03208_, _03206_);
  or _54682_ (_03210_, _03201_, _03175_);
  or _54683_ (_03211_, _03210_, _03158_);
  or _54684_ (_03212_, _03185_, _03169_);
  or _54685_ (_03213_, _03212_, _03158_);
  and _54686_ (_03214_, _03213_, _03211_);
  and _54687_ (_03215_, _03214_, _03209_);
  and _54688_ (_03216_, _03215_, _03204_);
  not _54689_ (_03217_, _03157_);
  not _54690_ (_03218_, _03147_);
  and _54691_ (_03219_, _03218_, _03113_);
  and _54692_ (_03220_, _03219_, _03217_);
  and _54693_ (_03221_, _03220_, _03186_);
  nor _54694_ (_03222_, _03185_, _03008_);
  and _54695_ (_03223_, _03222_, _03159_);
  nor _54696_ (_03224_, _03223_, _03221_);
  and _54697_ (_03225_, _03224_, _03216_);
  and _54698_ (_03226_, _03225_, _03198_);
  or _54699_ (_03227_, _03226_, _03155_);
  or _54700_ (_03228_, _03078_, _03043_);
  or _54701_ (_03229_, _03228_, _03148_);
  not _54702_ (_03230_, _03229_);
  and _54703_ (_03231_, _03230_, _03186_);
  not _54704_ (_03232_, _03231_);
  not _54705_ (_03233_, \oc8051_golden_model_1.ACC [1]);
  and _54706_ (_03234_, _02888_, _02861_);
  nor _54707_ (_03235_, _03234_, _03233_);
  and _54708_ (_03236_, \oc8051_golden_model_1.ACC [0], _02887_);
  and _54709_ (_03237_, _03234_, _03233_);
  nor _54710_ (_03238_, _03237_, _03235_);
  and _54711_ (_03239_, _03238_, _03236_);
  nor _54712_ (_03240_, _03239_, _03235_);
  nor _54713_ (_03241_, _02855_, _02865_);
  and _54714_ (_03242_, _02855_, _02865_);
  nor _54715_ (_03243_, _03242_, _03241_);
  and _54716_ (_03244_, _03243_, \oc8051_golden_model_1.ACC [2]);
  nor _54717_ (_03245_, _03243_, \oc8051_golden_model_1.ACC [2]);
  nor _54718_ (_03246_, _03245_, _03244_);
  not _54719_ (_03247_, _03246_);
  and _54720_ (_03248_, _03247_, _03240_);
  nor _54721_ (_03249_, _03247_, _03240_);
  nor _54722_ (_03250_, _03249_, _03248_);
  nor _54723_ (_03251_, _03250_, _03232_);
  and _54724_ (_03252_, _03232_, _03224_);
  not _54725_ (_03253_, _03222_);
  or _54726_ (_03254_, _03229_, _03253_);
  and _54727_ (_03255_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and _54728_ (_03256_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _54729_ (_03257_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _54730_ (_03258_, _03257_, _03255_);
  and _54731_ (_03259_, _03258_, _03256_);
  nor _54732_ (_03260_, _03259_, _03255_);
  and _54733_ (_03261_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _54734_ (_03262_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _54735_ (_03263_, _03262_, _03261_);
  not _54736_ (_03264_, _03263_);
  nor _54737_ (_03265_, _03264_, _03260_);
  and _54738_ (_03266_, _03264_, _03260_);
  nor _54739_ (_03267_, _03266_, _03265_);
  or _54740_ (_03268_, _03267_, _03254_);
  not _54741_ (_03270_, _03243_);
  and _54742_ (_03271_, _03254_, _03270_);
  nand _54743_ (_03272_, _03271_, _03216_);
  nand _54744_ (_03273_, _03272_, _03268_);
  and _54745_ (_03274_, _03273_, _03252_);
  or _54746_ (_03275_, _03274_, _03251_);
  nand _54747_ (_03276_, _03275_, _03198_);
  nand _54748_ (_03277_, _03276_, _03227_);
  nor _54749_ (_03278_, _02873_, _02860_);
  nor _54750_ (_03279_, _03153_, \oc8051_golden_model_1.PC [3]);
  nor _54751_ (_03280_, _03279_, _03278_);
  or _54752_ (_03281_, _03280_, _03226_);
  nor _54753_ (_03282_, _03265_, _03261_);
  and _54754_ (_03283_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _54755_ (_03284_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _54756_ (_03285_, _03284_, _03283_);
  not _54757_ (_03286_, _03285_);
  nor _54758_ (_03287_, _03286_, _03282_);
  and _54759_ (_03288_, _03286_, _03282_);
  nor _54760_ (_03289_, _03288_, _03287_);
  or _54761_ (_03290_, _03289_, _03254_);
  not _54762_ (_03291_, _02867_);
  nor _54763_ (_03292_, _03241_, _02856_);
  nor _54764_ (_03293_, _03292_, _03291_);
  and _54765_ (_03294_, _03254_, _03293_);
  nand _54766_ (_03295_, _03294_, _03216_);
  nand _54767_ (_03296_, _03295_, _03290_);
  and _54768_ (_03297_, _03296_, _03252_);
  nor _54769_ (_03298_, _03249_, _03244_);
  nor _54770_ (_03299_, _03293_, \oc8051_golden_model_1.ACC [3]);
  and _54771_ (_03300_, _03293_, \oc8051_golden_model_1.ACC [3]);
  nor _54772_ (_03301_, _03300_, _03299_);
  and _54773_ (_03302_, _03301_, _03298_);
  nor _54774_ (_03303_, _03301_, _03298_);
  nor _54775_ (_03304_, _03303_, _03302_);
  nor _54776_ (_03305_, _03304_, _03232_);
  or _54777_ (_03306_, _03305_, _03297_);
  nand _54778_ (_03307_, _03306_, _03198_);
  nand _54779_ (_03308_, _03307_, _03281_);
  or _54780_ (_03309_, _03308_, _03277_);
  or _54781_ (_03310_, _03225_, _02887_);
  not _54782_ (_03311_, _03254_);
  nor _54783_ (_03312_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _54784_ (_03313_, _03312_, _03256_);
  nand _54785_ (_03314_, _03313_, _03311_);
  and _54786_ (_03315_, _03254_, _02887_);
  nand _54787_ (_03316_, _03315_, _03216_);
  nand _54788_ (_03317_, _03316_, _03314_);
  nand _54789_ (_03318_, _03317_, _03224_);
  nand _54790_ (_03319_, _03318_, _03310_);
  nand _54791_ (_03320_, _03319_, _03232_);
  not _54792_ (_03321_, \oc8051_golden_model_1.ACC [0]);
  and _54793_ (_03322_, _03321_, \oc8051_golden_model_1.PC [0]);
  nor _54794_ (_03323_, _03322_, _03236_);
  and _54795_ (_03324_, _03323_, _03231_);
  not _54796_ (_03325_, _03324_);
  and _54797_ (_03326_, _03325_, _03198_);
  nand _54798_ (_03327_, _03326_, _03320_);
  or _54799_ (_03328_, _03198_, \oc8051_golden_model_1.PC [0]);
  nand _54800_ (_03329_, _03328_, _03327_);
  or _54801_ (_03330_, _03226_, _02860_);
  nor _54802_ (_03331_, _03258_, _03256_);
  nor _54803_ (_03332_, _03331_, _03259_);
  or _54804_ (_03333_, _03332_, _03254_);
  and _54805_ (_03334_, _03254_, _03234_);
  nand _54806_ (_03335_, _03334_, _03216_);
  nand _54807_ (_03336_, _03335_, _03333_);
  and _54808_ (_03337_, _03336_, _03252_);
  nor _54809_ (_03338_, _03238_, _03236_);
  nor _54810_ (_03339_, _03338_, _03239_);
  nor _54811_ (_03340_, _03339_, _03232_);
  or _54812_ (_03341_, _03340_, _03337_);
  nand _54813_ (_03342_, _03341_, _03198_);
  nand _54814_ (_03343_, _03342_, _03330_);
  or _54815_ (_03344_, _03343_, _03329_);
  or _54816_ (_03345_, _03344_, _03309_);
  or _54817_ (_03346_, _03345_, _42240_);
  and _54818_ (_03347_, _03342_, _03330_);
  or _54819_ (_03348_, _03347_, _03329_);
  and _54820_ (_03349_, _03276_, _03227_);
  or _54821_ (_03350_, _03308_, _03349_);
  or _54822_ (_03351_, _03350_, _03348_);
  or _54823_ (_03352_, _03351_, _41994_);
  and _54824_ (_03353_, _03352_, _03346_);
  and _54825_ (_03354_, _03307_, _03281_);
  or _54826_ (_03355_, _03354_, _03277_);
  or _54827_ (_03356_, _03355_, _03348_);
  or _54828_ (_03357_, _03356_, _41830_);
  or _54829_ (_03358_, _03354_, _03349_);
  or _54830_ (_03359_, _03358_, _03344_);
  or _54831_ (_03360_, _03359_, _41740_);
  and _54832_ (_03361_, _03360_, _03357_);
  and _54833_ (_03362_, _03361_, _03353_);
  and _54834_ (_03363_, _03328_, _03327_);
  or _54835_ (_03364_, _03343_, _03363_);
  or _54836_ (_03365_, _03364_, _03309_);
  or _54837_ (_03366_, _03365_, _42199_);
  or _54838_ (_03367_, _03348_, _03309_);
  or _54839_ (_03368_, _03367_, _42158_);
  and _54840_ (_03369_, _03368_, _03366_);
  or _54841_ (_03370_, _03355_, _03344_);
  or _54842_ (_03371_, _03370_, _41912_);
  or _54843_ (_03372_, _03347_, _03363_);
  or _54844_ (_03373_, _03355_, _03372_);
  or _54845_ (_03374_, _03373_, _41789_);
  and _54846_ (_03375_, _03374_, _03371_);
  and _54847_ (_03376_, _03375_, _03369_);
  and _54848_ (_03377_, _03376_, _03362_);
  or _54849_ (_03378_, _03350_, _03364_);
  or _54850_ (_03379_, _03378_, _42035_);
  or _54851_ (_03380_, _03350_, _03372_);
  or _54852_ (_03381_, _03380_, _41953_);
  and _54853_ (_03382_, _03381_, _03379_);
  or _54854_ (_03383_, _03358_, _03372_);
  or _54855_ (_03384_, _03383_, _41610_);
  or _54856_ (_03385_, _03358_, _03348_);
  or _54857_ (_03386_, _03385_, _41651_);
  and _54858_ (_03387_, _03386_, _03384_);
  and _54859_ (_03388_, _03387_, _03382_);
  or _54860_ (_03389_, _03372_, _03309_);
  or _54861_ (_03390_, _03389_, _42117_);
  or _54862_ (_03391_, _03355_, _03364_);
  or _54863_ (_03392_, _03391_, _41871_);
  and _54864_ (_03393_, _03392_, _03390_);
  or _54865_ (_03394_, _03350_, _03344_);
  or _54866_ (_03395_, _03394_, _42076_);
  or _54867_ (_03396_, _03358_, _03364_);
  or _54868_ (_03397_, _03396_, _41692_);
  and _54869_ (_03398_, _03397_, _03395_);
  and _54870_ (_03399_, _03398_, _03393_);
  and _54871_ (_03400_, _03399_, _03388_);
  nand _54872_ (_03401_, _03400_, _03377_);
  or _54873_ (_03402_, _03367_, _42178_);
  or _54874_ (_03403_, _03370_, _41932_);
  and _54875_ (_03404_, _03403_, _03402_);
  or _54876_ (_03405_, _03356_, _41850_);
  or _54877_ (_03406_, _03383_, _41630_);
  and _54878_ (_03407_, _03406_, _03405_);
  and _54879_ (_03408_, _03407_, _03404_);
  or _54880_ (_03409_, _03394_, _42096_);
  or _54881_ (_03410_, _03359_, _41768_);
  and _54882_ (_03411_, _03410_, _03409_);
  or _54883_ (_03412_, _03378_, _42055_);
  or _54884_ (_03413_, _03380_, _41973_);
  and _54885_ (_03414_, _03413_, _03412_);
  and _54886_ (_03415_, _03414_, _03411_);
  and _54887_ (_03416_, _03415_, _03408_);
  or _54888_ (_03417_, _03391_, _41891_);
  or _54889_ (_03418_, _03373_, _41809_);
  and _54890_ (_03419_, _03418_, _03417_);
  or _54891_ (_03420_, _03345_, _42260_);
  or _54892_ (_03421_, _03385_, _41671_);
  and _54893_ (_03422_, _03421_, _03420_);
  and _54894_ (_03423_, _03422_, _03419_);
  or _54895_ (_03424_, _03365_, _42219_);
  or _54896_ (_03425_, _03396_, _41719_);
  and _54897_ (_03426_, _03425_, _03424_);
  or _54898_ (_03427_, _03389_, _42137_);
  or _54899_ (_03428_, _03351_, _42014_);
  and _54900_ (_03429_, _03428_, _03427_);
  and _54901_ (_03430_, _03429_, _03426_);
  and _54902_ (_03431_, _03430_, _03423_);
  and _54903_ (_03432_, _03431_, _03416_);
  or _54904_ (_03433_, _03432_, _03401_);
  nor _54905_ (_03434_, _03433_, _03152_);
  nor _54906_ (_03435_, _03401_, _03152_);
  not _54907_ (_03436_, _03435_);
  and _54908_ (_03437_, _03220_, _03188_);
  not _54909_ (_03438_, _03437_);
  nor _54910_ (_03439_, _03438_, _03401_);
  or _54911_ (_03440_, _03391_, _41876_);
  or _54912_ (_03441_, _03356_, _41835_);
  and _54913_ (_03442_, _03441_, _03440_);
  or _54914_ (_03443_, _03359_, _41749_);
  or _54915_ (_03444_, _03396_, _41697_);
  and _54916_ (_03445_, _03444_, _03443_);
  and _54917_ (_03446_, _03445_, _03442_);
  or _54918_ (_03447_, _03367_, _42163_);
  or _54919_ (_03448_, _03380_, _41958_);
  and _54920_ (_03449_, _03448_, _03447_);
  or _54921_ (_03450_, _03394_, _42081_);
  or _54922_ (_03451_, _03351_, _41999_);
  and _54923_ (_03452_, _03451_, _03450_);
  and _54924_ (_03453_, _03452_, _03449_);
  and _54925_ (_03454_, _03453_, _03446_);
  or _54926_ (_03455_, _03383_, _41615_);
  or _54927_ (_03456_, _03385_, _41656_);
  and _54928_ (_03457_, _03456_, _03455_);
  or _54929_ (_03458_, _03370_, _41917_);
  or _54930_ (_03459_, _03373_, _41794_);
  and _54931_ (_03460_, _03459_, _03458_);
  and _54932_ (_03461_, _03460_, _03457_);
  or _54933_ (_03462_, _03345_, _42245_);
  or _54934_ (_03463_, _03365_, _42204_);
  and _54935_ (_03464_, _03463_, _03462_);
  or _54936_ (_03465_, _03389_, _42122_);
  or _54937_ (_03466_, _03378_, _42040_);
  and _54938_ (_03467_, _03466_, _03465_);
  and _54939_ (_03468_, _03467_, _03464_);
  and _54940_ (_03469_, _03468_, _03461_);
  and _54941_ (_03471_, _03469_, _03454_);
  not _54942_ (_03472_, _03471_);
  and _54943_ (_03473_, _03472_, _03439_);
  not _54944_ (_03474_, _03221_);
  nor _54945_ (_03475_, _03218_, _03113_);
  and _54946_ (_03476_, _03475_, _03078_);
  and _54947_ (_03477_, _03476_, _03186_);
  and _54948_ (_03478_, _03219_, _03077_);
  and _54949_ (_03479_, _03478_, _03186_);
  nor _54950_ (_03480_, _03479_, _03477_);
  and _54951_ (_03481_, _03147_, _03113_);
  and _54952_ (_03482_, _03481_, _03077_);
  and _54953_ (_03483_, _03481_, _03217_);
  or _54954_ (_03484_, _03483_, _03482_);
  and _54955_ (_03485_, _03484_, _03186_);
  not _54956_ (_03486_, _03485_);
  and _54957_ (_03487_, _03481_, _03079_);
  and _54958_ (_03488_, _03487_, _03186_);
  and _54959_ (_03489_, _03475_, _03077_);
  and _54960_ (_03490_, _03489_, _03186_);
  nor _54961_ (_03491_, _03490_, _03488_);
  and _54962_ (_03492_, _03491_, _03486_);
  and _54963_ (_03493_, _03492_, _03480_);
  and _54964_ (_03494_, _03493_, _03474_);
  nor _54965_ (_03495_, _03494_, _03401_);
  and _54966_ (_03496_, _03495_, _03471_);
  and _54967_ (_03497_, _03077_, _03043_);
  and _54968_ (_03498_, _03497_, _03149_);
  and _54969_ (_03499_, _03498_, _03222_);
  not _54970_ (_03500_, _03499_);
  nor _54971_ (_03501_, _03500_, _03433_);
  not _54972_ (_03502_, \oc8051_golden_model_1.SP [0]);
  nor _54973_ (_03503_, _03200_, _03502_);
  not _54974_ (_03504_, _03199_);
  and _54975_ (_03505_, _03498_, _03504_);
  not _54976_ (_03506_, _03505_);
  nor _54977_ (_03507_, _03506_, _03433_);
  nor _54978_ (_03508_, _03506_, _03401_);
  not _54979_ (_03509_, _03508_);
  not _54980_ (_03510_, _03205_);
  and _54981_ (_03511_, _03510_, _03150_);
  and _54982_ (_03512_, _03498_, _03510_);
  not _54983_ (_03513_, _03512_);
  nor _54984_ (_03514_, _03513_, _03433_);
  not _54985_ (_03515_, _03202_);
  and _54986_ (_03516_, _03498_, _03515_);
  not _54987_ (_03517_, _03516_);
  or _54988_ (_03518_, _03517_, _03433_);
  not _54989_ (_03519_, _03211_);
  and _54990_ (_03520_, _03220_, _03165_);
  not _54991_ (_03521_, _03520_);
  and _54992_ (_03522_, _03498_, _03171_);
  not _54993_ (_03523_, _03522_);
  and _54994_ (_03524_, _03220_, _03171_);
  and _54995_ (_03525_, _03524_, _03432_);
  not _54996_ (_03526_, _03524_);
  and _54997_ (_03527_, _03220_, _03504_);
  nor _54998_ (_03528_, _03527_, _03511_);
  not _54999_ (_03529_, _03528_);
  and _55000_ (_03530_, _03529_, _03432_);
  nor _55001_ (_03531_, _03345_, _42275_);
  nor _55002_ (_03532_, _03365_, _42234_);
  nor _55003_ (_03533_, _03532_, _03531_);
  nor _55004_ (_03534_, _03367_, _42193_);
  nor _55005_ (_03535_, _03394_, _42111_);
  nor _55006_ (_03536_, _03535_, _03534_);
  and _55007_ (_03537_, _03536_, _03533_);
  nor _55008_ (_03538_, _03370_, _41947_);
  nor _55009_ (_03539_, _03391_, _41906_);
  nor _55010_ (_03540_, _03539_, _03538_);
  nor _55011_ (_03541_, _03356_, _41865_);
  nor _55012_ (_03542_, _03396_, _41734_);
  nor _55013_ (_03543_, _03542_, _03541_);
  and _55014_ (_03544_, _03543_, _03540_);
  and _55015_ (_03545_, _03544_, _03537_);
  nor _55016_ (_03546_, _03380_, _41988_);
  nor _55017_ (_03547_, _03385_, _41686_);
  nor _55018_ (_03548_, _03547_, _03546_);
  nor _55019_ (_03549_, _03351_, _42029_);
  nor _55020_ (_03550_, _03359_, _41783_);
  nor _55021_ (_03551_, _03550_, _03549_);
  and _55022_ (_03552_, _03551_, _03548_);
  nor _55023_ (_03553_, _03389_, _42152_);
  nor _55024_ (_03554_, _03383_, _41645_);
  nor _55025_ (_03555_, _03554_, _03553_);
  nor _55026_ (_03556_, _03378_, _42070_);
  nor _55027_ (_03557_, _03373_, _41824_);
  nor _55028_ (_03558_, _03557_, _03556_);
  and _55029_ (_03559_, _03558_, _03555_);
  and _55030_ (_03560_, _03559_, _03552_);
  and _55031_ (_03561_, _03560_, _03545_);
  nor _55032_ (_03562_, _03561_, _03401_);
  not _55033_ (_03563_, _03432_);
  and _55034_ (_03564_, _03563_, _03401_);
  nor _55035_ (_03565_, _03564_, _03562_);
  and _55036_ (_03566_, _03565_, _03516_);
  not _55037_ (_03567_, \oc8051_golden_model_1.SP [3]);
  and _55038_ (_03568_, _03515_, _03150_);
  and _55039_ (_03569_, _03568_, _03567_);
  and _55040_ (_03570_, _03220_, _03515_);
  not _55041_ (_03571_, _03207_);
  and _55042_ (_03572_, _03220_, _03571_);
  nor _55043_ (_03573_, _03572_, _03570_);
  or _55044_ (_03574_, _03573_, _03432_);
  and _55045_ (_03575_, _03220_, _03510_);
  nor _55046_ (_03576_, _03568_, _03516_);
  nand _55047_ (_03577_, _03573_, \oc8051_golden_model_1.PSW [3]);
  and _55048_ (_03578_, _03577_, _03576_);
  or _55049_ (_03579_, _03578_, _03575_);
  and _55050_ (_03580_, _03579_, _03574_);
  or _55051_ (_03581_, _03580_, _03569_);
  nor _55052_ (_03582_, _03581_, _03566_);
  not _55053_ (_03583_, _03575_);
  nor _55054_ (_03584_, _03583_, _03432_);
  nor _55055_ (_03585_, _03584_, _03582_);
  nor _55056_ (_03586_, _03585_, _03512_);
  nor _55057_ (_03587_, _03565_, _03513_);
  nor _55058_ (_03588_, _03587_, _03529_);
  not _55059_ (_03589_, _03588_);
  nor _55060_ (_03590_, _03589_, _03586_);
  nor _55061_ (_03591_, _03590_, _03530_);
  and _55062_ (_03592_, _03504_, _03150_);
  nor _55063_ (_03593_, _03592_, _03505_);
  not _55064_ (_03594_, _03593_);
  or _55065_ (_03595_, _03594_, _03591_);
  not _55066_ (_03596_, _03212_);
  and _55067_ (_03597_, _03484_, _03596_);
  not _55068_ (_03598_, _03597_);
  and _55069_ (_03599_, _03487_, _03596_);
  and _55070_ (_03600_, _03475_, _03596_);
  nor _55071_ (_03601_, _03600_, _03599_);
  and _55072_ (_03602_, _03601_, _03598_);
  nand _55073_ (_03603_, _03594_, _03565_);
  and _55074_ (_03604_, _03603_, _03602_);
  and _55075_ (_03605_, _03604_, _03595_);
  and _55076_ (_03606_, _03596_, _03150_);
  and _55077_ (_03607_, _03498_, _03596_);
  nor _55078_ (_03608_, _03607_, _03606_);
  not _55079_ (_03609_, _03608_);
  nor _55080_ (_03610_, _03602_, _03432_);
  nor _55081_ (_03611_, _03610_, _03609_);
  not _55082_ (_03612_, _03611_);
  nor _55083_ (_03613_, _03612_, _03605_);
  and _55084_ (_03614_, _03222_, _03220_);
  and _55085_ (_03615_, _03609_, _03565_);
  nor _55086_ (_03616_, _03615_, _03614_);
  not _55087_ (_03617_, _03616_);
  or _55088_ (_03618_, _03617_, _03613_);
  not _55089_ (_03619_, _03614_);
  nor _55090_ (_03620_, _03619_, _03432_);
  nor _55091_ (_03621_, _03620_, _03499_);
  nand _55092_ (_03622_, _03621_, _03618_);
  and _55093_ (_03623_, _03565_, _03499_);
  nor _55094_ (_03624_, _03623_, _03221_);
  nand _55095_ (_03625_, _03624_, _03622_);
  not _55096_ (_03626_, _03155_);
  and _55097_ (_03627_, _03177_, _03150_);
  and _55098_ (_03628_, _03171_, _03150_);
  nor _55099_ (_03629_, _03628_, _03627_);
  and _55100_ (_03630_, _03629_, _03152_);
  and _55101_ (_03631_, _03630_, _03438_);
  and _55102_ (_03632_, _03222_, _03150_);
  and _55103_ (_03633_, _03481_, _03497_);
  and _55104_ (_03634_, _03633_, _03504_);
  nor _55105_ (_03635_, _03634_, _03632_);
  and _55106_ (_03636_, _03230_, _03193_);
  and _55107_ (_03637_, _03219_, _03079_);
  and _55108_ (_03638_, _03637_, _03504_);
  nor _55109_ (_03639_, _03638_, _03636_);
  and _55110_ (_03640_, _03639_, _03635_);
  and _55111_ (_03641_, _03498_, _03010_);
  nor _55112_ (_03642_, _03641_, _03527_);
  and _55113_ (_03643_, _03181_, _03168_);
  and _55114_ (_03644_, _03230_, _03643_);
  and _55115_ (_03645_, _03498_, _03165_);
  nor _55116_ (_03646_, _03645_, _03644_);
  and _55117_ (_03647_, _03646_, _03642_);
  and _55118_ (_03648_, _03647_, _03640_);
  and _55119_ (_03649_, _03648_, _03631_);
  and _55120_ (_03650_, _03475_, _03079_);
  or _55121_ (_03651_, _03650_, _03483_);
  and _55122_ (_03652_, _03651_, _03504_);
  not _55123_ (_03653_, _03652_);
  not _55124_ (_03654_, _03228_);
  and _55125_ (_03655_, _03481_, _03654_);
  and _55126_ (_03656_, _03655_, _03504_);
  and _55127_ (_03657_, _03478_, _03504_);
  or _55128_ (_03658_, _03657_, _03570_);
  nor _55129_ (_03659_, _03658_, _03656_);
  and _55130_ (_03660_, _03659_, _03653_);
  and _55131_ (_03661_, _03475_, _03654_);
  nor _55132_ (_03662_, _03661_, _03487_);
  and _55133_ (_03663_, _03475_, _03497_);
  and _55134_ (_03664_, _03475_, _03217_);
  nor _55135_ (_03665_, _03664_, _03663_);
  and _55136_ (_03666_, _03665_, _03662_);
  nor _55137_ (_03667_, _03666_, _03199_);
  not _55138_ (_03668_, _03667_);
  and _55139_ (_03669_, _03668_, _03660_);
  and _55140_ (_03670_, _03669_, _03649_);
  nor _55141_ (_03672_, _03670_, _03626_);
  and _55142_ (_03673_, _03670_, _03243_);
  nor _55143_ (_03674_, _03673_, _03672_);
  not _55144_ (_03675_, _03280_);
  nor _55145_ (_03676_, _03670_, _03675_);
  not _55146_ (_03677_, _03293_);
  and _55147_ (_03678_, _03670_, _03677_);
  nor _55148_ (_03679_, _03678_, _03676_);
  nor _55149_ (_03680_, _03679_, _03674_);
  nor _55150_ (_03681_, _03670_, _02887_);
  and _55151_ (_03682_, _03670_, _02887_);
  nor _55152_ (_03683_, _03682_, _03681_);
  not _55153_ (_03684_, _03683_);
  nor _55154_ (_03685_, _03682_, _02860_);
  and _55155_ (_03686_, _03682_, _02860_);
  nor _55156_ (_03687_, _03686_, _03685_);
  and _55157_ (_03688_, _03687_, _03684_);
  and _55158_ (_03689_, _03688_, _03680_);
  and _55159_ (_03690_, _03689_, _02000_);
  nor _55160_ (_03691_, _03687_, _03683_);
  and _55161_ (_03692_, _03679_, _03674_);
  and _55162_ (_03693_, _03692_, _03691_);
  and _55163_ (_03694_, _03693_, _02013_);
  nor _55164_ (_03695_, _03694_, _03690_);
  not _55165_ (_03696_, _03674_);
  nor _55166_ (_03697_, _03679_, _03696_);
  and _55167_ (_03698_, _03697_, _03688_);
  and _55168_ (_03699_, _03698_, _02032_);
  and _55169_ (_03700_, _03692_, _03688_);
  and _55170_ (_03701_, _03700_, _02024_);
  nor _55171_ (_03702_, _03701_, _03699_);
  and _55172_ (_03703_, _03702_, _03695_);
  and _55173_ (_03704_, _03697_, _03691_);
  and _55174_ (_03705_, _03704_, _02017_);
  and _55175_ (_03706_, _03687_, _03683_);
  and _55176_ (_03707_, _03692_, _03706_);
  and _55177_ (_03708_, _03707_, _02026_);
  nor _55178_ (_03709_, _03708_, _03705_);
  and _55179_ (_03710_, _03679_, _03696_);
  and _55180_ (_03711_, _03710_, _03688_);
  and _55181_ (_03712_, _03711_, _01997_);
  and _55182_ (_03713_, _03710_, _03691_);
  and _55183_ (_03714_, _03713_, _02010_);
  nor _55184_ (_03715_, _03714_, _03712_);
  and _55185_ (_03716_, _03715_, _03709_);
  and _55186_ (_03717_, _03716_, _03703_);
  nor _55187_ (_03718_, _03687_, _03684_);
  and _55188_ (_03719_, _03710_, _03718_);
  and _55189_ (_03720_, _03719_, _02008_);
  and _55190_ (_03721_, _03692_, _03718_);
  and _55191_ (_03722_, _03721_, _02002_);
  nor _55192_ (_03723_, _03722_, _03720_);
  and _55193_ (_03724_, _03706_, _03680_);
  and _55194_ (_03725_, _03724_, _02043_);
  and _55195_ (_03726_, _03697_, _03706_);
  and _55196_ (_03727_, _03726_, _02034_);
  nor _55197_ (_03728_, _03727_, _03725_);
  and _55198_ (_03729_, _03728_, _03723_);
  and _55199_ (_03730_, _03691_, _03680_);
  and _55200_ (_03731_, _03730_, _02019_);
  and _55201_ (_03732_, _03718_, _03697_);
  and _55202_ (_03733_, _03732_, _02030_);
  nor _55203_ (_03734_, _03733_, _03731_);
  and _55204_ (_03735_, _03718_, _03680_);
  and _55205_ (_03736_, _03735_, _02036_);
  and _55206_ (_03737_, _03710_, _03706_);
  and _55207_ (_03738_, _03737_, _02046_);
  nor _55208_ (_03739_, _03738_, _03736_);
  and _55209_ (_03740_, _03739_, _03734_);
  and _55210_ (_03741_, _03740_, _03729_);
  and _55211_ (_03742_, _03741_, _03717_);
  nor _55212_ (_03743_, _03742_, _03474_);
  and _55213_ (_03744_, _03498_, _03188_);
  and _55214_ (_03745_, _03498_, _03186_);
  nor _55215_ (_03746_, _03745_, _03744_);
  not _55216_ (_03747_, _03746_);
  nor _55217_ (_03748_, _03747_, _03743_);
  and _55218_ (_03749_, _03748_, _03625_);
  and _55219_ (_03750_, _03747_, _03565_);
  or _55220_ (_03751_, _03750_, _03749_);
  and _55221_ (_03752_, _03498_, _03191_);
  not _55222_ (_03753_, _03752_);
  and _55223_ (_03754_, _03230_, _03191_);
  and _55224_ (_03755_, _03220_, _03191_);
  nor _55225_ (_03756_, _03755_, _03754_);
  and _55226_ (_03757_, _03756_, _03753_);
  and _55227_ (_03758_, _03230_, _03182_);
  not _55228_ (_03759_, _03758_);
  and _55229_ (_03760_, _03498_, _03182_);
  and _55230_ (_03761_, _03220_, _03182_);
  nor _55231_ (_03762_, _03761_, _03760_);
  and _55232_ (_03763_, _03762_, _03759_);
  and _55233_ (_03764_, _03763_, _03757_);
  and _55234_ (_03765_, _03220_, _03177_);
  not _55235_ (_03766_, _03765_);
  and _55236_ (_03767_, _03220_, _03193_);
  not _55237_ (_03768_, _03767_);
  and _55238_ (_03769_, _03498_, _03193_);
  nor _55239_ (_03770_, _03769_, _03636_);
  and _55240_ (_03771_, _03770_, _03768_);
  and _55241_ (_03772_, _03771_, _03766_);
  and _55242_ (_03773_, _03772_, _03764_);
  nand _55243_ (_03774_, _03773_, _03751_);
  and _55244_ (_03775_, _03498_, _03177_);
  nor _55245_ (_03776_, _03773_, _03563_);
  nor _55246_ (_03777_, _03776_, _03775_);
  and _55247_ (_03778_, _03777_, _03774_);
  and _55248_ (_03779_, _03775_, \oc8051_golden_model_1.SP [3]);
  or _55249_ (_03780_, _03779_, _03627_);
  nor _55250_ (_03781_, _03780_, _03778_);
  and _55251_ (_03782_, _03565_, _03627_);
  or _55252_ (_03783_, _03782_, _03781_);
  and _55253_ (_03784_, _03783_, _03526_);
  or _55254_ (_03785_, _03784_, _03525_);
  nand _55255_ (_03786_, _03785_, _03523_);
  and _55256_ (_03787_, _03522_, _03567_);
  nor _55257_ (_03788_, _03787_, _03628_);
  nand _55258_ (_03789_, _03788_, _03786_);
  and _55259_ (_03790_, _03220_, _03010_);
  not _55260_ (_03791_, _03628_);
  nor _55261_ (_03792_, _03791_, _03565_);
  nor _55262_ (_03793_, _03792_, _03790_);
  nand _55263_ (_03794_, _03793_, _03789_);
  and _55264_ (_03795_, _03790_, _03432_);
  nor _55265_ (_03796_, _03795_, _03151_);
  and _55266_ (_03797_, _03796_, _03794_);
  nor _55267_ (_03798_, _03565_, _03152_);
  or _55268_ (_03799_, _03798_, _03797_);
  nand _55269_ (_03800_, _03799_, _03521_);
  nor _55270_ (_03801_, _03521_, _03432_);
  not _55271_ (_03802_, _03801_);
  and _55272_ (_03803_, _03802_, _03800_);
  nor _55273_ (_03804_, _03383_, _41640_);
  nor _55274_ (_03805_, _03396_, _41729_);
  nor _55275_ (_03806_, _03805_, _03804_);
  nor _55276_ (_03807_, _03365_, _42229_);
  nor _55277_ (_03808_, _03391_, _41901_);
  nor _55278_ (_03809_, _03808_, _03807_);
  and _55279_ (_03810_, _03809_, _03806_);
  nor _55280_ (_03811_, _03394_, _42106_);
  nor _55281_ (_03812_, _03380_, _41983_);
  nor _55282_ (_03813_, _03812_, _03811_);
  nor _55283_ (_03814_, _03373_, _41819_);
  nor _55284_ (_03815_, _03385_, _41681_);
  nor _55285_ (_03816_, _03815_, _03814_);
  and _55286_ (_03817_, _03816_, _03813_);
  and _55287_ (_03818_, _03817_, _03810_);
  nor _55288_ (_03819_, _03389_, _42147_);
  nor _55289_ (_03820_, _03351_, _42024_);
  nor _55290_ (_03821_, _03820_, _03819_);
  nor _55291_ (_03822_, _03345_, _42270_);
  nor _55292_ (_03823_, _03367_, _42188_);
  nor _55293_ (_03824_, _03823_, _03822_);
  and _55294_ (_03825_, _03824_, _03821_);
  nor _55295_ (_03826_, _03378_, _42065_);
  nor _55296_ (_03827_, _03359_, _41778_);
  nor _55297_ (_03828_, _03827_, _03826_);
  nor _55298_ (_03829_, _03370_, _41942_);
  nor _55299_ (_03830_, _03356_, _41860_);
  nor _55300_ (_03831_, _03830_, _03829_);
  and _55301_ (_03832_, _03831_, _03828_);
  and _55302_ (_03833_, _03832_, _03825_);
  and _55303_ (_03834_, _03833_, _03818_);
  nor _55304_ (_03835_, _03834_, _03401_);
  and _55305_ (_03836_, _03835_, _03499_);
  not _55306_ (_03837_, _03836_);
  not _55307_ (_03838_, _03835_);
  and _55308_ (_03839_, _03608_, _03513_);
  and _55309_ (_03840_, _03839_, _03593_);
  and _55310_ (_03841_, _03746_, _03517_);
  and _55311_ (_03842_, _03841_, _03630_);
  and _55312_ (_03843_, _03842_, _03840_);
  nor _55313_ (_03844_, _03843_, _03838_);
  not _55314_ (_03845_, _03844_);
  nor _55315_ (_03846_, _03345_, _42255_);
  nor _55316_ (_03847_, _03359_, _41763_);
  nor _55317_ (_03848_, _03847_, _03846_);
  nor _55318_ (_03849_, _03365_, _42214_);
  nor _55319_ (_03850_, _03380_, _41968_);
  nor _55320_ (_03851_, _03850_, _03849_);
  and _55321_ (_03852_, _03851_, _03848_);
  nor _55322_ (_03853_, _03394_, _42091_);
  nor _55323_ (_03854_, _03370_, _41927_);
  nor _55324_ (_03855_, _03854_, _03853_);
  nor _55325_ (_03856_, _03391_, _41886_);
  nor _55326_ (_03857_, _03385_, _41666_);
  nor _55327_ (_03858_, _03857_, _03856_);
  and _55328_ (_03859_, _03858_, _03855_);
  and _55329_ (_03860_, _03859_, _03852_);
  nor _55330_ (_03861_, _03367_, _42173_);
  nor _55331_ (_03862_, _03389_, _42132_);
  nor _55332_ (_03863_, _03862_, _03861_);
  nor _55333_ (_03864_, _03351_, _42009_);
  nor _55334_ (_03865_, _03373_, _41804_);
  nor _55335_ (_03866_, _03865_, _03864_);
  and _55336_ (_03867_, _03866_, _03863_);
  nor _55337_ (_03868_, _03378_, _42050_);
  nor _55338_ (_03869_, _03396_, _41714_);
  nor _55339_ (_03870_, _03869_, _03868_);
  nor _55340_ (_03871_, _03356_, _41845_);
  nor _55341_ (_03873_, _03383_, _41625_);
  nor _55342_ (_03874_, _03873_, _03871_);
  and _55343_ (_03875_, _03874_, _03870_);
  and _55344_ (_03876_, _03875_, _03867_);
  and _55345_ (_03877_, _03876_, _03860_);
  nor _55346_ (_03878_, _03614_, _03575_);
  and _55347_ (_03879_, _03878_, _03528_);
  and _55348_ (_03880_, _03879_, _03573_);
  and _55349_ (_03881_, _03880_, _03602_);
  nor _55350_ (_03882_, _03790_, _03520_);
  nor _55351_ (_03883_, _03765_, _03524_);
  and _55352_ (_03884_, _03883_, _03882_);
  and _55353_ (_03885_, _03884_, _03771_);
  and _55354_ (_03886_, _03885_, _03764_);
  and _55355_ (_03887_, _03886_, _03881_);
  nor _55356_ (_03888_, _03887_, _03877_);
  not _55357_ (_03889_, _03888_);
  and _55358_ (_03890_, _03711_, _01983_);
  and _55359_ (_03891_, _03700_, _01962_);
  nor _55360_ (_03892_, _03891_, _03890_);
  and _55361_ (_03893_, _03724_, _01941_);
  and _55362_ (_03894_, _03735_, _01944_);
  nor _55363_ (_03895_, _03894_, _03893_);
  and _55364_ (_03896_, _03895_, _03892_);
  and _55365_ (_03897_, _03737_, _01971_);
  and _55366_ (_03898_, _03713_, _01966_);
  nor _55367_ (_03899_, _03898_, _03897_);
  and _55368_ (_03900_, _03707_, _01978_);
  and _55369_ (_03901_, _03693_, _01969_);
  nor _55370_ (_03902_, _03901_, _03900_);
  and _55371_ (_03903_, _03902_, _03899_);
  and _55372_ (_03904_, _03903_, _03896_);
  and _55373_ (_03905_, _03726_, _01989_);
  and _55374_ (_03906_, _03732_, _01954_);
  nor _55375_ (_03907_, _03906_, _03905_);
  and _55376_ (_03908_, _03689_, _01952_);
  and _55377_ (_03909_, _03730_, _01976_);
  nor _55378_ (_03910_, _03909_, _03908_);
  and _55379_ (_03911_, _03910_, _03907_);
  and _55380_ (_03912_, _03719_, _01960_);
  and _55381_ (_03913_, _03721_, _01980_);
  nor _55382_ (_03914_, _03913_, _03912_);
  and _55383_ (_03915_, _03698_, _01946_);
  and _55384_ (_03916_, _03704_, _01986_);
  nor _55385_ (_03917_, _03916_, _03915_);
  and _55386_ (_03918_, _03917_, _03914_);
  and _55387_ (_03919_, _03918_, _03911_);
  and _55388_ (_03920_, _03919_, _03904_);
  nor _55389_ (_03921_, _03920_, _03474_);
  and _55390_ (_03922_, _03482_, _03571_);
  and _55391_ (_03923_, _03483_, _03571_);
  or _55392_ (_03924_, _03923_, _03922_);
  and _55393_ (_03925_, _03481_, _03078_);
  and _55394_ (_03926_, _03925_, _03182_);
  nor _55395_ (_03927_, _03926_, _03924_);
  and _55396_ (_03928_, _03925_, _03191_);
  and _55397_ (_03929_, _03925_, _03504_);
  nor _55398_ (_03930_, _03929_, _03928_);
  and _55399_ (_03931_, _03930_, _03927_);
  and _55400_ (_03932_, _03487_, _03193_);
  not _55401_ (_03933_, _03932_);
  and _55402_ (_03934_, _03482_, _03193_);
  and _55403_ (_03935_, _03483_, _03193_);
  nor _55404_ (_03936_, _03935_, _03934_);
  and _55405_ (_03937_, _03936_, _03933_);
  and _55406_ (_03938_, _03482_, _03186_);
  and _55407_ (_03939_, _03925_, _03171_);
  nor _55408_ (_03940_, _03939_, _03938_);
  and _55409_ (_03941_, _03940_, _03937_);
  and _55410_ (_03942_, _03941_, _03931_);
  and _55411_ (_03943_, _03482_, _03510_);
  not _55412_ (_03944_, _03943_);
  and _55413_ (_03945_, _03482_, _03010_);
  and _55414_ (_03946_, _03482_, _03182_);
  nor _55415_ (_03947_, _03946_, _03945_);
  and _55416_ (_03948_, _03947_, _03944_);
  and _55417_ (_03949_, _03482_, _03165_);
  and _55418_ (_03950_, _03482_, _03191_);
  nor _55419_ (_03951_, _03950_, _03949_);
  and _55420_ (_03952_, _03482_, _03171_);
  and _55421_ (_03953_, _03482_, _03177_);
  nor _55422_ (_03954_, _03953_, _03952_);
  and _55423_ (_03955_, _03954_, _03951_);
  and _55424_ (_03956_, _03955_, _03948_);
  and _55425_ (_03957_, _03956_, _03942_);
  and _55426_ (_03958_, _03483_, _03177_);
  and _55427_ (_03959_, _03487_, _03571_);
  nor _55428_ (_03960_, _03959_, _03958_);
  and _55429_ (_03961_, _03482_, _03222_);
  and _55430_ (_03962_, _03482_, _03504_);
  or _55431_ (_03963_, _03962_, _03961_);
  nor _55432_ (_03964_, _03185_, _03007_);
  and _55433_ (_03965_, _03964_, _03483_);
  nor _55434_ (_03966_, _03965_, _03963_);
  and _55435_ (_03967_, _03966_, _03960_);
  not _55436_ (_03968_, _03488_);
  and _55437_ (_03969_, _03925_, _03165_);
  and _55438_ (_03970_, _03925_, _03010_);
  nor _55439_ (_03971_, _03970_, _03969_);
  and _55440_ (_03972_, _03971_, _03968_);
  and _55441_ (_03973_, _03487_, _03177_);
  and _55442_ (_03974_, _03487_, _03222_);
  nor _55443_ (_03975_, _03974_, _03973_);
  and _55444_ (_03976_, _03975_, _03972_);
  and _55445_ (_03977_, _03976_, _03967_);
  and _55446_ (_03978_, _03925_, _03510_);
  and _55447_ (_03979_, _03481_, _03515_);
  nor _55448_ (_03980_, _03979_, _03978_);
  not _55449_ (_03981_, _03980_);
  not _55450_ (_03982_, \oc8051_golden_model_1.SP [2]);
  not _55451_ (_03983_, _03568_);
  nor _55452_ (_03984_, _03775_, _03522_);
  and _55453_ (_03985_, _03984_, _03983_);
  nor _55454_ (_03986_, _03985_, _03982_);
  nor _55455_ (_03987_, _03986_, _03981_);
  and _55456_ (_03988_, _03987_, _03977_);
  and _55457_ (_03989_, _03988_, _03957_);
  not _55458_ (_03990_, _03989_);
  nor _55459_ (_03991_, _03990_, _03921_);
  and _55460_ (_03992_, _03991_, _03889_);
  and _55461_ (_03993_, _03992_, _03845_);
  and _55462_ (_03994_, _03993_, _03837_);
  nor _55463_ (_03995_, _03521_, _03471_);
  not _55464_ (_03996_, _03995_);
  nor _55465_ (_03997_, _03619_, _03471_);
  not _55466_ (_03998_, _03527_);
  nor _55467_ (_03999_, _03998_, _03471_);
  or _55468_ (_04000_, _03583_, _03471_);
  nor _55469_ (_04001_, _03573_, _03471_);
  not _55470_ (_04002_, _03663_);
  nor _55471_ (_04003_, _03487_, _03220_);
  and _55472_ (_04004_, _03497_, _03219_);
  nor _55473_ (_04005_, _04004_, _03650_);
  and _55474_ (_04006_, _04005_, _04003_);
  and _55475_ (_04007_, _04006_, _04002_);
  nor _55476_ (_04008_, _04007_, _03207_);
  not _55477_ (_04009_, _04008_);
  not _55478_ (_04010_, _03210_);
  and _55479_ (_04011_, _04004_, _04010_);
  and _55480_ (_04012_, _03633_, _03571_);
  nor _55481_ (_04013_, _04012_, _04011_);
  nor _55482_ (_04014_, _04003_, _03202_);
  not _55483_ (_04015_, _04014_);
  and _55484_ (_04016_, _04004_, _03515_);
  not _55485_ (_04017_, _04016_);
  and _55486_ (_04018_, _03633_, _03515_);
  and _55487_ (_04019_, _03475_, _03043_);
  and _55488_ (_04020_, _04019_, _03515_);
  nor _55489_ (_04021_, _04020_, _04018_);
  and _55490_ (_04022_, _04021_, _04017_);
  and _55491_ (_04023_, _04022_, _04015_);
  and _55492_ (_04024_, _04023_, _04013_);
  and _55493_ (_04025_, _04024_, _04009_);
  or _55494_ (_04026_, _04025_, _04001_);
  nand _55495_ (_04027_, _04026_, _03517_);
  nand _55496_ (_04028_, _03518_, _04027_);
  nor _55497_ (_04029_, _04006_, _03205_);
  not _55498_ (_04030_, _04029_);
  and _55499_ (_04031_, _03568_, _03502_);
  not _55500_ (_04032_, _03043_);
  and _55501_ (_04033_, _03489_, _03510_);
  nor _55502_ (_04034_, _04033_, _03943_);
  nor _55503_ (_04035_, _04034_, _04032_);
  nor _55504_ (_04036_, _04035_, _04031_);
  and _55505_ (_04037_, _04036_, _04030_);
  nand _55506_ (_04038_, _04037_, _04028_);
  nand _55507_ (_04039_, _04038_, _04000_);
  and _55508_ (_04040_, _04039_, _03513_);
  or _55509_ (_04041_, _03514_, _04040_);
  and _55510_ (_04042_, _03511_, _03471_);
  nor _55511_ (_04043_, _03663_, _03633_);
  and _55512_ (_04044_, _04043_, _04005_);
  and _55513_ (_04045_, _04044_, _04003_);
  nor _55514_ (_04046_, _04045_, _03199_);
  nor _55515_ (_04047_, _04046_, _04042_);
  and _55516_ (_04048_, _04047_, _04041_);
  or _55517_ (_04049_, _04048_, _03999_);
  and _55518_ (_04050_, _04049_, _03593_);
  nor _55519_ (_04051_, _03593_, _03433_);
  or _55520_ (_04052_, _04051_, _04050_);
  not _55521_ (_04053_, _03602_);
  and _55522_ (_04054_, _04053_, _03471_);
  and _55523_ (_04055_, _04004_, _03596_);
  nor _55524_ (_04056_, _04055_, _03609_);
  not _55525_ (_04057_, _04056_);
  nor _55526_ (_04058_, _04057_, _04054_);
  and _55527_ (_04059_, _04058_, _04052_);
  nor _55528_ (_04060_, _03608_, _03433_);
  nor _55529_ (_04061_, _04060_, _04059_);
  nor _55530_ (_04062_, _04045_, _03253_);
  nor _55531_ (_04063_, _04062_, _04061_);
  or _55532_ (_04064_, _04063_, _03997_);
  and _55533_ (_04065_, _04064_, _03500_);
  or _55534_ (_04066_, _04065_, _03501_);
  and _55535_ (_04067_, _03663_, _03186_);
  nor _55536_ (_04068_, _04067_, _03488_);
  and _55537_ (_04069_, _04004_, _03186_);
  and _55538_ (_04070_, _03650_, _03186_);
  not _55539_ (_04071_, _03186_);
  nor _55540_ (_04072_, _03633_, _03220_);
  nor _55541_ (_04074_, _04072_, _04071_);
  or _55542_ (_04075_, _04074_, _04070_);
  nor _55543_ (_04076_, _04075_, _04069_);
  and _55544_ (_04077_, _04076_, _04068_);
  and _55545_ (_04078_, _04077_, _04066_);
  and _55546_ (_04079_, _03732_, _01840_);
  and _55547_ (_04080_, _03719_, _01853_);
  nor _55548_ (_04081_, _04080_, _04079_);
  and _55549_ (_04082_, _03689_, _01842_);
  and _55550_ (_04083_, _03711_, _01873_);
  nor _55551_ (_04084_, _04083_, _04082_);
  and _55552_ (_04085_, _04084_, _04081_);
  and _55553_ (_04086_, _03704_, _01875_);
  and _55554_ (_04087_, _03713_, _01848_);
  nor _55555_ (_04088_, _04087_, _04086_);
  and _55556_ (_04089_, _03721_, _01868_);
  and _55557_ (_04090_, _03693_, _01858_);
  nor _55558_ (_04091_, _04090_, _04089_);
  and _55559_ (_04092_, _04091_, _04088_);
  and _55560_ (_04093_, _04092_, _04085_);
  and _55561_ (_04094_, _03730_, _01866_);
  and _55562_ (_04095_, _03698_, _01829_);
  nor _55563_ (_04096_, _04095_, _04094_);
  and _55564_ (_04097_, _03737_, _01861_);
  and _55565_ (_04098_, _03707_, _01870_);
  nor _55566_ (_04099_, _04098_, _04097_);
  and _55567_ (_04100_, _04099_, _04096_);
  and _55568_ (_04101_, _03735_, _01832_);
  and _55569_ (_04102_, _03726_, _01877_);
  nor _55570_ (_04103_, _04102_, _04101_);
  and _55571_ (_04104_, _03724_, _01836_);
  and _55572_ (_04105_, _03700_, _01850_);
  nor _55573_ (_04106_, _04105_, _04104_);
  and _55574_ (_04107_, _04106_, _04103_);
  and _55575_ (_04108_, _04107_, _04100_);
  and _55576_ (_04109_, _04108_, _04093_);
  nor _55577_ (_04110_, _04109_, _03474_);
  or _55578_ (_04111_, _04110_, _04078_);
  and _55579_ (_04112_, _03745_, _03433_);
  and _55580_ (_04113_, _04004_, _03188_);
  nor _55581_ (_04114_, _04113_, _03744_);
  not _55582_ (_04115_, _04114_);
  nor _55583_ (_04116_, _04115_, _04112_);
  and _55584_ (_04117_, _04116_, _04111_);
  not _55585_ (_04118_, _03744_);
  nor _55586_ (_04119_, _04118_, _03433_);
  or _55587_ (_04120_, _04119_, _04117_);
  not _55588_ (_04121_, _03193_);
  nor _55589_ (_04122_, _03663_, _03487_);
  nor _55590_ (_04123_, _04122_, _04121_);
  not _55591_ (_04124_, _04123_);
  and _55592_ (_04125_, _04004_, _03193_);
  not _55593_ (_04126_, _04125_);
  and _55594_ (_04127_, _03934_, _03043_);
  and _55595_ (_04128_, _03476_, _03193_);
  and _55596_ (_04129_, _04128_, _03043_);
  nor _55597_ (_04130_, _04129_, _04127_);
  and _55598_ (_04131_, _04130_, _04126_);
  and _55599_ (_04132_, _04131_, _04124_);
  and _55600_ (_04133_, _04132_, _04120_);
  nor _55601_ (_04134_, _03771_, _03472_);
  and _55602_ (_04135_, _03476_, _03191_);
  and _55603_ (_04136_, _04135_, _03043_);
  not _55604_ (_04137_, _04136_);
  and _55605_ (_04138_, _04004_, _03191_);
  not _55606_ (_04139_, _04138_);
  and _55607_ (_04140_, _03663_, _03191_);
  and _55608_ (_04141_, _03147_, _03043_);
  and _55609_ (_04142_, _04141_, _03113_);
  and _55610_ (_04143_, _04142_, _03191_);
  nor _55611_ (_04144_, _04143_, _04140_);
  and _55612_ (_04145_, _04144_, _04139_);
  and _55613_ (_04146_, _04145_, _04137_);
  not _55614_ (_04147_, _04146_);
  nor _55615_ (_04148_, _04147_, _04134_);
  and _55616_ (_04149_, _04148_, _04133_);
  nor _55617_ (_04150_, _03764_, _03472_);
  and _55618_ (_04151_, _03663_, _03177_);
  nor _55619_ (_04152_, _04151_, _03973_);
  and _55620_ (_04153_, _04004_, _03177_);
  not _55621_ (_04154_, _04153_);
  and _55622_ (_04155_, _03650_, _03177_);
  not _55623_ (_04156_, _03177_);
  nor _55624_ (_04157_, _04072_, _04156_);
  nor _55625_ (_04158_, _04157_, _04155_);
  and _55626_ (_04159_, _04158_, _04154_);
  and _55627_ (_04160_, _04159_, _04152_);
  and _55628_ (_04161_, _03650_, _03182_);
  and _55629_ (_04162_, _04142_, _03182_);
  nor _55630_ (_04163_, _04162_, _04161_);
  and _55631_ (_04164_, _03663_, _03182_);
  and _55632_ (_04165_, _04004_, _03182_);
  nor _55633_ (_04166_, _04165_, _04164_);
  and _55634_ (_04167_, _04166_, _04163_);
  and _55635_ (_04168_, _04167_, _04160_);
  not _55636_ (_04169_, _04168_);
  nor _55637_ (_04170_, _04169_, _04150_);
  and _55638_ (_04171_, _04170_, _04149_);
  nor _55639_ (_04172_, _03766_, _03471_);
  nor _55640_ (_04173_, _04172_, _04171_);
  and _55641_ (_04175_, _03775_, _03502_);
  nor _55642_ (_04176_, _04175_, _04173_);
  and _55643_ (_04177_, _03627_, _03433_);
  not _55644_ (_04178_, _03171_);
  nor _55645_ (_04179_, _04045_, _04178_);
  nor _55646_ (_04180_, _04179_, _04177_);
  and _55647_ (_04181_, _04180_, _04176_);
  nor _55648_ (_04182_, _03526_, _03471_);
  nor _55649_ (_04183_, _04182_, _04181_);
  and _55650_ (_04184_, _03522_, _03502_);
  nor _55651_ (_04185_, _04184_, _04183_);
  and _55652_ (_04186_, _03628_, _03433_);
  and _55653_ (_04187_, _03487_, _03010_);
  and _55654_ (_04188_, _03663_, _03010_);
  or _55655_ (_04189_, _04188_, _04187_);
  and _55656_ (_04190_, _04004_, _03010_);
  nor _55657_ (_04191_, _04190_, _04189_);
  not _55658_ (_04192_, _03790_);
  and _55659_ (_04193_, _03633_, _03010_);
  and _55660_ (_04194_, _03650_, _03010_);
  nor _55661_ (_04195_, _04194_, _04193_);
  and _55662_ (_04196_, _04195_, _04192_);
  and _55663_ (_04197_, _04196_, _04191_);
  not _55664_ (_04198_, _04197_);
  nor _55665_ (_04199_, _04198_, _04186_);
  and _55666_ (_04200_, _04199_, _04185_);
  nor _55667_ (_04201_, _04192_, _03471_);
  or _55668_ (_04202_, _04201_, _04200_);
  and _55669_ (_04203_, _04202_, _03152_);
  or _55670_ (_04204_, _04203_, _03434_);
  and _55671_ (_04205_, _03489_, _03165_);
  and _55672_ (_04206_, _04205_, _03043_);
  and _55673_ (_04207_, _03969_, _03043_);
  nor _55674_ (_04208_, _04207_, _04206_);
  and _55675_ (_04209_, _03650_, _03165_);
  nor _55676_ (_04210_, _04209_, _03520_);
  and _55677_ (_04211_, _03633_, _03165_);
  and _55678_ (_04212_, _04004_, _03165_);
  nor _55679_ (_04213_, _04212_, _04211_);
  and _55680_ (_04214_, _04213_, _04210_);
  and _55681_ (_04215_, _04214_, _04208_);
  nand _55682_ (_04216_, _04215_, _04204_);
  and _55683_ (_04217_, _04216_, _03996_);
  nand _55684_ (_04218_, _04217_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _55685_ (_04219_, _03385_, _41676_);
  nor _55686_ (_04220_, _03396_, _41724_);
  nor _55687_ (_04221_, _04220_, _04219_);
  nor _55688_ (_04222_, _03367_, _42183_);
  nor _55689_ (_04223_, _03391_, _41896_);
  nor _55690_ (_04224_, _04223_, _04222_);
  and _55691_ (_04225_, _04224_, _04221_);
  nor _55692_ (_04226_, _03359_, _41773_);
  nor _55693_ (_04227_, _03373_, _41814_);
  nor _55694_ (_04228_, _04227_, _04226_);
  nor _55695_ (_04229_, _03394_, _42101_);
  nor _55696_ (_04230_, _03380_, _41978_);
  nor _55697_ (_04231_, _04230_, _04229_);
  and _55698_ (_04232_, _04231_, _04228_);
  and _55699_ (_04233_, _04232_, _04225_);
  nor _55700_ (_04234_, _03345_, _42265_);
  nor _55701_ (_04235_, _03365_, _42224_);
  nor _55702_ (_04236_, _04235_, _04234_);
  nor _55703_ (_04237_, _03389_, _42142_);
  nor _55704_ (_04238_, _03351_, _42019_);
  nor _55705_ (_04239_, _04238_, _04237_);
  and _55706_ (_04240_, _04239_, _04236_);
  nor _55707_ (_04241_, _03378_, _42060_);
  nor _55708_ (_04242_, _03383_, _41635_);
  nor _55709_ (_04243_, _04242_, _04241_);
  nor _55710_ (_04244_, _03370_, _41937_);
  nor _55711_ (_04245_, _03356_, _41855_);
  nor _55712_ (_04246_, _04245_, _04244_);
  and _55713_ (_04247_, _04246_, _04243_);
  and _55714_ (_04248_, _04247_, _04240_);
  and _55715_ (_04249_, _04248_, _04233_);
  nor _55716_ (_04250_, _04249_, _03401_);
  and _55717_ (_04251_, _04250_, _03151_);
  not _55718_ (_04252_, _04251_);
  nor _55719_ (_04253_, _03365_, _42209_);
  nor _55720_ (_04254_, _03367_, _42168_);
  nor _55721_ (_04255_, _04254_, _04253_);
  nor _55722_ (_04256_, _03370_, _41922_);
  nor _55723_ (_04257_, _03359_, _41758_);
  nor _55724_ (_04258_, _04257_, _04256_);
  and _55725_ (_04259_, _04258_, _04255_);
  nor _55726_ (_04260_, _03391_, _41881_);
  nor _55727_ (_04261_, _03373_, _41799_);
  nor _55728_ (_04262_, _04261_, _04260_);
  nor _55729_ (_04263_, _03356_, _41840_);
  nor _55730_ (_04264_, _03383_, _41620_);
  nor _55731_ (_04265_, _04264_, _04263_);
  and _55732_ (_04266_, _04265_, _04262_);
  and _55733_ (_04267_, _04266_, _04259_);
  nor _55734_ (_04268_, _03378_, _42045_);
  nor _55735_ (_04269_, _03380_, _41963_);
  nor _55736_ (_04270_, _04269_, _04268_);
  nor _55737_ (_04271_, _03345_, _42250_);
  nor _55738_ (_04272_, _03389_, _42127_);
  nor _55739_ (_04273_, _04272_, _04271_);
  and _55740_ (_04274_, _04273_, _04270_);
  nor _55741_ (_04276_, _03396_, _41706_);
  nor _55742_ (_04277_, _03385_, _41661_);
  nor _55743_ (_04278_, _04277_, _04276_);
  nor _55744_ (_04279_, _03394_, _42086_);
  nor _55745_ (_04280_, _03351_, _42004_);
  nor _55746_ (_04281_, _04280_, _04279_);
  and _55747_ (_04282_, _04281_, _04278_);
  and _55748_ (_04283_, _04282_, _04274_);
  and _55749_ (_04284_, _04283_, _04267_);
  nor _55750_ (_04285_, _04284_, _03887_);
  not _55751_ (_04286_, _04285_);
  and _55752_ (_04287_, _03698_, _01931_);
  and _55753_ (_04288_, _03721_, _01890_);
  nor _55754_ (_04289_, _04288_, _04287_);
  and _55755_ (_04290_, _03689_, _01888_);
  and _55756_ (_04291_, _03737_, _01925_);
  nor _55757_ (_04292_, _04291_, _04290_);
  and _55758_ (_04293_, _04292_, _04289_);
  and _55759_ (_04294_, _03726_, _01929_);
  and _55760_ (_04295_, _03704_, _01912_);
  nor _55761_ (_04296_, _04295_, _04294_);
  and _55762_ (_04297_, _03724_, _01885_);
  and _55763_ (_04298_, _03700_, _01896_);
  nor _55764_ (_04299_, _04298_, _04297_);
  and _55765_ (_04300_, _04299_, _04296_);
  and _55766_ (_04301_, _04300_, _04293_);
  and _55767_ (_04302_, _03719_, _01898_);
  and _55768_ (_04303_, _03693_, _01908_);
  nor _55769_ (_04304_, _04303_, _04302_);
  and _55770_ (_04305_, _03711_, _01920_);
  and _55771_ (_04306_, _03713_, _01905_);
  nor _55772_ (_04307_, _04306_, _04305_);
  and _55773_ (_04308_, _04307_, _04304_);
  and _55774_ (_04309_, _03732_, _01922_);
  and _55775_ (_04310_, _03707_, _01902_);
  nor _55776_ (_04311_, _04310_, _04309_);
  and _55777_ (_04312_, _03730_, _01914_);
  and _55778_ (_04313_, _03735_, _01927_);
  nor _55779_ (_04314_, _04313_, _04312_);
  and _55780_ (_04315_, _04314_, _04311_);
  and _55781_ (_04316_, _04315_, _04308_);
  and _55782_ (_04317_, _04316_, _04301_);
  nor _55783_ (_04318_, _04317_, _03474_);
  and _55784_ (_04319_, _03489_, _03182_);
  not _55785_ (_04320_, _04319_);
  and _55786_ (_04321_, _03482_, _03515_);
  and _55787_ (_04322_, _03489_, _03171_);
  nor _55788_ (_04323_, _04322_, _04321_);
  and _55789_ (_04324_, _04323_, _04320_);
  and _55790_ (_04325_, _03661_, _03193_);
  nor _55791_ (_04326_, _04325_, _04151_);
  and _55792_ (_04327_, _03661_, _03177_);
  and _55793_ (_04328_, _03489_, _03010_);
  nor _55794_ (_04329_, _04328_, _04327_);
  and _55795_ (_04330_, _04329_, _04326_);
  and _55796_ (_04331_, _04330_, _04324_);
  and _55797_ (_04332_, _04331_, _03956_);
  not _55798_ (_04333_, \oc8051_golden_model_1.SP [1]);
  nor _55799_ (_04334_, _03985_, _04333_);
  not _55800_ (_04335_, _04334_);
  not _55801_ (_04336_, _03489_);
  and _55802_ (_04337_, _03253_, _03207_);
  nor _55803_ (_04338_, _04337_, _04336_);
  not _55804_ (_04339_, _04338_);
  and _55805_ (_04340_, _03489_, _03515_);
  nor _55806_ (_04341_, _04340_, _04205_);
  not _55807_ (_04342_, _04341_);
  nor _55808_ (_04343_, _04342_, _03963_);
  and _55809_ (_04344_, _04343_, _04339_);
  and _55810_ (_04345_, _03489_, _03191_);
  nor _55811_ (_04346_, _04345_, _03938_);
  and _55812_ (_04347_, _03663_, _03193_);
  and _55813_ (_04348_, _03489_, _03504_);
  nor _55814_ (_04349_, _04348_, _04347_);
  and _55815_ (_04350_, _04349_, _04346_);
  nor _55816_ (_04351_, _03490_, _03922_);
  nor _55817_ (_04352_, _04033_, _03934_);
  and _55818_ (_04353_, _04352_, _04351_);
  and _55819_ (_04354_, _04353_, _04350_);
  and _55820_ (_04355_, _04354_, _04344_);
  and _55821_ (_04356_, _04355_, _04335_);
  and _55822_ (_04357_, _04356_, _04332_);
  not _55823_ (_04358_, _04357_);
  nor _55824_ (_04359_, _04358_, _04318_);
  and _55825_ (_04360_, _04359_, _04286_);
  and _55826_ (_04361_, _04360_, _04252_);
  and _55827_ (_04362_, _04250_, _03499_);
  and _55828_ (_04363_, _03841_, _03629_);
  and _55829_ (_04364_, _04363_, _03840_);
  not _55830_ (_04365_, _04364_);
  and _55831_ (_04366_, _04365_, _04250_);
  nor _55832_ (_04367_, _04366_, _04362_);
  and _55833_ (_04368_, _04367_, _04361_);
  not _55834_ (_04369_, \oc8051_golden_model_1.IRAM[1] [0]);
  or _55835_ (_04370_, _04217_, _04369_);
  and _55836_ (_04371_, _04370_, _04368_);
  nand _55837_ (_04372_, _04371_, _04218_);
  nand _55838_ (_04373_, _04216_, _03996_);
  nand _55839_ (_04374_, _04373_, \oc8051_golden_model_1.IRAM[3] [0]);
  not _55840_ (_04375_, _04368_);
  nand _55841_ (_04377_, _04217_, \oc8051_golden_model_1.IRAM[2] [0]);
  and _55842_ (_04378_, _04377_, _04375_);
  nand _55843_ (_04379_, _04378_, _04374_);
  nand _55844_ (_04380_, _04379_, _04372_);
  nand _55845_ (_04381_, _04380_, _03994_);
  not _55846_ (_04382_, _03994_);
  nand _55847_ (_04383_, _04373_, \oc8051_golden_model_1.IRAM[7] [0]);
  nand _55848_ (_04384_, _04217_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _55849_ (_04385_, _04384_, _04375_);
  nand _55850_ (_04386_, _04385_, _04383_);
  nand _55851_ (_04387_, _04217_, \oc8051_golden_model_1.IRAM[4] [0]);
  not _55852_ (_04388_, \oc8051_golden_model_1.IRAM[5] [0]);
  or _55853_ (_04389_, _04217_, _04388_);
  and _55854_ (_04390_, _04389_, _04368_);
  nand _55855_ (_04391_, _04390_, _04387_);
  nand _55856_ (_04392_, _04391_, _04386_);
  nand _55857_ (_04393_, _04392_, _04382_);
  nand _55858_ (_04394_, _04393_, _04381_);
  nand _55859_ (_04395_, _04394_, _03803_);
  not _55860_ (_04396_, _03803_);
  nand _55861_ (_04397_, _04373_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _55862_ (_04398_, _04217_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _55863_ (_04399_, _04398_, _04375_);
  nand _55864_ (_04400_, _04399_, _04397_);
  nand _55865_ (_04401_, _04217_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand _55866_ (_04402_, _04373_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _55867_ (_04403_, _04402_, _04368_);
  nand _55868_ (_04404_, _04403_, _04401_);
  nand _55869_ (_04405_, _04404_, _04400_);
  nand _55870_ (_04406_, _04405_, _03994_);
  nand _55871_ (_04407_, _04373_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _55872_ (_04408_, _04217_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _55873_ (_04409_, _04408_, _04375_);
  nand _55874_ (_04410_, _04409_, _04407_);
  nand _55875_ (_04411_, _04217_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand _55876_ (_04412_, _04373_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _55877_ (_04413_, _04412_, _04368_);
  nand _55878_ (_04414_, _04413_, _04411_);
  nand _55879_ (_04415_, _04414_, _04410_);
  nand _55880_ (_04416_, _04415_, _04382_);
  nand _55881_ (_04417_, _04416_, _04406_);
  nand _55882_ (_04418_, _04417_, _04396_);
  and _55883_ (_04419_, _04418_, _04395_);
  and _55884_ (_04420_, _04419_, _03519_);
  nor _55885_ (_04421_, _03637_, _03159_);
  and _55886_ (_04422_, _04421_, _04005_);
  nor _55887_ (_04423_, _04422_, _03210_);
  not _55888_ (_04424_, _04423_);
  nor _55889_ (_04425_, _04424_, _04420_);
  and _55890_ (_04426_, _03655_, _03571_);
  not _55891_ (_04427_, _04426_);
  nor _55892_ (_04428_, _04427_, _03401_);
  and _55893_ (_04429_, _04428_, _03471_);
  nor _55894_ (_04430_, _04429_, _04425_);
  and _55895_ (_04431_, _03923_, \oc8051_golden_model_1.SP [0]);
  not _55896_ (_04432_, _04431_);
  and _55897_ (_04433_, _03487_, _03515_);
  not _55898_ (_04434_, _04433_);
  and _55899_ (_04435_, _04021_, _04434_);
  and _55900_ (_04436_, _04435_, _04432_);
  and _55901_ (_04437_, _04436_, _04430_);
  and _55902_ (_04438_, _03478_, _03515_);
  nand _55903_ (_04439_, _04418_, _04395_);
  and _55904_ (_04440_, _04439_, _04438_);
  not _55905_ (_04441_, _04440_);
  and _55906_ (_04442_, _04441_, _04437_);
  nor _55907_ (_04443_, _03517_, _03401_);
  not _55908_ (_04444_, _03570_);
  nor _55909_ (_04445_, _04444_, _03401_);
  and _55910_ (_04446_, _04445_, _03471_);
  nor _55911_ (_04447_, _04446_, _04443_);
  and _55912_ (_04448_, _04447_, _04442_);
  not _55913_ (_04449_, _04448_);
  and _55914_ (_04450_, _04449_, _03518_);
  nor _55915_ (_04451_, _03203_, _03502_);
  nor _55916_ (_04452_, _04451_, _04450_);
  and _55917_ (_04453_, _04141_, _03510_);
  nor _55918_ (_04454_, _03983_, _03401_);
  and _55919_ (_04455_, _04454_, _03471_);
  nor _55920_ (_04456_, _04455_, _04453_);
  and _55921_ (_04457_, _04456_, _04452_);
  and _55922_ (_04458_, _03478_, _03510_);
  and _55923_ (_04459_, _04458_, _04439_);
  not _55924_ (_04460_, _04459_);
  and _55925_ (_04461_, _04460_, _04457_);
  nor _55926_ (_04462_, _03513_, _03401_);
  nor _55927_ (_04463_, _03583_, _03401_);
  and _55928_ (_04464_, _04463_, _03471_);
  nor _55929_ (_04465_, _04464_, _04462_);
  and _55930_ (_04466_, _04465_, _04461_);
  nor _55931_ (_04467_, _04466_, _03514_);
  or _55932_ (_04468_, _04467_, _03511_);
  nand _55933_ (_04469_, _03511_, _03502_);
  nand _55934_ (_04470_, _04469_, _04468_);
  and _55935_ (_04471_, _04470_, _03509_);
  nor _55936_ (_04472_, _04471_, _03507_);
  and _55937_ (_04473_, _04141_, _03596_);
  or _55938_ (_04474_, _04473_, _04472_);
  nor _55939_ (_04475_, _04474_, _03503_);
  nor _55940_ (_04476_, _03500_, _03401_);
  and _55941_ (_04478_, _03478_, _03596_);
  and _55942_ (_04479_, _04439_, _04478_);
  nor _55943_ (_04480_, _04479_, _04476_);
  and _55944_ (_04481_, _04480_, _04475_);
  nor _55945_ (_04482_, _04481_, _03501_);
  nor _55946_ (_04483_, _04482_, _03223_);
  and _55947_ (_04484_, _03223_, _03502_);
  nor _55948_ (_04485_, _04484_, _04483_);
  and _55949_ (_04486_, _04141_, _03188_);
  or _55950_ (_04487_, _04486_, _04485_);
  nor _55951_ (_04488_, _04487_, _03496_);
  and _55952_ (_04489_, _03478_, _03188_);
  and _55953_ (_04490_, _04489_, _04439_);
  nor _55954_ (_04491_, _04490_, _03439_);
  and _55955_ (_04492_, _04491_, _04488_);
  nor _55956_ (_04493_, _04492_, _03473_);
  nor _55957_ (_04494_, _04493_, _03189_);
  and _55958_ (_04495_, _03189_, _03502_);
  nor _55959_ (_04496_, _04495_, _04494_);
  nor _55960_ (_04497_, _03753_, _03401_);
  not _55961_ (_04498_, _04497_);
  not _55962_ (_04499_, _03636_);
  nor _55963_ (_04500_, _04499_, _03401_);
  not _55964_ (_04501_, _03769_);
  nor _55965_ (_04502_, _04501_, _03401_);
  nor _55966_ (_04503_, _04502_, _04500_);
  and _55967_ (_04504_, _03644_, _03162_);
  not _55968_ (_04505_, _04504_);
  nor _55969_ (_04506_, _04505_, _03401_);
  not _55970_ (_04507_, _04506_);
  and _55971_ (_04508_, _04507_, _04503_);
  and _55972_ (_04509_, _04508_, _04498_);
  nor _55973_ (_04510_, _04509_, _03472_);
  nor _55974_ (_04511_, _04510_, _03192_);
  not _55975_ (_04512_, _04511_);
  nor _55976_ (_04513_, _04512_, _04496_);
  and _55977_ (_04514_, _03192_, _03502_);
  nor _55978_ (_04515_, _04514_, _04513_);
  nor _55979_ (_04516_, _03759_, _03401_);
  not _55980_ (_04517_, _03760_);
  nor _55981_ (_04518_, _04517_, _03401_);
  nor _55982_ (_04519_, _04518_, _04516_);
  nor _55983_ (_04520_, _04519_, _03472_);
  nor _55984_ (_04521_, _04520_, _04515_);
  and _55985_ (_04522_, _04141_, _03010_);
  and _55986_ (_04523_, _03179_, \oc8051_golden_model_1.SP [0]);
  nor _55987_ (_04524_, _04523_, _04522_);
  and _55988_ (_04525_, _04524_, _04521_);
  nor _55989_ (_04526_, _04192_, _03401_);
  and _55990_ (_04527_, _03478_, _03010_);
  and _55991_ (_04528_, _04439_, _04527_);
  nor _55992_ (_04529_, _04528_, _04526_);
  and _55993_ (_04530_, _04529_, _04525_);
  and _55994_ (_04531_, _04526_, _03472_);
  nor _55995_ (_04532_, _04531_, _04530_);
  nor _55996_ (_04533_, _03641_, _03160_);
  nor _55997_ (_04534_, _04533_, _03502_);
  nor _55998_ (_04535_, _04534_, _04532_);
  and _55999_ (_04536_, _04535_, _03436_);
  nor _56000_ (_04537_, _04536_, _03434_);
  and _56001_ (_04538_, _04141_, _03165_);
  nor _56002_ (_04539_, _04538_, _04537_);
  and _56003_ (_04540_, _03478_, _03165_);
  and _56004_ (_04541_, _04540_, _04439_);
  not _56005_ (_04542_, _04541_);
  and _56006_ (_04543_, _04542_, _04539_);
  nor _56007_ (_04544_, _03521_, _03401_);
  and _56008_ (_04545_, _04544_, _03471_);
  not _56009_ (_04546_, _04545_);
  and _56010_ (_04547_, _04546_, _04543_);
  not _56011_ (_04548_, _04284_);
  and _56012_ (_04549_, _04544_, _04548_);
  and _56013_ (_04550_, _04333_, \oc8051_golden_model_1.SP [0]);
  and _56014_ (_04551_, \oc8051_golden_model_1.SP [1], _03502_);
  nor _56015_ (_04552_, _04551_, _04550_);
  not _56016_ (_04553_, _04552_);
  nor _56017_ (_04554_, _04553_, _04533_);
  and _56018_ (_04555_, _04553_, _03179_);
  and _56019_ (_04556_, _04548_, _03439_);
  and _56020_ (_04557_, _03478_, _04010_);
  nand _56021_ (_04558_, _04217_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand _56022_ (_04559_, _04373_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _56023_ (_04560_, _04559_, _04368_);
  nand _56024_ (_04561_, _04560_, _04558_);
  nand _56025_ (_04562_, _04373_, \oc8051_golden_model_1.IRAM[3] [1]);
  nand _56026_ (_04563_, _04217_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _56027_ (_04564_, _04563_, _04375_);
  nand _56028_ (_04565_, _04564_, _04562_);
  nand _56029_ (_04566_, _04565_, _04561_);
  nand _56030_ (_04567_, _04566_, _03994_);
  nand _56031_ (_04568_, _04373_, \oc8051_golden_model_1.IRAM[7] [1]);
  nand _56032_ (_04569_, _04217_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _56033_ (_04570_, _04569_, _04375_);
  nand _56034_ (_04571_, _04570_, _04568_);
  nand _56035_ (_04572_, _04217_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand _56036_ (_04573_, _04373_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _56037_ (_04574_, _04573_, _04368_);
  nand _56038_ (_04575_, _04574_, _04572_);
  nand _56039_ (_04576_, _04575_, _04571_);
  nand _56040_ (_04577_, _04576_, _04382_);
  nand _56041_ (_04579_, _04577_, _04567_);
  nand _56042_ (_04580_, _04579_, _03803_);
  nand _56043_ (_04581_, _04373_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _56044_ (_04582_, _04217_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _56045_ (_04583_, _04582_, _04375_);
  nand _56046_ (_04584_, _04583_, _04581_);
  nand _56047_ (_04585_, _04217_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand _56048_ (_04586_, _04373_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _56049_ (_04587_, _04586_, _04368_);
  nand _56050_ (_04588_, _04587_, _04585_);
  nand _56051_ (_04589_, _04588_, _04584_);
  nand _56052_ (_04590_, _04589_, _03994_);
  nand _56053_ (_04591_, _04373_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _56054_ (_04592_, _04217_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _56055_ (_04593_, _04592_, _04375_);
  nand _56056_ (_04594_, _04593_, _04591_);
  nand _56057_ (_04595_, _04217_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand _56058_ (_04596_, _04373_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _56059_ (_04597_, _04596_, _04368_);
  nand _56060_ (_04598_, _04597_, _04595_);
  nand _56061_ (_04599_, _04598_, _04594_);
  nand _56062_ (_04600_, _04599_, _04382_);
  nand _56063_ (_04601_, _04600_, _04590_);
  nand _56064_ (_04602_, _04601_, _04396_);
  nand _56065_ (_04603_, _04602_, _04580_);
  and _56066_ (_04604_, _04603_, _03519_);
  or _56067_ (_04605_, _04604_, _04557_);
  and _56068_ (_04606_, _04428_, _04284_);
  or _56069_ (_04607_, _04606_, _04605_);
  and _56070_ (_04608_, _04552_, _03923_);
  not _56071_ (_04609_, _04608_);
  and _56072_ (_04610_, _03476_, _03515_);
  and _56073_ (_04611_, _03925_, _03515_);
  nor _56074_ (_04612_, _04611_, _04610_);
  and _56075_ (_04613_, _04612_, _04609_);
  not _56076_ (_04614_, _04613_);
  nor _56077_ (_04615_, _04614_, _04607_);
  and _56078_ (_04616_, _04603_, _04438_);
  nor _56079_ (_04617_, _04616_, _04445_);
  and _56080_ (_04618_, _04617_, _04615_);
  and _56081_ (_04619_, _04445_, _04548_);
  nor _56082_ (_04620_, _04619_, _04618_);
  and _56083_ (_04621_, _04249_, _04443_);
  nor _56084_ (_04622_, _04621_, _04620_);
  or _56085_ (_04623_, _04553_, _03203_);
  nand _56086_ (_04624_, _04623_, _04622_);
  and _56087_ (_04625_, _04454_, _04284_);
  and _56088_ (_04626_, _03476_, _03510_);
  nor _56089_ (_04627_, _04626_, _03978_);
  not _56090_ (_04628_, _04627_);
  nor _56091_ (_04629_, _04628_, _04625_);
  not _56092_ (_04630_, _04629_);
  nor _56093_ (_04631_, _04630_, _04624_);
  and _56094_ (_04632_, _04603_, _04458_);
  nor _56095_ (_04633_, _04632_, _04463_);
  and _56096_ (_04634_, _04633_, _04631_);
  and _56097_ (_04635_, _04463_, _04548_);
  nor _56098_ (_04636_, _04635_, _04634_);
  and _56099_ (_04637_, _04249_, _04462_);
  or _56100_ (_04638_, _04637_, _03511_);
  nor _56101_ (_04639_, _04638_, _04636_);
  and _56102_ (_04640_, _04553_, _03511_);
  nor _56103_ (_04641_, _04640_, _04639_);
  and _56104_ (_04642_, _03508_, _04249_);
  nor _56105_ (_04643_, _04642_, _04641_);
  nor _56106_ (_04644_, _04553_, _03200_);
  nor _56107_ (_04645_, _03476_, _03925_);
  nor _56108_ (_04646_, _04645_, _03212_);
  nor _56109_ (_04647_, _04646_, _04644_);
  and _56110_ (_04648_, _04647_, _04643_);
  and _56111_ (_04649_, _04603_, _04478_);
  nor _56112_ (_04650_, _04649_, _04476_);
  and _56113_ (_04651_, _04650_, _04648_);
  nor _56114_ (_04652_, _04651_, _04362_);
  nor _56115_ (_04653_, _04652_, _03223_);
  and _56116_ (_04654_, _04553_, _03223_);
  nor _56117_ (_04655_, _04654_, _04653_);
  and _56118_ (_04656_, _03495_, _04284_);
  not _56119_ (_04657_, _03188_);
  nor _56120_ (_04658_, _04645_, _04657_);
  nor _56121_ (_04659_, _04658_, _04656_);
  not _56122_ (_04660_, _04659_);
  nor _56123_ (_04661_, _04660_, _04655_);
  and _56124_ (_04662_, _04603_, _04489_);
  nor _56125_ (_04663_, _04662_, _03439_);
  and _56126_ (_04664_, _04663_, _04661_);
  nor _56127_ (_04665_, _04664_, _04556_);
  nor _56128_ (_04666_, _04665_, _03189_);
  and _56129_ (_04667_, _04553_, _03189_);
  nor _56130_ (_04668_, _04667_, _04666_);
  nor _56131_ (_04669_, _04509_, _04548_);
  nor _56132_ (_04670_, _04669_, _03192_);
  not _56133_ (_04671_, _04670_);
  nor _56134_ (_04672_, _04671_, _04668_);
  and _56135_ (_04673_, _04553_, _03192_);
  nor _56136_ (_04674_, _04673_, _04672_);
  nor _56137_ (_04675_, _04519_, _04548_);
  nor _56138_ (_04676_, _04675_, _03179_);
  not _56139_ (_04677_, _04676_);
  nor _56140_ (_04678_, _04677_, _04674_);
  nor _56141_ (_04680_, _04678_, _04555_);
  and _56142_ (_04681_, _03476_, _03010_);
  nor _56143_ (_04682_, _04681_, _03970_);
  not _56144_ (_04683_, _04682_);
  nor _56145_ (_04684_, _04683_, _04680_);
  and _56146_ (_04685_, _04603_, _04527_);
  nor _56147_ (_04686_, _04685_, _04526_);
  and _56148_ (_04687_, _04686_, _04684_);
  and _56149_ (_04688_, _04526_, _04548_);
  nor _56150_ (_04689_, _04688_, _04687_);
  or _56151_ (_04690_, _04689_, _03435_);
  nor _56152_ (_04691_, _04690_, _04554_);
  nor _56153_ (_04692_, _04691_, _04251_);
  and _56154_ (_04693_, _03476_, _03165_);
  nor _56155_ (_04694_, _04693_, _03969_);
  not _56156_ (_04695_, _04694_);
  nor _56157_ (_04696_, _04695_, _04692_);
  and _56158_ (_04697_, _04603_, _04540_);
  nor _56159_ (_04698_, _04697_, _04544_);
  and _56160_ (_04699_, _04698_, _04696_);
  nor _56161_ (_04700_, _04699_, _04549_);
  not _56162_ (_04701_, _00000_);
  nor _56163_ (_04702_, _03508_, _04454_);
  nor _56164_ (_04703_, _04463_, _04428_);
  and _56165_ (_04704_, _04703_, _04702_);
  and _56166_ (_04705_, _03484_, _03010_);
  not _56167_ (_04706_, _04705_);
  and _56168_ (_04707_, _03661_, _03010_);
  nor _56169_ (_04708_, _04707_, _04189_);
  and _56170_ (_04709_, _04708_, _04706_);
  and _56171_ (_04710_, _03664_, _03510_);
  nor _56172_ (_04711_, _04710_, _04033_);
  nor _56173_ (_04712_, _03478_, _03476_);
  nor _56174_ (_04713_, _04712_, _03210_);
  nor _56175_ (_04714_, _04713_, _04342_);
  and _56176_ (_04715_, _04714_, _04711_);
  and _56177_ (_04716_, _04715_, _04709_);
  and _56178_ (_04717_, _04716_, _03980_);
  not _56179_ (_04718_, _03220_);
  and _56180_ (_04719_, _04421_, _04718_);
  nor _56181_ (_04720_, _04719_, _03210_);
  nor _56182_ (_04721_, _04540_, _04209_);
  not _56183_ (_04722_, _04721_);
  nor _56184_ (_04723_, _04722_, _04720_);
  and _56185_ (_04724_, _04142_, _03188_);
  and _56186_ (_04725_, _03483_, _03188_);
  or _56187_ (_04726_, _04725_, _04724_);
  not _56188_ (_04727_, _04726_);
  nand _56189_ (_04728_, _03489_, _03188_);
  nand _56190_ (_04729_, _03476_, _03188_);
  or _56191_ (_04730_, _04729_, _03043_);
  and _56192_ (_04731_, _04730_, _04728_);
  and _56193_ (_04732_, _04731_, _04727_);
  and _56194_ (_04733_, _04732_, _04723_);
  nor _56195_ (_04734_, _04610_, _04681_);
  and _56196_ (_04735_, _03476_, _03596_);
  nor _56197_ (_04736_, _04438_, _04735_);
  and _56198_ (_04737_, _04736_, _04734_);
  nor _56199_ (_04738_, _04489_, _04527_);
  and _56200_ (_04739_, _03655_, _03188_);
  nor _56201_ (_04740_, _04739_, _03943_);
  and _56202_ (_04741_, _04740_, _04738_);
  and _56203_ (_04742_, _04741_, _04737_);
  not _56204_ (_04743_, _03200_);
  or _56205_ (_04744_, _03223_, _04743_);
  not _56206_ (_04745_, _04744_);
  not _56207_ (_04746_, _03203_);
  nor _56208_ (_04747_, _04746_, _03189_);
  and _56209_ (_04748_, _04747_, _04745_);
  and _56210_ (_04749_, _03650_, _03510_);
  not _56211_ (_04750_, _04749_);
  nor _56212_ (_04751_, _04458_, _03511_);
  and _56213_ (_04752_, _04751_, _04750_);
  and _56214_ (_04753_, _04752_, _04748_);
  and _56215_ (_04754_, _04753_, _04742_);
  nor _56216_ (_04755_, _03192_, _03179_);
  not _56217_ (_04756_, _03599_);
  and _56218_ (_04757_, _04756_, _04755_);
  and _56219_ (_04758_, _03650_, _03188_);
  and _56220_ (_04759_, _03664_, _03165_);
  nor _56221_ (_04760_, _04759_, _04758_);
  and _56222_ (_04761_, _04760_, _04757_);
  not _56223_ (_04762_, _03923_);
  and _56224_ (_04763_, _04533_, _04762_);
  and _56225_ (_04764_, _03489_, _03596_);
  nor _56226_ (_04765_, _04764_, _03597_);
  and _56227_ (_04766_, _03481_, _03165_);
  nor _56228_ (_04767_, _04478_, _04766_);
  and _56229_ (_04768_, _04767_, _04765_);
  and _56230_ (_04769_, _04768_, _04763_);
  and _56231_ (_04770_, _04769_, _04761_);
  and _56232_ (_04771_, _04770_, _04754_);
  and _56233_ (_04772_, _04771_, _04733_);
  and _56234_ (_04773_, _04772_, _04717_);
  not _56235_ (_04774_, _04773_);
  nor _56236_ (_04775_, _03752_, _03520_);
  and _56237_ (_04776_, _04775_, _03486_);
  and _56238_ (_04777_, _04776_, _03480_);
  and _56239_ (_04778_, _04777_, _03491_);
  nor _56240_ (_04779_, _04778_, _03401_);
  nor _56241_ (_04781_, _04779_, _04774_);
  and _56242_ (_04782_, _04781_, _04519_);
  and _56243_ (_04783_, _04782_, _04704_);
  nor _56244_ (_04784_, _03401_, _03474_);
  nor _56245_ (_04785_, _04784_, _04462_);
  nor _56246_ (_04786_, _04445_, _04476_);
  and _56247_ (_04787_, _04786_, _04785_);
  nor _56248_ (_04788_, _04526_, _03435_);
  nor _56249_ (_04789_, _04443_, _03439_);
  and _56250_ (_04790_, _04789_, _04788_);
  and _56251_ (_04791_, _04790_, _04787_);
  and _56252_ (_04792_, _04791_, _04508_);
  and _56253_ (_04793_, _04792_, _04783_);
  nor _56254_ (_04794_, _04793_, _04701_);
  not _56255_ (_04795_, _04794_);
  nor _56256_ (_04796_, _04795_, _04700_);
  and _56257_ (_04797_, _04796_, _04547_);
  not _56258_ (_04798_, \oc8051_golden_model_1.IRAM[0] [3]);
  or _56259_ (_04799_, _04373_, _04798_);
  nand _56260_ (_04800_, _04373_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _56261_ (_04801_, _04800_, _04368_);
  nand _56262_ (_04802_, _04801_, _04799_);
  nand _56263_ (_04803_, _04373_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand _56264_ (_04804_, _04217_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _56265_ (_04805_, _04804_, _04375_);
  nand _56266_ (_04806_, _04805_, _04803_);
  nand _56267_ (_04807_, _04806_, _04802_);
  nand _56268_ (_04808_, _04807_, _03994_);
  nand _56269_ (_04809_, _04373_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand _56270_ (_04810_, _04217_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _56271_ (_04811_, _04810_, _04375_);
  nand _56272_ (_04812_, _04811_, _04809_);
  nand _56273_ (_04813_, _04217_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand _56274_ (_04814_, _04373_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _56275_ (_04815_, _04814_, _04368_);
  nand _56276_ (_04816_, _04815_, _04813_);
  nand _56277_ (_04817_, _04816_, _04812_);
  nand _56278_ (_04818_, _04817_, _04382_);
  nand _56279_ (_04819_, _04818_, _04808_);
  nand _56280_ (_04820_, _04819_, _03803_);
  nand _56281_ (_04821_, _04373_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _56282_ (_04822_, _04217_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _56283_ (_04823_, _04822_, _04375_);
  nand _56284_ (_04824_, _04823_, _04821_);
  nand _56285_ (_04825_, _04217_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand _56286_ (_04826_, _04373_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _56287_ (_04827_, _04826_, _04368_);
  nand _56288_ (_04828_, _04827_, _04825_);
  nand _56289_ (_04829_, _04828_, _04824_);
  nand _56290_ (_04830_, _04829_, _03994_);
  nand _56291_ (_04831_, _04373_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _56292_ (_04832_, _04217_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _56293_ (_04833_, _04832_, _04375_);
  nand _56294_ (_04834_, _04833_, _04831_);
  nand _56295_ (_04835_, _04217_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand _56296_ (_04836_, _04373_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _56297_ (_04837_, _04836_, _04368_);
  nand _56298_ (_04838_, _04837_, _04835_);
  nand _56299_ (_04839_, _04838_, _04834_);
  nand _56300_ (_04840_, _04839_, _04382_);
  nand _56301_ (_04841_, _04840_, _04830_);
  nand _56302_ (_04842_, _04841_, _04396_);
  nand _56303_ (_04843_, _04842_, _04820_);
  and _56304_ (_04844_, _04843_, _04540_);
  and _56305_ (_04845_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _56306_ (_04846_, _04845_, \oc8051_golden_model_1.SP [2]);
  nor _56307_ (_04847_, _04846_, \oc8051_golden_model_1.SP [3]);
  and _56308_ (_04848_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _56309_ (_04849_, _04848_, \oc8051_golden_model_1.SP [3]);
  and _56310_ (_04850_, _04849_, \oc8051_golden_model_1.SP [0]);
  nor _56311_ (_04851_, _04850_, _04847_);
  and _56312_ (_04852_, _04851_, _03223_);
  not _56313_ (_04853_, _03223_);
  nand _56314_ (_04854_, _04443_, _03561_);
  nand _56315_ (_04855_, _04843_, _03519_);
  not _56316_ (_04856_, \oc8051_golden_model_1.PSW [3]);
  nand _56317_ (_04857_, _03211_, _04856_);
  and _56318_ (_04858_, _04857_, _04855_);
  or _56319_ (_04859_, _04858_, _04428_);
  nand _56320_ (_04860_, _04428_, _03432_);
  and _56321_ (_04861_, _04860_, _04762_);
  and _56322_ (_04862_, _04861_, _04859_);
  and _56323_ (_04863_, _04851_, _03923_);
  or _56324_ (_04864_, _04863_, _04438_);
  or _56325_ (_04865_, _04864_, _04862_);
  not _56326_ (_04866_, _04445_);
  nand _56327_ (_04867_, _04843_, _04438_);
  and _56328_ (_04868_, _04867_, _04866_);
  and _56329_ (_04869_, _04868_, _04865_);
  and _56330_ (_04870_, _04445_, _03563_);
  or _56331_ (_04871_, _04870_, _04443_);
  or _56332_ (_04872_, _04871_, _04869_);
  and _56333_ (_04873_, _04872_, _04854_);
  or _56334_ (_04874_, _04873_, _04746_);
  nor _56335_ (_04875_, _04851_, _03203_);
  nor _56336_ (_04876_, _04875_, _04454_);
  and _56337_ (_04877_, _04876_, _04874_);
  and _56338_ (_04878_, _04454_, _03563_);
  or _56339_ (_04879_, _04878_, _04458_);
  or _56340_ (_04880_, _04879_, _04877_);
  and _56341_ (_04881_, _04843_, _04458_);
  nor _56342_ (_04882_, _04881_, _04463_);
  and _56343_ (_04883_, _04882_, _04880_);
  and _56344_ (_04884_, _04463_, _03563_);
  or _56345_ (_04885_, _04884_, _04462_);
  or _56346_ (_04886_, _04885_, _04883_);
  not _56347_ (_04887_, _03511_);
  nand _56348_ (_04888_, _03561_, _04462_);
  and _56349_ (_04889_, _04888_, _04887_);
  and _56350_ (_04890_, _04889_, _04886_);
  and _56351_ (_04891_, _04851_, _03511_);
  or _56352_ (_04892_, _04891_, _03508_);
  or _56353_ (_04893_, _04892_, _04890_);
  nand _56354_ (_04894_, _03508_, _03561_);
  and _56355_ (_04895_, _04894_, _03200_);
  and _56356_ (_04896_, _04895_, _04893_);
  nor _56357_ (_04897_, _04478_, _04743_);
  nor _56358_ (_04898_, _04851_, _04478_);
  nor _56359_ (_04899_, _04898_, _04897_);
  or _56360_ (_04900_, _04899_, _04896_);
  not _56361_ (_04901_, _04476_);
  nand _56362_ (_04902_, _04843_, _04478_);
  and _56363_ (_04903_, _04902_, _04901_);
  and _56364_ (_04904_, _04903_, _04900_);
  nor _56365_ (_04905_, _04901_, _03565_);
  or _56366_ (_04906_, _04905_, _04904_);
  and _56367_ (_04907_, _04906_, _04853_);
  nor _56368_ (_04908_, _04907_, _04852_);
  or _56369_ (_04909_, _04908_, _03495_);
  not _56370_ (_04910_, _04489_);
  nand _56371_ (_04911_, _03495_, _03563_);
  and _56372_ (_04912_, _04911_, _04910_);
  and _56373_ (_04913_, _04912_, _04909_);
  and _56374_ (_04914_, _04843_, _04489_);
  nor _56375_ (_04915_, _04914_, _03439_);
  not _56376_ (_04916_, _04915_);
  nor _56377_ (_04917_, _04916_, _04913_);
  nor _56378_ (_04918_, _03438_, _03433_);
  nor _56379_ (_04919_, _04918_, _04917_);
  nor _56380_ (_04920_, _04919_, _03189_);
  and _56381_ (_04921_, _04851_, _03189_);
  not _56382_ (_04922_, _04921_);
  and _56383_ (_04923_, _04922_, _04509_);
  not _56384_ (_04924_, _04923_);
  nor _56385_ (_04925_, _04924_, _04920_);
  nor _56386_ (_04926_, _04509_, _03563_);
  nor _56387_ (_04927_, _04926_, _03192_);
  not _56388_ (_04928_, _04927_);
  nor _56389_ (_04929_, _04928_, _04925_);
  and _56390_ (_04930_, _04851_, _03192_);
  not _56391_ (_04931_, _04930_);
  and _56392_ (_04932_, _04931_, _04519_);
  not _56393_ (_04933_, _04932_);
  nor _56394_ (_04934_, _04933_, _04929_);
  nor _56395_ (_04935_, _04519_, _03563_);
  nor _56396_ (_04936_, _04935_, _03179_);
  not _56397_ (_04937_, _04936_);
  nor _56398_ (_04938_, _04937_, _04934_);
  and _56399_ (_04939_, _04851_, _03179_);
  nor _56400_ (_04940_, _04939_, _04527_);
  not _56401_ (_04941_, _04940_);
  nor _56402_ (_04942_, _04941_, _04938_);
  and _56403_ (_04943_, _04843_, _04527_);
  nor _56404_ (_04944_, _04943_, _04526_);
  not _56405_ (_04945_, _04944_);
  nor _56406_ (_04946_, _04945_, _04942_);
  not _56407_ (_04947_, _04533_);
  and _56408_ (_04948_, _04526_, _03563_);
  nor _56409_ (_04949_, _04948_, _04947_);
  not _56410_ (_04950_, _04949_);
  nor _56411_ (_04951_, _04950_, _04946_);
  nor _56412_ (_04952_, _04851_, _04533_);
  nor _56413_ (_04953_, _04952_, _03435_);
  not _56414_ (_04954_, _04953_);
  nor _56415_ (_04955_, _04954_, _04951_);
  not _56416_ (_04956_, _03561_);
  and _56417_ (_04957_, _03435_, _04956_);
  nor _56418_ (_04958_, _04957_, _04540_);
  not _56419_ (_04959_, _04958_);
  nor _56420_ (_04960_, _04959_, _04955_);
  or _56421_ (_04961_, _04960_, _04544_);
  nor _56422_ (_04962_, _04961_, _04844_);
  and _56423_ (_04963_, _04544_, _03563_);
  nor _56424_ (_04964_, _04963_, _04962_);
  not _56425_ (_04965_, _03877_);
  and _56426_ (_04966_, _04544_, _04965_);
  and _56427_ (_04967_, _03475_, _03165_);
  and _56428_ (_04968_, _03835_, _03151_);
  nor _56429_ (_04969_, _04845_, \oc8051_golden_model_1.SP [2]);
  nor _56430_ (_04970_, _04969_, _04846_);
  and _56431_ (_04971_, _04970_, _03179_);
  and _56432_ (_04972_, _04965_, _03439_);
  and _56433_ (_04973_, _03495_, _03877_);
  nor _56434_ (_04974_, _04970_, _03200_);
  nor _56435_ (_04975_, _04974_, _03600_);
  and _56436_ (_04976_, _04445_, _04965_);
  not _56437_ (_04977_, _04970_);
  and _56438_ (_04978_, _04977_, _03923_);
  and _56439_ (_04979_, _03475_, _03515_);
  nor _56440_ (_04980_, _04979_, _04978_);
  not _56441_ (_04981_, _04720_);
  nand _56442_ (_04982_, _04217_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand _56443_ (_04983_, _04373_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _56444_ (_04984_, _04983_, _04368_);
  nand _56445_ (_04985_, _04984_, _04982_);
  nand _56446_ (_04986_, _04373_, \oc8051_golden_model_1.IRAM[3] [2]);
  nand _56447_ (_04987_, _04217_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _56448_ (_04988_, _04987_, _04375_);
  nand _56449_ (_04989_, _04988_, _04986_);
  nand _56450_ (_04990_, _04989_, _04985_);
  nand _56451_ (_04991_, _04990_, _03994_);
  nand _56452_ (_04992_, _04373_, \oc8051_golden_model_1.IRAM[7] [2]);
  nand _56453_ (_04993_, _04217_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _56454_ (_04994_, _04993_, _04375_);
  nand _56455_ (_04995_, _04994_, _04992_);
  nand _56456_ (_04996_, _04217_, \oc8051_golden_model_1.IRAM[4] [2]);
  nand _56457_ (_04997_, _04373_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _56458_ (_04998_, _04997_, _04368_);
  nand _56459_ (_04999_, _04998_, _04996_);
  nand _56460_ (_05000_, _04999_, _04995_);
  nand _56461_ (_05001_, _05000_, _04382_);
  nand _56462_ (_05002_, _05001_, _04991_);
  nand _56463_ (_05003_, _05002_, _03803_);
  nand _56464_ (_05004_, _04373_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _56465_ (_05005_, _04217_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _56466_ (_05006_, _05005_, _04375_);
  nand _56467_ (_05007_, _05006_, _05004_);
  nand _56468_ (_05008_, _04217_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand _56469_ (_05009_, _04373_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _56470_ (_05010_, _05009_, _04368_);
  nand _56471_ (_05011_, _05010_, _05008_);
  nand _56472_ (_05012_, _05011_, _05007_);
  nand _56473_ (_05013_, _05012_, _03994_);
  nand _56474_ (_05014_, _04373_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _56475_ (_05015_, _04217_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _56476_ (_05016_, _05015_, _04375_);
  nand _56477_ (_05017_, _05016_, _05014_);
  nand _56478_ (_05018_, _04217_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand _56479_ (_05019_, _04373_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _56480_ (_05020_, _05019_, _04368_);
  nand _56481_ (_05021_, _05020_, _05018_);
  nand _56482_ (_05022_, _05021_, _05017_);
  nand _56483_ (_05023_, _05022_, _04382_);
  nand _56484_ (_05024_, _05023_, _05013_);
  nand _56485_ (_05025_, _05024_, _04396_);
  nand _56486_ (_05026_, _05025_, _05003_);
  nor _56487_ (_05027_, _05026_, _03158_);
  nor _56488_ (_05028_, _05027_, _04981_);
  and _56489_ (_05029_, _04428_, _03877_);
  nor _56490_ (_05030_, _05029_, _05028_);
  and _56491_ (_05031_, _05030_, _04980_);
  and _56492_ (_05032_, _05026_, _04438_);
  nor _56493_ (_05033_, _05032_, _04445_);
  and _56494_ (_05034_, _05033_, _05031_);
  nor _56495_ (_05035_, _05034_, _04976_);
  and _56496_ (_05036_, _04443_, _03834_);
  or _56497_ (_05037_, _05036_, _05035_);
  nor _56498_ (_05038_, _04970_, _03203_);
  or _56499_ (_05039_, _05038_, _05037_);
  and _56500_ (_05040_, _04454_, _03877_);
  and _56501_ (_05041_, _03475_, _03510_);
  nor _56502_ (_05042_, _05041_, _05040_);
  not _56503_ (_05043_, _05042_);
  nor _56504_ (_05044_, _05043_, _05039_);
  and _56505_ (_05045_, _05026_, _04458_);
  nor _56506_ (_05046_, _05045_, _04463_);
  and _56507_ (_05047_, _05046_, _05044_);
  and _56508_ (_05048_, _04463_, _04965_);
  nor _56509_ (_05049_, _05048_, _05047_);
  and _56510_ (_05050_, _03834_, _04462_);
  or _56511_ (_05051_, _05050_, _03511_);
  nor _56512_ (_05052_, _05051_, _05049_);
  and _56513_ (_05053_, _04970_, _03511_);
  nor _56514_ (_05054_, _05053_, _05052_);
  and _56515_ (_05055_, _03508_, _03834_);
  nor _56516_ (_05056_, _05055_, _05054_);
  and _56517_ (_05057_, _05056_, _04975_);
  and _56518_ (_05058_, _05026_, _04478_);
  nor _56519_ (_05059_, _05058_, _04476_);
  and _56520_ (_05060_, _05059_, _05057_);
  nor _56521_ (_05061_, _05060_, _03836_);
  nor _56522_ (_05062_, _05061_, _03223_);
  and _56523_ (_05063_, _04970_, _03223_);
  nor _56524_ (_05064_, _05063_, _05062_);
  and _56525_ (_05065_, _03475_, _03188_);
  or _56526_ (_05066_, _05065_, _05064_);
  nor _56527_ (_05067_, _05066_, _04973_);
  and _56528_ (_05068_, _05026_, _04489_);
  nor _56529_ (_05069_, _05068_, _03439_);
  and _56530_ (_05070_, _05069_, _05067_);
  nor _56531_ (_05071_, _05070_, _04972_);
  nor _56532_ (_05072_, _05071_, _03189_);
  and _56533_ (_05073_, _04970_, _03189_);
  nor _56534_ (_05074_, _05073_, _05072_);
  nor _56535_ (_05075_, _04509_, _04965_);
  nor _56536_ (_05076_, _05075_, _03192_);
  not _56537_ (_05077_, _05076_);
  nor _56538_ (_05078_, _05077_, _05074_);
  and _56539_ (_05079_, _04970_, _03192_);
  nor _56540_ (_05080_, _05079_, _05078_);
  nor _56541_ (_05081_, _04519_, _04965_);
  nor _56542_ (_05082_, _05081_, _03179_);
  not _56543_ (_05083_, _05082_);
  nor _56544_ (_05084_, _05083_, _05080_);
  nor _56545_ (_05085_, _05084_, _04971_);
  and _56546_ (_05086_, _03475_, _03010_);
  nor _56547_ (_05087_, _05086_, _05085_);
  and _56548_ (_05088_, _05026_, _04527_);
  nor _56549_ (_05089_, _05088_, _04526_);
  and _56550_ (_05090_, _05089_, _05087_);
  and _56551_ (_05091_, _04526_, _04965_);
  nor _56552_ (_05092_, _05091_, _05090_);
  nor _56553_ (_05093_, _04970_, _04533_);
  nor _56554_ (_05094_, _05093_, _03435_);
  not _56555_ (_05095_, _05094_);
  nor _56556_ (_05096_, _05095_, _05092_);
  nor _56557_ (_05097_, _05096_, _04968_);
  nor _56558_ (_05098_, _05097_, _04967_);
  and _56559_ (_05099_, _05026_, _04540_);
  nor _56560_ (_05100_, _05099_, _04544_);
  and _56561_ (_05101_, _05100_, _05098_);
  nor _56562_ (_05102_, _05101_, _04966_);
  nor _56563_ (_05103_, _05102_, _04795_);
  not _56564_ (_05104_, _05103_);
  nor _56565_ (_05105_, _05104_, _04964_);
  and _56566_ (_05106_, _05105_, _04797_);
  or _56567_ (_05107_, _05106_, \oc8051_golden_model_1.IRAM[15] [7]);
  and _56568_ (_05108_, _04848_, _03502_);
  nor _56569_ (_05109_, _04970_, _04551_);
  nor _56570_ (_05110_, _05109_, _05108_);
  and _56571_ (_05111_, _04849_, _03502_);
  nor _56572_ (_05112_, _05108_, _04851_);
  nor _56573_ (_05113_, _05112_, _05111_);
  and _56574_ (_05114_, _04533_, _04755_);
  and _56575_ (_05115_, _05114_, _04748_);
  and _56576_ (_05116_, _05115_, _04762_);
  nor _56577_ (_05117_, _05116_, _04701_);
  and _56578_ (_05118_, _05117_, _05113_);
  and _56579_ (_05119_, _05118_, _05110_);
  and _56580_ (_05120_, _05119_, _04550_);
  not _56581_ (_05121_, _05120_);
  and _56582_ (_05122_, _05121_, _05107_);
  not _56583_ (_05123_, _05106_);
  not _56584_ (_05124_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _56585_ (_05125_, _04373_, _05124_);
  not _56586_ (_05126_, \oc8051_golden_model_1.IRAM[1] [7]);
  or _56587_ (_05127_, _04217_, _05126_);
  and _56588_ (_05128_, _05127_, _04368_);
  nand _56589_ (_05129_, _05128_, _05125_);
  not _56590_ (_05130_, \oc8051_golden_model_1.IRAM[3] [7]);
  or _56591_ (_05131_, _04217_, _05130_);
  not _56592_ (_05132_, \oc8051_golden_model_1.IRAM[2] [7]);
  or _56593_ (_05133_, _04373_, _05132_);
  and _56594_ (_05134_, _05133_, _04375_);
  nand _56595_ (_05135_, _05134_, _05131_);
  nand _56596_ (_05136_, _05135_, _05129_);
  nand _56597_ (_05137_, _05136_, _03994_);
  not _56598_ (_05138_, \oc8051_golden_model_1.IRAM[7] [7]);
  or _56599_ (_05139_, _04217_, _05138_);
  not _56600_ (_05140_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _56601_ (_05141_, _04373_, _05140_);
  and _56602_ (_05142_, _05141_, _04375_);
  nand _56603_ (_05143_, _05142_, _05139_);
  not _56604_ (_05144_, \oc8051_golden_model_1.IRAM[4] [7]);
  or _56605_ (_05145_, _04373_, _05144_);
  not _56606_ (_05146_, \oc8051_golden_model_1.IRAM[5] [7]);
  or _56607_ (_05147_, _04217_, _05146_);
  and _56608_ (_05148_, _05147_, _04368_);
  nand _56609_ (_05149_, _05148_, _05145_);
  nand _56610_ (_05150_, _05149_, _05143_);
  nand _56611_ (_05151_, _05150_, _04382_);
  nand _56612_ (_05152_, _05151_, _05137_);
  nand _56613_ (_05153_, _05152_, _03803_);
  nand _56614_ (_05154_, _04373_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand _56615_ (_05155_, _04217_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _56616_ (_05156_, _05155_, _04375_);
  nand _56617_ (_05157_, _05156_, _05154_);
  nand _56618_ (_05158_, _04217_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand _56619_ (_05159_, _04373_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _56620_ (_05160_, _05159_, _04368_);
  nand _56621_ (_05161_, _05160_, _05158_);
  nand _56622_ (_05162_, _05161_, _05157_);
  nand _56623_ (_05163_, _05162_, _03994_);
  nand _56624_ (_05164_, _04373_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand _56625_ (_05165_, _04217_, \oc8051_golden_model_1.IRAM[14] [7]);
  and _56626_ (_05166_, _05165_, _04375_);
  nand _56627_ (_05167_, _05166_, _05164_);
  nand _56628_ (_05168_, _04217_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand _56629_ (_05169_, _04373_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _56630_ (_05170_, _05169_, _04368_);
  nand _56631_ (_05171_, _05170_, _05168_);
  nand _56632_ (_05172_, _05171_, _05167_);
  nand _56633_ (_05173_, _05172_, _04382_);
  nand _56634_ (_05174_, _05173_, _05163_);
  nand _56635_ (_05175_, _05174_, _04396_);
  nand _56636_ (_05176_, _05175_, _05153_);
  or _56637_ (_05177_, _05176_, _03401_);
  and _56638_ (_05178_, _04284_, _03472_);
  and _56639_ (_05179_, _05178_, _03877_);
  and _56640_ (_05180_, _05179_, _03563_);
  and _56641_ (_05181_, _03561_, _03401_);
  not _56642_ (_05182_, _04249_);
  and _56643_ (_05183_, _05182_, _03834_);
  and _56644_ (_05184_, _05183_, _05181_);
  and _56645_ (_05185_, _05184_, _05180_);
  and _56646_ (_05186_, _05185_, \oc8051_golden_model_1.SBUF [7]);
  and _56647_ (_05187_, _04284_, _03471_);
  and _56648_ (_05188_, _05187_, _03877_);
  and _56649_ (_05189_, _05188_, _03563_);
  not _56650_ (_05190_, _03834_);
  and _56651_ (_05191_, _04249_, _05190_);
  and _56652_ (_05192_, _05191_, _05181_);
  and _56653_ (_05193_, _05192_, _05189_);
  and _56654_ (_05194_, _05193_, \oc8051_golden_model_1.IE [7]);
  nor _56655_ (_05195_, _05194_, _05186_);
  and _56656_ (_05196_, _03877_, _03432_);
  and _56657_ (_05197_, _05187_, _05196_);
  nor _56658_ (_05198_, _04249_, _03834_);
  and _56659_ (_05199_, _05198_, _05181_);
  and _56660_ (_05200_, _05199_, _05197_);
  and _56661_ (_05201_, _05200_, \oc8051_golden_model_1.P3 [7]);
  not _56662_ (_05202_, _05201_);
  and _56663_ (_05203_, _05181_, _03834_);
  and _56664_ (_05204_, _05203_, _04249_);
  and _56665_ (_05205_, _05204_, _03432_);
  nor _56666_ (_05206_, _04284_, _03471_);
  and _56667_ (_05207_, _05206_, _04965_);
  and _56668_ (_05208_, _05207_, _05205_);
  and _56669_ (_05209_, _05208_, \oc8051_golden_model_1.PCON [7]);
  and _56670_ (_05210_, _05197_, _05192_);
  and _56671_ (_05211_, _05210_, \oc8051_golden_model_1.P2 [7]);
  nor _56672_ (_05212_, _05211_, _05209_);
  and _56673_ (_05213_, _05212_, _05202_);
  and _56674_ (_05214_, _05213_, _05195_);
  not _56675_ (_05215_, _03401_);
  nor _56676_ (_05216_, _03561_, _05215_);
  and _56677_ (_05217_, _05216_, _05183_);
  and _56678_ (_05218_, _05217_, _05197_);
  and _56679_ (_05219_, _05218_, \oc8051_golden_model_1.PSW [7]);
  and _56680_ (_05220_, _05198_, _05216_);
  and _56681_ (_05221_, _05220_, _05197_);
  and _56682_ (_05222_, _05221_, \oc8051_golden_model_1.B [7]);
  nor _56683_ (_05223_, _05222_, _05219_);
  and _56684_ (_05224_, _05199_, _05189_);
  and _56685_ (_05225_, _05224_, \oc8051_golden_model_1.IP [7]);
  and _56686_ (_05226_, _05216_, _05191_);
  and _56687_ (_05227_, _05226_, _05197_);
  and _56688_ (_05228_, _05227_, \oc8051_golden_model_1.ACC [7]);
  nor _56689_ (_05229_, _05228_, _05225_);
  and _56690_ (_05230_, _05229_, _05223_);
  not _56691_ (_05231_, _05204_);
  nor _56692_ (_05232_, _03877_, _03432_);
  nand _56693_ (_05233_, _05232_, _05187_);
  nor _56694_ (_05234_, _05233_, _05231_);
  and _56695_ (_05235_, _05234_, \oc8051_golden_model_1.TH0 [7]);
  and _56696_ (_05236_, _05189_, _05204_);
  and _56697_ (_05237_, _05236_, \oc8051_golden_model_1.TCON [7]);
  nor _56698_ (_05238_, _05237_, _05235_);
  not _56699_ (_05239_, _05206_);
  nand _56700_ (_05240_, _03877_, _03563_);
  or _56701_ (_05241_, _05240_, _05239_);
  nor _56702_ (_05242_, _05241_, _05231_);
  and _56703_ (_05243_, _05242_, \oc8051_golden_model_1.TL1 [7]);
  and _56704_ (_05244_, _05197_, _05184_);
  and _56705_ (_05245_, _05244_, \oc8051_golden_model_1.P1 [7]);
  nor _56706_ (_05246_, _05245_, _05243_);
  and _56707_ (_05247_, _05246_, _05238_);
  and _56708_ (_05248_, _05184_, _05189_);
  and _56709_ (_05249_, _05248_, \oc8051_golden_model_1.SCON [7]);
  nand _56710_ (_05250_, _05232_, _05178_);
  nor _56711_ (_05251_, _05250_, _05231_);
  and _56712_ (_05252_, _05251_, \oc8051_golden_model_1.TH1 [7]);
  nor _56713_ (_05253_, _05252_, _05249_);
  and _56714_ (_05254_, _05180_, _05204_);
  and _56715_ (_05255_, _05254_, \oc8051_golden_model_1.TMOD [7]);
  nor _56716_ (_05256_, _04284_, _03472_);
  nor _56717_ (_05257_, _05240_, _05231_);
  and _56718_ (_05258_, _05257_, _05256_);
  and _56719_ (_05259_, _05258_, \oc8051_golden_model_1.TL0 [7]);
  nor _56720_ (_05260_, _05259_, _05255_);
  and _56721_ (_05261_, _05260_, _05253_);
  and _56722_ (_05262_, _05261_, _05247_);
  and _56723_ (_05263_, _05262_, _05230_);
  and _56724_ (_05264_, _05263_, _05214_);
  and _56725_ (_05265_, _05206_, _03877_);
  and _56726_ (_05266_, _05265_, _05205_);
  and _56727_ (_05267_, _05266_, \oc8051_golden_model_1.DPH [7]);
  not _56728_ (_05268_, _05267_);
  and _56729_ (_05269_, _05179_, _05205_);
  and _56730_ (_05270_, _05269_, \oc8051_golden_model_1.SP [7]);
  and _56731_ (_05271_, _05256_, _03877_);
  and _56732_ (_05272_, _05271_, _05205_);
  and _56733_ (_05273_, _05272_, \oc8051_golden_model_1.DPL [7]);
  nor _56734_ (_05274_, _05273_, _05270_);
  and _56735_ (_05275_, _05274_, _05268_);
  and _56736_ (_05276_, _05197_, _05204_);
  and _56737_ (_05277_, _05276_, \oc8051_golden_model_1.P0 [7]);
  not _56738_ (_05278_, _05277_);
  and _56739_ (_05279_, _05278_, _05275_);
  and _56740_ (_05280_, _05279_, _05264_);
  and _56741_ (_05281_, _05280_, _05177_);
  not _56742_ (_05282_, _05281_);
  nand _56743_ (_05283_, _04217_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand _56744_ (_05284_, _04373_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _56745_ (_05285_, _05284_, _04368_);
  nand _56746_ (_05286_, _05285_, _05283_);
  nand _56747_ (_05287_, _04373_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand _56748_ (_05288_, _04217_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _56749_ (_05289_, _05288_, _04375_);
  nand _56750_ (_05290_, _05289_, _05287_);
  nand _56751_ (_05291_, _05290_, _05286_);
  nand _56752_ (_05292_, _05291_, _03994_);
  nand _56753_ (_05293_, _04373_, \oc8051_golden_model_1.IRAM[7] [6]);
  nand _56754_ (_05294_, _04217_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _56755_ (_05295_, _05294_, _04375_);
  nand _56756_ (_05296_, _05295_, _05293_);
  nand _56757_ (_05297_, _04217_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand _56758_ (_05298_, _04373_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _56759_ (_05299_, _05298_, _04368_);
  nand _56760_ (_05300_, _05299_, _05297_);
  nand _56761_ (_05301_, _05300_, _05296_);
  nand _56762_ (_05302_, _05301_, _04382_);
  nand _56763_ (_05303_, _05302_, _05292_);
  nand _56764_ (_05304_, _05303_, _03803_);
  nand _56765_ (_05305_, _04373_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _56766_ (_05306_, _04217_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _56767_ (_05307_, _05306_, _04375_);
  nand _56768_ (_05308_, _05307_, _05305_);
  nand _56769_ (_05309_, _04217_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand _56770_ (_05310_, _04373_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _56771_ (_05311_, _05310_, _04368_);
  nand _56772_ (_05312_, _05311_, _05309_);
  nand _56773_ (_05313_, _05312_, _05308_);
  nand _56774_ (_05314_, _05313_, _03994_);
  nand _56775_ (_05315_, _04373_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _56776_ (_05316_, _04217_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _56777_ (_05317_, _05316_, _04375_);
  nand _56778_ (_05318_, _05317_, _05315_);
  nand _56779_ (_05319_, _04217_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand _56780_ (_05320_, _04373_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _56781_ (_05321_, _05320_, _04368_);
  nand _56782_ (_05322_, _05321_, _05319_);
  nand _56783_ (_05323_, _05322_, _05318_);
  nand _56784_ (_05324_, _05323_, _04382_);
  nand _56785_ (_05325_, _05324_, _05314_);
  nand _56786_ (_05326_, _05325_, _04396_);
  nand _56787_ (_05327_, _05326_, _05304_);
  or _56788_ (_05328_, _05327_, _03401_);
  and _56789_ (_05329_, _05266_, \oc8051_golden_model_1.DPH [6]);
  not _56790_ (_05330_, _05329_);
  and _56791_ (_05331_, _05269_, \oc8051_golden_model_1.SP [6]);
  and _56792_ (_05332_, _05258_, \oc8051_golden_model_1.TL0 [6]);
  nor _56793_ (_05333_, _05332_, _05331_);
  and _56794_ (_05334_, _05333_, _05330_);
  and _56795_ (_05335_, _05248_, \oc8051_golden_model_1.SCON [6]);
  not _56796_ (_05336_, _05335_);
  and _56797_ (_05337_, _05251_, \oc8051_golden_model_1.TH1 [6]);
  and _56798_ (_05338_, _05185_, \oc8051_golden_model_1.SBUF [6]);
  nor _56799_ (_05339_, _05338_, _05337_);
  and _56800_ (_05340_, _05339_, _05336_);
  and _56801_ (_05341_, _05272_, \oc8051_golden_model_1.DPL [6]);
  not _56802_ (_05342_, _05341_);
  and _56803_ (_05343_, _05254_, \oc8051_golden_model_1.TMOD [6]);
  and _56804_ (_05344_, _05193_, \oc8051_golden_model_1.IE [6]);
  nor _56805_ (_05345_, _05344_, _05343_);
  and _56806_ (_05346_, _05345_, _05342_);
  and _56807_ (_05347_, _05346_, _05340_);
  and _56808_ (_05348_, _05347_, _05334_);
  not _56809_ (_05349_, _05348_);
  and _56810_ (_05350_, _05208_, \oc8051_golden_model_1.PCON [6]);
  and _56811_ (_05351_, _05276_, \oc8051_golden_model_1.P0 [6]);
  not _56812_ (_05352_, _05351_);
  and _56813_ (_05353_, _05224_, \oc8051_golden_model_1.IP [6]);
  and _56814_ (_05354_, _05227_, \oc8051_golden_model_1.ACC [6]);
  nor _56815_ (_05355_, _05354_, _05353_);
  and _56816_ (_05356_, _05218_, \oc8051_golden_model_1.PSW [6]);
  and _56817_ (_05357_, _05221_, \oc8051_golden_model_1.B [6]);
  nor _56818_ (_05358_, _05357_, _05356_);
  and _56819_ (_05359_, _05358_, _05355_);
  nand _56820_ (_05360_, _05359_, _05352_);
  or _56821_ (_05361_, _05360_, _05350_);
  and _56822_ (_05362_, _05234_, \oc8051_golden_model_1.TH0 [6]);
  and _56823_ (_05363_, _05242_, \oc8051_golden_model_1.TL1 [6]);
  nor _56824_ (_05364_, _05363_, _05362_);
  and _56825_ (_05365_, _05236_, \oc8051_golden_model_1.TCON [6]);
  not _56826_ (_05366_, _05365_);
  and _56827_ (_05367_, _05244_, \oc8051_golden_model_1.P1 [6]);
  and _56828_ (_05368_, _05210_, \oc8051_golden_model_1.P2 [6]);
  and _56829_ (_05369_, _05200_, \oc8051_golden_model_1.P3 [6]);
  or _56830_ (_05370_, _05369_, _05368_);
  nor _56831_ (_05371_, _05370_, _05367_);
  and _56832_ (_05372_, _05371_, _05366_);
  nand _56833_ (_05373_, _05372_, _05364_);
  or _56834_ (_05374_, _05373_, _05361_);
  nor _56835_ (_05375_, _05374_, _05349_);
  and _56836_ (_05376_, _05375_, _05328_);
  not _56837_ (_05377_, _05376_);
  nand _56838_ (_05378_, _04217_, \oc8051_golden_model_1.IRAM[0] [5]);
  nand _56839_ (_05379_, _04373_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _56840_ (_05380_, _05379_, _04368_);
  nand _56841_ (_05381_, _05380_, _05378_);
  nand _56842_ (_05382_, _04373_, \oc8051_golden_model_1.IRAM[3] [5]);
  nand _56843_ (_05383_, _04217_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _56844_ (_05384_, _05383_, _04375_);
  nand _56845_ (_05385_, _05384_, _05382_);
  nand _56846_ (_05386_, _05385_, _05381_);
  nand _56847_ (_05387_, _05386_, _03994_);
  nand _56848_ (_05388_, _04373_, \oc8051_golden_model_1.IRAM[7] [5]);
  nand _56849_ (_05389_, _04217_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _56850_ (_05390_, _05389_, _04375_);
  nand _56851_ (_05391_, _05390_, _05388_);
  nand _56852_ (_05392_, _04217_, \oc8051_golden_model_1.IRAM[4] [5]);
  nand _56853_ (_05393_, _04373_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _56854_ (_05394_, _05393_, _04368_);
  nand _56855_ (_05395_, _05394_, _05392_);
  nand _56856_ (_05396_, _05395_, _05391_);
  nand _56857_ (_05397_, _05396_, _04382_);
  nand _56858_ (_05398_, _05397_, _05387_);
  nand _56859_ (_05399_, _05398_, _03803_);
  nand _56860_ (_05400_, _04373_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _56861_ (_05401_, _04217_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _56862_ (_05402_, _05401_, _04375_);
  nand _56863_ (_05403_, _05402_, _05400_);
  nand _56864_ (_05404_, _04217_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand _56865_ (_05405_, _04373_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _56866_ (_05406_, _05405_, _04368_);
  nand _56867_ (_05407_, _05406_, _05404_);
  nand _56868_ (_05408_, _05407_, _05403_);
  nand _56869_ (_05409_, _05408_, _03994_);
  nand _56870_ (_05410_, _04373_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _56871_ (_05411_, _04217_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _56872_ (_05412_, _05411_, _04375_);
  nand _56873_ (_05413_, _05412_, _05410_);
  nand _56874_ (_05414_, _04217_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand _56875_ (_05415_, _04373_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _56876_ (_05416_, _05415_, _04368_);
  nand _56877_ (_05417_, _05416_, _05414_);
  nand _56878_ (_05418_, _05417_, _05413_);
  nand _56879_ (_05419_, _05418_, _04382_);
  nand _56880_ (_05420_, _05419_, _05409_);
  nand _56881_ (_05421_, _05420_, _04396_);
  nand _56882_ (_05422_, _05421_, _05399_);
  or _56883_ (_05423_, _05422_, _03401_);
  and _56884_ (_05424_, _05272_, \oc8051_golden_model_1.DPL [5]);
  not _56885_ (_05425_, _05424_);
  and _56886_ (_05426_, _05266_, \oc8051_golden_model_1.DPH [5]);
  and _56887_ (_05427_, _05258_, \oc8051_golden_model_1.TL0 [5]);
  nor _56888_ (_05428_, _05427_, _05426_);
  and _56889_ (_05429_, _05428_, _05425_);
  and _56890_ (_05430_, _05236_, \oc8051_golden_model_1.TCON [5]);
  not _56891_ (_05431_, _05430_);
  and _56892_ (_05432_, _05251_, \oc8051_golden_model_1.TH1 [5]);
  and _56893_ (_05433_, _05248_, \oc8051_golden_model_1.SCON [5]);
  nor _56894_ (_05434_, _05433_, _05432_);
  and _56895_ (_05435_, _05434_, _05431_);
  and _56896_ (_05436_, _05254_, \oc8051_golden_model_1.TMOD [5]);
  and _56897_ (_05437_, _05193_, \oc8051_golden_model_1.IE [5]);
  nor _56898_ (_05438_, _05437_, _05436_);
  and _56899_ (_05439_, _05234_, \oc8051_golden_model_1.TH0 [5]);
  and _56900_ (_05440_, _05185_, \oc8051_golden_model_1.SBUF [5]);
  nor _56901_ (_05441_, _05440_, _05439_);
  and _56902_ (_05442_, _05441_, _05438_);
  and _56903_ (_05443_, _05269_, \oc8051_golden_model_1.SP [5]);
  and _56904_ (_05444_, _05257_, _05206_);
  and _56905_ (_05445_, _05444_, \oc8051_golden_model_1.TL1 [5]);
  nor _56906_ (_05446_, _05445_, _05443_);
  and _56907_ (_05447_, _05446_, _05442_);
  and _56908_ (_05448_, _05447_, _05435_);
  and _56909_ (_05449_, _05448_, _05429_);
  and _56910_ (_05450_, _05208_, \oc8051_golden_model_1.PCON [5]);
  not _56911_ (_05451_, _05450_);
  and _56912_ (_05452_, _05218_, \oc8051_golden_model_1.PSW [5]);
  and _56913_ (_05453_, _05227_, \oc8051_golden_model_1.ACC [5]);
  nor _56914_ (_05454_, _05453_, _05452_);
  and _56915_ (_05455_, _05224_, \oc8051_golden_model_1.IP [5]);
  and _56916_ (_05456_, _05221_, \oc8051_golden_model_1.B [5]);
  nor _56917_ (_05457_, _05456_, _05455_);
  and _56918_ (_05458_, _05457_, _05454_);
  and _56919_ (_05459_, _05458_, _05451_);
  and _56920_ (_05460_, _05276_, \oc8051_golden_model_1.P0 [5]);
  not _56921_ (_05461_, _05460_);
  and _56922_ (_05462_, _05244_, \oc8051_golden_model_1.P1 [5]);
  not _56923_ (_05463_, _05462_);
  and _56924_ (_05464_, _05210_, \oc8051_golden_model_1.P2 [5]);
  and _56925_ (_05465_, _05200_, \oc8051_golden_model_1.P3 [5]);
  nor _56926_ (_05466_, _05465_, _05464_);
  and _56927_ (_05467_, _05466_, _05463_);
  and _56928_ (_05468_, _05467_, _05461_);
  and _56929_ (_05469_, _05468_, _05459_);
  and _56930_ (_05470_, _05469_, _05449_);
  and _56931_ (_05471_, _05470_, _05423_);
  not _56932_ (_05472_, _05471_);
  or _56933_ (_05473_, _04843_, _03401_);
  and _56934_ (_05474_, _05208_, \oc8051_golden_model_1.PCON [3]);
  not _56935_ (_05475_, _05474_);
  and _56936_ (_05476_, _05185_, \oc8051_golden_model_1.SBUF [3]);
  and _56937_ (_05477_, _05193_, \oc8051_golden_model_1.IE [3]);
  nor _56938_ (_05478_, _05477_, _05476_);
  and _56939_ (_05479_, _05478_, _05475_);
  and _56940_ (_05480_, _05210_, \oc8051_golden_model_1.P2 [3]);
  and _56941_ (_05481_, _05200_, \oc8051_golden_model_1.P3 [3]);
  nor _56942_ (_05482_, _05481_, _05480_);
  and _56943_ (_05483_, _05482_, _05479_);
  and _56944_ (_05484_, _05218_, \oc8051_golden_model_1.PSW [3]);
  not _56945_ (_05485_, _05484_);
  and _56946_ (_05486_, _05224_, \oc8051_golden_model_1.IP [3]);
  not _56947_ (_05487_, _05486_);
  and _56948_ (_05488_, _05227_, \oc8051_golden_model_1.ACC [3]);
  and _56949_ (_05489_, _05221_, \oc8051_golden_model_1.B [3]);
  nor _56950_ (_05490_, _05489_, _05488_);
  and _56951_ (_05491_, _05490_, _05487_);
  and _56952_ (_05492_, _05491_, _05485_);
  and _56953_ (_05493_, _05236_, \oc8051_golden_model_1.TCON [3]);
  and _56954_ (_05494_, _05234_, \oc8051_golden_model_1.TH0 [3]);
  nor _56955_ (_05495_, _05494_, _05493_);
  and _56956_ (_05496_, _05244_, \oc8051_golden_model_1.P1 [3]);
  and _56957_ (_05497_, _05242_, \oc8051_golden_model_1.TL1 [3]);
  nor _56958_ (_05498_, _05497_, _05496_);
  and _56959_ (_05499_, _05498_, _05495_);
  and _56960_ (_05500_, _05248_, \oc8051_golden_model_1.SCON [3]);
  and _56961_ (_05501_, _05251_, \oc8051_golden_model_1.TH1 [3]);
  nor _56962_ (_05502_, _05501_, _05500_);
  and _56963_ (_05503_, _05254_, \oc8051_golden_model_1.TMOD [3]);
  and _56964_ (_05504_, _05258_, \oc8051_golden_model_1.TL0 [3]);
  nor _56965_ (_05505_, _05504_, _05503_);
  and _56966_ (_05506_, _05505_, _05502_);
  and _56967_ (_05507_, _05506_, _05499_);
  and _56968_ (_05508_, _05507_, _05492_);
  and _56969_ (_05509_, _05508_, _05483_);
  and _56970_ (_05510_, _05276_, \oc8051_golden_model_1.P0 [3]);
  not _56971_ (_05511_, _05510_);
  and _56972_ (_05512_, _05266_, \oc8051_golden_model_1.DPH [3]);
  not _56973_ (_05513_, _05512_);
  and _56974_ (_05514_, _05269_, \oc8051_golden_model_1.SP [3]);
  and _56975_ (_05515_, _05272_, \oc8051_golden_model_1.DPL [3]);
  nor _56976_ (_05516_, _05515_, _05514_);
  and _56977_ (_05517_, _05516_, _05513_);
  and _56978_ (_05518_, _05517_, _05511_);
  and _56979_ (_05519_, _05518_, _05509_);
  and _56980_ (_05520_, _05519_, _05473_);
  not _56981_ (_05521_, _05520_);
  or _56982_ (_05522_, _04603_, _03401_);
  and _56983_ (_05523_, _05266_, \oc8051_golden_model_1.DPH [1]);
  not _56984_ (_05524_, _05523_);
  and _56985_ (_05525_, _05269_, \oc8051_golden_model_1.SP [1]);
  and _56986_ (_05526_, _05272_, \oc8051_golden_model_1.DPL [1]);
  nor _56987_ (_05527_, _05526_, _05525_);
  and _56988_ (_05528_, _05527_, _05524_);
  and _56989_ (_05529_, _05254_, \oc8051_golden_model_1.TMOD [1]);
  not _56990_ (_05530_, _05529_);
  and _56991_ (_05531_, _05248_, \oc8051_golden_model_1.SCON [1]);
  and _56992_ (_05532_, _05185_, \oc8051_golden_model_1.SBUF [1]);
  nor _56993_ (_05533_, _05532_, _05531_);
  and _56994_ (_05534_, _05533_, _05530_);
  and _56995_ (_05535_, _05258_, \oc8051_golden_model_1.TL0 [1]);
  not _56996_ (_05536_, _05535_);
  and _56997_ (_05537_, _05251_, \oc8051_golden_model_1.TH1 [1]);
  and _56998_ (_05538_, _05193_, \oc8051_golden_model_1.IE [1]);
  nor _56999_ (_05539_, _05538_, _05537_);
  and _57000_ (_05540_, _05539_, _05536_);
  and _57001_ (_05541_, _05540_, _05534_);
  and _57002_ (_05542_, _05541_, _05528_);
  and _57003_ (_05543_, _05236_, \oc8051_golden_model_1.TCON [1]);
  and _57004_ (_05544_, _05234_, \oc8051_golden_model_1.TH0 [1]);
  nor _57005_ (_05545_, _05544_, _05543_);
  and _57006_ (_05546_, _05444_, \oc8051_golden_model_1.TL1 [1]);
  not _57007_ (_05547_, _05546_);
  and _57008_ (_05548_, _05547_, _05545_);
  and _57009_ (_05549_, _05224_, \oc8051_golden_model_1.IP [1]);
  and _57010_ (_05550_, _05227_, \oc8051_golden_model_1.ACC [1]);
  nor _57011_ (_05551_, _05550_, _05549_);
  and _57012_ (_05552_, _05218_, \oc8051_golden_model_1.PSW [1]);
  and _57013_ (_05553_, _05221_, \oc8051_golden_model_1.B [1]);
  nor _57014_ (_05554_, _05553_, _05552_);
  and _57015_ (_05555_, _05554_, _05551_);
  and _57016_ (_05556_, _05244_, \oc8051_golden_model_1.P1 [1]);
  not _57017_ (_05557_, _05556_);
  and _57018_ (_05558_, _05210_, \oc8051_golden_model_1.P2 [1]);
  and _57019_ (_05559_, _05200_, \oc8051_golden_model_1.P3 [1]);
  nor _57020_ (_05560_, _05559_, _05558_);
  and _57021_ (_05561_, _05560_, _05557_);
  and _57022_ (_05562_, _05561_, _05555_);
  and _57023_ (_05563_, _05276_, \oc8051_golden_model_1.P0 [1]);
  and _57024_ (_05564_, _05208_, \oc8051_golden_model_1.PCON [1]);
  nor _57025_ (_05565_, _05564_, _05563_);
  and _57026_ (_05566_, _05565_, _05562_);
  and _57027_ (_05567_, _05566_, _05548_);
  and _57028_ (_05568_, _05567_, _05542_);
  nand _57029_ (_05569_, _05568_, _05522_);
  or _57030_ (_05570_, _04439_, _03401_);
  and _57031_ (_05571_, _05224_, \oc8051_golden_model_1.IP [0]);
  and _57032_ (_05572_, _05221_, \oc8051_golden_model_1.B [0]);
  nor _57033_ (_05573_, _05572_, _05571_);
  and _57034_ (_05574_, _05218_, \oc8051_golden_model_1.PSW [0]);
  and _57035_ (_05575_, _05227_, \oc8051_golden_model_1.ACC [0]);
  nor _57036_ (_05576_, _05575_, _05574_);
  and _57037_ (_05577_, _05576_, _05573_);
  and _57038_ (_05578_, _05276_, \oc8051_golden_model_1.P0 [0]);
  not _57039_ (_05579_, _05578_);
  and _57040_ (_05580_, _05244_, \oc8051_golden_model_1.P1 [0]);
  not _57041_ (_05581_, _05580_);
  and _57042_ (_05582_, _05210_, \oc8051_golden_model_1.P2 [0]);
  and _57043_ (_05583_, _05200_, \oc8051_golden_model_1.P3 [0]);
  nor _57044_ (_05584_, _05583_, _05582_);
  and _57045_ (_05585_, _05584_, _05581_);
  and _57046_ (_05586_, _05585_, _05579_);
  and _57047_ (_05587_, _05586_, _05577_);
  and _57048_ (_05588_, _05269_, \oc8051_golden_model_1.SP [0]);
  and _57049_ (_05589_, _05272_, \oc8051_golden_model_1.DPL [0]);
  nor _57050_ (_05590_, _05589_, _05588_);
  and _57051_ (_05591_, _05208_, \oc8051_golden_model_1.PCON [0]);
  not _57052_ (_05592_, _05591_);
  and _57053_ (_05593_, _05185_, \oc8051_golden_model_1.SBUF [0]);
  and _57054_ (_05594_, _05193_, \oc8051_golden_model_1.IE [0]);
  nor _57055_ (_05595_, _05594_, _05593_);
  and _57056_ (_05596_, _05595_, _05592_);
  and _57057_ (_05597_, _05596_, _05590_);
  and _57058_ (_05598_, _05597_, _05587_);
  and _57059_ (_05599_, _05258_, \oc8051_golden_model_1.TL0 [0]);
  not _57060_ (_05600_, _05599_);
  and _57061_ (_05601_, _05254_, \oc8051_golden_model_1.TMOD [0]);
  and _57062_ (_05602_, _05248_, \oc8051_golden_model_1.SCON [0]);
  nor _57063_ (_05603_, _05602_, _05601_);
  and _57064_ (_05604_, _05236_, \oc8051_golden_model_1.TCON [0]);
  and _57065_ (_05605_, _05251_, \oc8051_golden_model_1.TH1 [0]);
  nor _57066_ (_05606_, _05605_, _05604_);
  and _57067_ (_05607_, _05606_, _05603_);
  and _57068_ (_05608_, _05607_, _05600_);
  and _57069_ (_05609_, _05444_, \oc8051_golden_model_1.TL1 [0]);
  not _57070_ (_05610_, _05609_);
  and _57071_ (_05611_, _05266_, \oc8051_golden_model_1.DPH [0]);
  and _57072_ (_05612_, _05234_, \oc8051_golden_model_1.TH0 [0]);
  nor _57073_ (_05613_, _05612_, _05611_);
  and _57074_ (_05614_, _05613_, _05610_);
  and _57075_ (_05615_, _05614_, _05608_);
  and _57076_ (_05616_, _05615_, _05598_);
  nand _57077_ (_05617_, _05616_, _05570_);
  and _57078_ (_05618_, _05617_, _05569_);
  or _57079_ (_05619_, _05026_, _03401_);
  and _57080_ (_05620_, _05269_, \oc8051_golden_model_1.SP [2]);
  and _57081_ (_05621_, _05272_, \oc8051_golden_model_1.DPL [2]);
  nor _57082_ (_05622_, _05621_, _05620_);
  and _57083_ (_05623_, _05236_, \oc8051_golden_model_1.TCON [2]);
  and _57084_ (_05624_, _05234_, \oc8051_golden_model_1.TH0 [2]);
  nor _57085_ (_05625_, _05624_, _05623_);
  and _57086_ (_05626_, _05244_, \oc8051_golden_model_1.P1 [2]);
  and _57087_ (_05627_, _05242_, \oc8051_golden_model_1.TL1 [2]);
  nor _57088_ (_05628_, _05627_, _05626_);
  and _57089_ (_05629_, _05628_, _05625_);
  and _57090_ (_05630_, _05248_, \oc8051_golden_model_1.SCON [2]);
  and _57091_ (_05631_, _05251_, \oc8051_golden_model_1.TH1 [2]);
  nor _57092_ (_05632_, _05631_, _05630_);
  and _57093_ (_05633_, _05258_, \oc8051_golden_model_1.TL0 [2]);
  and _57094_ (_05634_, _05254_, \oc8051_golden_model_1.TMOD [2]);
  nor _57095_ (_05635_, _05634_, _05633_);
  and _57096_ (_05636_, _05635_, _05632_);
  and _57097_ (_05637_, _05636_, _05629_);
  and _57098_ (_05638_, _05637_, _05622_);
  and _57099_ (_05639_, _05210_, \oc8051_golden_model_1.P2 [2]);
  and _57100_ (_05640_, _05200_, \oc8051_golden_model_1.P3 [2]);
  nor _57101_ (_05641_, _05640_, _05639_);
  and _57102_ (_05642_, _05208_, \oc8051_golden_model_1.PCON [2]);
  not _57103_ (_05643_, _05642_);
  and _57104_ (_05644_, _05185_, \oc8051_golden_model_1.SBUF [2]);
  and _57105_ (_05645_, _05193_, \oc8051_golden_model_1.IE [2]);
  nor _57106_ (_05646_, _05645_, _05644_);
  and _57107_ (_05647_, _05646_, _05643_);
  and _57108_ (_05648_, _05647_, _05641_);
  and _57109_ (_05649_, _05224_, \oc8051_golden_model_1.IP [2]);
  not _57110_ (_05650_, _05649_);
  and _57111_ (_05651_, _05218_, \oc8051_golden_model_1.PSW [2]);
  not _57112_ (_05652_, _05651_);
  and _57113_ (_05653_, _05227_, \oc8051_golden_model_1.ACC [2]);
  and _57114_ (_05654_, _05221_, \oc8051_golden_model_1.B [2]);
  nor _57115_ (_05655_, _05654_, _05653_);
  and _57116_ (_05656_, _05655_, _05652_);
  and _57117_ (_05657_, _05656_, _05650_);
  and _57118_ (_05658_, _05276_, \oc8051_golden_model_1.P0 [2]);
  and _57119_ (_05659_, _05266_, \oc8051_golden_model_1.DPH [2]);
  nor _57120_ (_05660_, _05659_, _05658_);
  and _57121_ (_05661_, _05660_, _05657_);
  and _57122_ (_05662_, _05661_, _05648_);
  and _57123_ (_05663_, _05662_, _05638_);
  and _57124_ (_05664_, _05663_, _05619_);
  not _57125_ (_05665_, _05664_);
  and _57126_ (_05666_, _05665_, _05618_);
  and _57127_ (_05667_, _05666_, _05521_);
  nand _57128_ (_05668_, _04217_, \oc8051_golden_model_1.IRAM[0] [4]);
  nand _57129_ (_05669_, _04373_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _57130_ (_05670_, _05669_, _04368_);
  nand _57131_ (_05671_, _05670_, _05668_);
  nand _57132_ (_05672_, _04373_, \oc8051_golden_model_1.IRAM[3] [4]);
  nand _57133_ (_05673_, _04217_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _57134_ (_05674_, _05673_, _04375_);
  nand _57135_ (_05675_, _05674_, _05672_);
  nand _57136_ (_05676_, _05675_, _05671_);
  nand _57137_ (_05677_, _05676_, _03994_);
  nand _57138_ (_05678_, _04373_, \oc8051_golden_model_1.IRAM[7] [4]);
  nand _57139_ (_05679_, _04217_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _57140_ (_05680_, _05679_, _04375_);
  nand _57141_ (_05681_, _05680_, _05678_);
  nand _57142_ (_05682_, _04217_, \oc8051_golden_model_1.IRAM[4] [4]);
  nand _57143_ (_05683_, _04373_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _57144_ (_05684_, _05683_, _04368_);
  nand _57145_ (_05685_, _05684_, _05682_);
  nand _57146_ (_05686_, _05685_, _05681_);
  nand _57147_ (_05687_, _05686_, _04382_);
  nand _57148_ (_05688_, _05687_, _05677_);
  nand _57149_ (_05689_, _05688_, _03803_);
  nand _57150_ (_05690_, _04373_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _57151_ (_05691_, _04217_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _57152_ (_05692_, _05691_, _04375_);
  nand _57153_ (_05693_, _05692_, _05690_);
  nand _57154_ (_05694_, _04217_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand _57155_ (_05695_, _04373_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _57156_ (_05696_, _05695_, _04368_);
  nand _57157_ (_05697_, _05696_, _05694_);
  nand _57158_ (_05698_, _05697_, _05693_);
  nand _57159_ (_05699_, _05698_, _03994_);
  nand _57160_ (_05700_, _04373_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _57161_ (_05701_, _04217_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _57162_ (_05702_, _05701_, _04375_);
  nand _57163_ (_05703_, _05702_, _05700_);
  nand _57164_ (_05704_, _04217_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand _57165_ (_05705_, _04373_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _57166_ (_05706_, _05705_, _04368_);
  nand _57167_ (_05707_, _05706_, _05704_);
  nand _57168_ (_05708_, _05707_, _05703_);
  nand _57169_ (_05709_, _05708_, _04382_);
  nand _57170_ (_05710_, _05709_, _05699_);
  nand _57171_ (_05711_, _05710_, _04396_);
  nand _57172_ (_05712_, _05711_, _05689_);
  or _57173_ (_05713_, _05712_, _03401_);
  and _57174_ (_05714_, _05224_, \oc8051_golden_model_1.IP [4]);
  not _57175_ (_05715_, _05714_);
  and _57176_ (_05716_, _05218_, \oc8051_golden_model_1.PSW [4]);
  not _57177_ (_05717_, _05716_);
  and _57178_ (_05718_, _05221_, \oc8051_golden_model_1.B [4]);
  and _57179_ (_05719_, _05227_, \oc8051_golden_model_1.ACC [4]);
  nor _57180_ (_05720_, _05719_, _05718_);
  and _57181_ (_05721_, _05720_, _05717_);
  and _57182_ (_05722_, _05721_, _05715_);
  and _57183_ (_05723_, _05236_, \oc8051_golden_model_1.TCON [4]);
  and _57184_ (_05724_, _05234_, \oc8051_golden_model_1.TH0 [4]);
  nor _57185_ (_05725_, _05724_, _05723_);
  and _57186_ (_05726_, _05244_, \oc8051_golden_model_1.P1 [4]);
  and _57187_ (_05727_, _05242_, \oc8051_golden_model_1.TL1 [4]);
  nor _57188_ (_05728_, _05727_, _05726_);
  and _57189_ (_05729_, _05728_, _05725_);
  and _57190_ (_05730_, _05248_, \oc8051_golden_model_1.SCON [4]);
  and _57191_ (_05731_, _05251_, \oc8051_golden_model_1.TH1 [4]);
  nor _57192_ (_05732_, _05731_, _05730_);
  and _57193_ (_05733_, _05258_, \oc8051_golden_model_1.TL0 [4]);
  and _57194_ (_05734_, _05254_, \oc8051_golden_model_1.TMOD [4]);
  nor _57195_ (_05735_, _05734_, _05733_);
  and _57196_ (_05736_, _05735_, _05732_);
  and _57197_ (_05737_, _05736_, _05729_);
  and _57198_ (_05738_, _05208_, \oc8051_golden_model_1.PCON [4]);
  not _57199_ (_05739_, _05738_);
  and _57200_ (_05740_, _05185_, \oc8051_golden_model_1.SBUF [4]);
  and _57201_ (_05741_, _05193_, \oc8051_golden_model_1.IE [4]);
  nor _57202_ (_05742_, _05741_, _05740_);
  and _57203_ (_05743_, _05742_, _05739_);
  and _57204_ (_05744_, _05210_, \oc8051_golden_model_1.P2 [4]);
  and _57205_ (_05745_, _05200_, \oc8051_golden_model_1.P3 [4]);
  nor _57206_ (_05746_, _05745_, _05744_);
  and _57207_ (_05747_, _05746_, _05743_);
  and _57208_ (_05748_, _05276_, \oc8051_golden_model_1.P0 [4]);
  not _57209_ (_05749_, _05748_);
  and _57210_ (_05750_, _05266_, \oc8051_golden_model_1.DPH [4]);
  not _57211_ (_05751_, _05750_);
  and _57212_ (_05752_, _05269_, \oc8051_golden_model_1.SP [4]);
  and _57213_ (_05753_, _05272_, \oc8051_golden_model_1.DPL [4]);
  nor _57214_ (_05754_, _05753_, _05752_);
  and _57215_ (_05755_, _05754_, _05751_);
  and _57216_ (_05756_, _05755_, _05749_);
  and _57217_ (_05757_, _05756_, _05747_);
  and _57218_ (_05758_, _05757_, _05737_);
  and _57219_ (_05759_, _05758_, _05722_);
  and _57220_ (_05760_, _05759_, _05713_);
  not _57221_ (_05761_, _05760_);
  and _57222_ (_05762_, _05761_, _05667_);
  and _57223_ (_05763_, _05762_, _05472_);
  and _57224_ (_05764_, _05763_, _05377_);
  nor _57225_ (_05765_, _05764_, _05282_);
  and _57226_ (_05766_, _05764_, _05282_);
  nor _57227_ (_05767_, _05766_, _05765_);
  and _57228_ (_05768_, _05767_, _04544_);
  not _57229_ (_05769_, _03754_);
  nor _57230_ (_05770_, _05769_, _03401_);
  not _57231_ (_05771_, _05770_);
  not _57232_ (_05772_, _04502_);
  nor _57233_ (_05773_, _04739_, _04726_);
  nor _57234_ (_05774_, _05065_, _04489_);
  and _57235_ (_05775_, _05774_, _05773_);
  and _57236_ (_05776_, _05775_, _03438_);
  or _57237_ (_05777_, _05776_, _03401_);
  not _57238_ (_05778_, _04462_);
  not _57239_ (_05779_, _03433_);
  nor _57240_ (_05780_, _04250_, _05779_);
  and _57241_ (_05781_, _03838_, _03565_);
  and _57242_ (_05782_, _05781_, _05780_);
  and _57243_ (_05783_, _05217_, _05782_);
  and _57244_ (_05784_, _05783_, \oc8051_golden_model_1.PSW [7]);
  and _57245_ (_05785_, _05220_, _05782_);
  and _57246_ (_05786_, _05785_, \oc8051_golden_model_1.B [7]);
  nor _57247_ (_05787_, _05786_, _05784_);
  nor _57248_ (_05788_, _03835_, _03565_);
  and _57249_ (_05789_, _05788_, _05780_);
  and _57250_ (_05790_, _05789_, _05199_);
  and _57251_ (_05791_, _05790_, \oc8051_golden_model_1.IP [7]);
  and _57252_ (_05792_, _05226_, _05782_);
  and _57253_ (_05793_, _05792_, \oc8051_golden_model_1.ACC [7]);
  nor _57254_ (_05794_, _05793_, _05791_);
  and _57255_ (_05795_, _05794_, _05787_);
  and _57256_ (_05796_, _05199_, _05782_);
  and _57257_ (_05797_, _05796_, \oc8051_golden_model_1.P3 [7]);
  not _57258_ (_05798_, _05797_);
  and _57259_ (_05799_, _05789_, _05204_);
  and _57260_ (_05800_, _05799_, \oc8051_golden_model_1.TCON [7]);
  and _57261_ (_05801_, _05192_, _05782_);
  and _57262_ (_05802_, _05801_, \oc8051_golden_model_1.P2 [7]);
  nor _57263_ (_05803_, _05802_, _05800_);
  and _57264_ (_05804_, _05803_, _05798_);
  and _57265_ (_05805_, _05789_, _05184_);
  and _57266_ (_05806_, _05805_, \oc8051_golden_model_1.SCON [7]);
  and _57267_ (_05807_, _05789_, _05192_);
  and _57268_ (_05808_, _05807_, \oc8051_golden_model_1.IE [7]);
  nor _57269_ (_05809_, _05808_, _05806_);
  and _57270_ (_05810_, _05205_, \oc8051_golden_model_1.P0 [7]);
  and _57271_ (_05811_, _05184_, _05782_);
  and _57272_ (_05812_, _05811_, \oc8051_golden_model_1.P1 [7]);
  nor _57273_ (_05813_, _05812_, _05810_);
  and _57274_ (_05814_, _05813_, _05809_);
  and _57275_ (_05815_, _05814_, _05804_);
  and _57276_ (_05816_, _05815_, _05795_);
  and _57277_ (_05817_, _05816_, _05177_);
  nor _57278_ (_05818_, _05817_, _05207_);
  or _57279_ (_05819_, _05818_, _05778_);
  not _57280_ (_05820_, _04443_);
  not _57281_ (_05821_, _05176_);
  and _57282_ (_05822_, _05712_, _05422_);
  and _57283_ (_05823_, _04603_, _04439_);
  and _57284_ (_05824_, _05026_, _04843_);
  and _57285_ (_05825_, _05824_, _05823_);
  and _57286_ (_05826_, _05825_, _05822_);
  and _57287_ (_05827_, _05826_, _05327_);
  or _57288_ (_05828_, _05827_, _05821_);
  nand _57289_ (_05829_, _05827_, _05821_);
  and _57290_ (_05830_, _05829_, _05828_);
  or _57291_ (_05831_, _03202_, _03218_);
  or _57292_ (_05832_, _05831_, _05830_);
  not _57293_ (_05833_, _05831_);
  not _57294_ (_05834_, \oc8051_golden_model_1.ACC [7]);
  nor _57295_ (_05835_, _03923_, _05834_);
  and _57296_ (_05836_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and _57297_ (_05837_, _05836_, \oc8051_golden_model_1.PC [6]);
  and _57298_ (_05838_, _05837_, _03278_);
  and _57299_ (_05839_, _05838_, \oc8051_golden_model_1.PC [7]);
  nor _57300_ (_05840_, _05838_, \oc8051_golden_model_1.PC [7]);
  nor _57301_ (_05841_, _05840_, _05839_);
  and _57302_ (_05842_, _05841_, _03923_);
  or _57303_ (_05843_, _05842_, _05835_);
  or _57304_ (_05844_, _05843_, _05833_);
  and _57305_ (_05845_, _05844_, _05832_);
  or _57306_ (_05846_, _05845_, _04438_);
  not _57307_ (_05847_, _04438_);
  nor _57308_ (_05848_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _57309_ (_05849_, _05848_, _03982_);
  nor _57310_ (_05850_, _05849_, _03567_);
  nor _57311_ (_05851_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _57312_ (_05852_, _05851_, _03567_);
  and _57313_ (_05853_, _05852_, _03502_);
  nor _57314_ (_05854_, _05853_, _05850_);
  nor _57315_ (_05855_, _05854_, _03984_);
  not _57316_ (_05856_, _05855_);
  not _57317_ (_05857_, _04478_);
  nand _57318_ (_05858_, _04843_, _05857_);
  not _57319_ (_05859_, _03984_);
  and _57320_ (_05860_, _04478_, _03432_);
  nor _57321_ (_05861_, _05860_, _05859_);
  nand _57322_ (_05862_, _05861_, _05858_);
  and _57323_ (_05863_, _05862_, _05856_);
  not _57324_ (_05864_, _05863_);
  nor _57325_ (_05865_, _05848_, _03982_);
  nor _57326_ (_05866_, _05865_, _05849_);
  nor _57327_ (_05867_, _05866_, _03984_);
  not _57328_ (_05868_, _05867_);
  nand _57329_ (_05869_, _05026_, _05857_);
  and _57330_ (_05870_, _04478_, _03877_);
  nor _57331_ (_05871_, _05870_, _05859_);
  nand _57332_ (_05872_, _05871_, _05869_);
  and _57333_ (_05873_, _05872_, _05868_);
  or _57334_ (_05874_, _04419_, _04478_);
  and _57335_ (_05875_, _04478_, _03471_);
  nor _57336_ (_05876_, _05875_, _05859_);
  nand _57337_ (_05877_, _05876_, _05874_);
  nor _57338_ (_05878_, _03984_, \oc8051_golden_model_1.SP [0]);
  not _57339_ (_05879_, _05878_);
  and _57340_ (_05880_, _05879_, _05877_);
  or _57341_ (_05881_, _05880_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor _57342_ (_05882_, _04603_, _04478_);
  nor _57343_ (_05883_, _04284_, _05857_);
  or _57344_ (_05884_, _05883_, _05882_);
  nand _57345_ (_05885_, _05884_, _03984_);
  nor _57346_ (_05886_, _04553_, _03984_);
  not _57347_ (_05887_, _05886_);
  and _57348_ (_05888_, _05887_, _05885_);
  nand _57349_ (_05889_, _05879_, _05877_);
  or _57350_ (_05890_, _05889_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _57351_ (_05891_, _05890_, _05888_);
  and _57352_ (_05892_, _05891_, _05881_);
  or _57353_ (_05893_, _05889_, \oc8051_golden_model_1.IRAM[10] [7]);
  nand _57354_ (_05894_, _05887_, _05885_);
  or _57355_ (_05895_, _05880_, \oc8051_golden_model_1.IRAM[11] [7]);
  and _57356_ (_05896_, _05895_, _05894_);
  and _57357_ (_05897_, _05896_, _05893_);
  nor _57358_ (_05898_, _05897_, _05892_);
  nand _57359_ (_05899_, _05898_, _05873_);
  not _57360_ (_05900_, _05873_);
  or _57361_ (_05901_, _05880_, \oc8051_golden_model_1.IRAM[13] [7]);
  or _57362_ (_05902_, _05889_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _57363_ (_05903_, _05902_, _05888_);
  and _57364_ (_05904_, _05903_, _05901_);
  or _57365_ (_05905_, _05889_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _57366_ (_05906_, _05880_, \oc8051_golden_model_1.IRAM[15] [7]);
  and _57367_ (_05907_, _05906_, _05894_);
  and _57368_ (_05908_, _05907_, _05905_);
  nor _57369_ (_05909_, _05908_, _05904_);
  nand _57370_ (_05910_, _05909_, _05900_);
  nand _57371_ (_05911_, _05910_, _05899_);
  nand _57372_ (_05912_, _05911_, _05864_);
  or _57373_ (_05913_, _05889_, _05132_);
  or _57374_ (_05914_, _05880_, _05130_);
  and _57375_ (_05915_, _05914_, _05894_);
  nand _57376_ (_05916_, _05915_, _05913_);
  or _57377_ (_05917_, _05889_, _05124_);
  or _57378_ (_05918_, _05880_, _05126_);
  and _57379_ (_05919_, _05918_, _05888_);
  nand _57380_ (_05920_, _05919_, _05917_);
  nand _57381_ (_05921_, _05920_, _05916_);
  nand _57382_ (_05922_, _05921_, _05873_);
  or _57383_ (_05923_, _05889_, _05140_);
  or _57384_ (_05924_, _05880_, _05138_);
  and _57385_ (_05925_, _05924_, _05894_);
  nand _57386_ (_05926_, _05925_, _05923_);
  or _57387_ (_05927_, _05889_, _05144_);
  or _57388_ (_05928_, _05880_, _05146_);
  and _57389_ (_05929_, _05928_, _05888_);
  nand _57390_ (_05930_, _05929_, _05927_);
  nand _57391_ (_05931_, _05930_, _05926_);
  nand _57392_ (_05932_, _05931_, _05900_);
  nand _57393_ (_05933_, _05932_, _05922_);
  nand _57394_ (_05934_, _05933_, _05863_);
  and _57395_ (_05935_, _05934_, _05912_);
  or _57396_ (_05936_, _05935_, _05847_);
  and _57397_ (_05937_, _05936_, _05846_);
  and _57398_ (_05938_, _05937_, _04866_);
  and _57399_ (_05939_, _05760_, _05471_);
  and _57400_ (_05940_, _05568_, _05522_);
  and _57401_ (_05941_, _05616_, _05570_);
  and _57402_ (_05942_, _05941_, _05940_);
  and _57403_ (_05943_, _05664_, _05520_);
  and _57404_ (_05944_, _05943_, _05942_);
  and _57405_ (_05945_, _05944_, _05939_);
  and _57406_ (_05946_, _05945_, _05376_);
  nor _57407_ (_05947_, _05946_, _05282_);
  and _57408_ (_05948_, _05946_, _05282_);
  nor _57409_ (_05949_, _05948_, _05947_);
  and _57410_ (_05950_, _05949_, _04445_);
  or _57411_ (_05951_, _05950_, _05938_);
  and _57412_ (_05952_, _05951_, _05820_);
  not _57413_ (_05953_, _05207_);
  nand _57414_ (_05954_, _05817_, _05953_);
  and _57415_ (_05955_, _05954_, _04443_);
  or _57416_ (_05956_, _05955_, _04746_);
  or _57417_ (_05957_, _05956_, _05952_);
  nor _57418_ (_05958_, _05841_, _03203_);
  nor _57419_ (_05959_, _05958_, _04454_);
  and _57420_ (_05960_, _05959_, _05957_);
  and _57421_ (_05961_, _05821_, _04454_);
  or _57422_ (_05962_, _05961_, _04462_);
  or _57423_ (_05963_, _05962_, _05960_);
  and _57424_ (_05964_, _05963_, _05819_);
  or _57425_ (_05965_, _05964_, _03511_);
  not _57426_ (_05966_, _05237_);
  nor _57427_ (_05967_, _05243_, _05235_);
  and _57428_ (_05968_, _05260_, _05967_);
  and _57429_ (_05969_, _05968_, _05966_);
  and _57430_ (_05970_, _05969_, _05275_);
  not _57431_ (_05971_, _05209_);
  and _57432_ (_05972_, _05253_, _05971_);
  and _57433_ (_05973_, _05972_, _05195_);
  and _57434_ (_05974_, _05210_, \oc8051_golden_model_1.P2INREG [7]);
  and _57435_ (_05975_, _05200_, \oc8051_golden_model_1.P3INREG [7]);
  nor _57436_ (_05976_, _05975_, _05974_);
  and _57437_ (_05977_, _05276_, \oc8051_golden_model_1.P0INREG [7]);
  and _57438_ (_05978_, _05244_, \oc8051_golden_model_1.P1INREG [7]);
  nor _57439_ (_05979_, _05978_, _05977_);
  and _57440_ (_05980_, _05979_, _05976_);
  and _57441_ (_05981_, _05980_, _05230_);
  and _57442_ (_05982_, _05981_, _05973_);
  and _57443_ (_05983_, _05982_, _05970_);
  and _57444_ (_05984_, _05983_, _05177_);
  nand _57445_ (_05985_, _05984_, _03511_);
  and _57446_ (_05986_, _05985_, _03509_);
  and _57447_ (_05987_, _05986_, _05965_);
  nor _57448_ (_05988_, _05817_, _05953_);
  not _57449_ (_05989_, _05988_);
  and _57450_ (_05990_, _05989_, _05954_);
  and _57451_ (_05991_, _05990_, _03508_);
  or _57452_ (_05992_, _05991_, _05987_);
  and _57453_ (_05993_, _05992_, _03200_);
  not _57454_ (_05994_, _05841_);
  or _57455_ (_05995_, _05994_, _03200_);
  nand _57456_ (_05996_, _05995_, _03602_);
  or _57457_ (_05998_, _05996_, _05993_);
  nand _57458_ (_05999_, _05984_, _04053_);
  and _57459_ (_06001_, _05999_, _05998_);
  or _57460_ (_06002_, _06001_, _04478_);
  nand _57461_ (_06004_, _05934_, _05912_);
  or _57462_ (_06005_, _06004_, _03401_);
  and _57463_ (_06007_, _05983_, _04478_);
  nand _57464_ (_06008_, _06007_, _06005_);
  and _57465_ (_06010_, _06008_, _04901_);
  and _57466_ (_06011_, _06010_, _06002_);
  and _57467_ (_06013_, _05205_, \oc8051_golden_model_1.P0INREG [7]);
  not _57468_ (_06014_, _06013_);
  and _57469_ (_06016_, _05811_, \oc8051_golden_model_1.P1INREG [7]);
  and _57470_ (_06017_, _05801_, \oc8051_golden_model_1.P2INREG [7]);
  nor _57471_ (_06019_, _06017_, _06016_);
  and _57472_ (_06020_, _06019_, _06014_);
  and _57473_ (_06022_, _05796_, \oc8051_golden_model_1.P3INREG [7]);
  nor _57474_ (_06023_, _06022_, _05800_);
  and _57475_ (_06025_, _06023_, _05809_);
  and _57476_ (_06026_, _06025_, _06020_);
  and _57477_ (_06028_, _06026_, _05795_);
  and _57478_ (_06029_, _06028_, _05177_);
  nor _57479_ (_06031_, _06029_, _05207_);
  and _57480_ (_06032_, _05207_, \oc8051_golden_model_1.PSW [7]);
  nor _57481_ (_06034_, _06032_, _06031_);
  nor _57482_ (_06035_, _06034_, _04901_);
  or _57483_ (_06036_, _06035_, _03223_);
  or _57484_ (_06037_, _06036_, _06011_);
  not _57485_ (_06038_, _03477_);
  and _57486_ (_06039_, _03492_, _06038_);
  nor _57487_ (_06040_, _06039_, _03401_);
  and _57488_ (_06041_, _05994_, _03223_);
  nor _57489_ (_06042_, _06041_, _06040_);
  and _57490_ (_06043_, _06042_, _06037_);
  not _57491_ (_06044_, _03479_);
  nor _57492_ (_06045_, _06044_, _03401_);
  not _57493_ (_06046_, _06040_);
  nor _57494_ (_06047_, _05176_, _06046_);
  or _57495_ (_06048_, _06047_, _06045_);
  or _57496_ (_06049_, _06048_, _06043_);
  not _57497_ (_06050_, _04784_);
  not _57498_ (_06051_, _06045_);
  or _57499_ (_06052_, _05935_, _06051_);
  and _57500_ (_06053_, _06052_, _06050_);
  and _57501_ (_06054_, _06053_, _06049_);
  not _57502_ (_06055_, _05775_);
  and _57503_ (_06056_, _03704_, _01644_);
  and _57504_ (_06057_, _03713_, _01658_);
  nor _57505_ (_06058_, _06057_, _06056_);
  and _57506_ (_06059_, _03689_, _01662_);
  and _57507_ (_06060_, _03711_, _01670_);
  nor _57508_ (_06061_, _06060_, _06059_);
  and _57509_ (_06062_, _06061_, _06058_);
  and _57510_ (_06063_, _03732_, _01609_);
  and _57511_ (_06064_, _03719_, _01686_);
  nor _57512_ (_06065_, _06064_, _06063_);
  and _57513_ (_06066_, _03721_, _01711_);
  and _57514_ (_06067_, _03693_, _01714_);
  nor _57515_ (_06068_, _06067_, _06066_);
  and _57516_ (_06069_, _06068_, _06065_);
  and _57517_ (_06070_, _06069_, _06062_);
  and _57518_ (_06071_, _03730_, _01701_);
  and _57519_ (_06072_, _03726_, _01693_);
  nor _57520_ (_06073_, _06072_, _06071_);
  and _57521_ (_06074_, _03737_, _01682_);
  and _57522_ (_06075_, _03707_, _01649_);
  nor _57523_ (_06076_, _06075_, _06074_);
  and _57524_ (_06077_, _06076_, _06073_);
  and _57525_ (_06078_, _03698_, _01666_);
  and _57526_ (_06079_, _03735_, _01705_);
  nor _57527_ (_06080_, _06079_, _06078_);
  and _57528_ (_06081_, _03724_, _01697_);
  and _57529_ (_06082_, _03700_, _01674_);
  nor _57530_ (_06083_, _06082_, _06081_);
  and _57531_ (_06084_, _06083_, _06080_);
  and _57532_ (_06085_, _06084_, _06077_);
  and _57533_ (_06086_, _06085_, _06070_);
  not _57534_ (_06087_, _06086_);
  nor _57535_ (_06088_, _06087_, _05176_);
  and _57536_ (_06089_, _03920_, _03742_);
  and _57537_ (_06090_, _03732_, _02207_);
  and _57538_ (_06091_, _03713_, _02181_);
  nor _57539_ (_06093_, _06091_, _06090_);
  and _57540_ (_06095_, _03689_, _02177_);
  and _57541_ (_06096_, _03711_, _02175_);
  nor _57542_ (_06098_, _06096_, _06095_);
  and _57543_ (_06099_, _06098_, _06093_);
  and _57544_ (_06101_, _03704_, _02210_);
  and _57545_ (_06102_, _03719_, _02185_);
  nor _57546_ (_06104_, _06102_, _06101_);
  and _57547_ (_06105_, _03721_, _02201_);
  and _57548_ (_06107_, _03693_, _02189_);
  nor _57549_ (_06108_, _06107_, _06105_);
  and _57550_ (_06110_, _06108_, _06104_);
  and _57551_ (_06111_, _06110_, _06099_);
  and _57552_ (_06113_, _03735_, _02168_);
  and _57553_ (_06114_, _03698_, _02165_);
  nor _57554_ (_06116_, _06114_, _06113_);
  and _57555_ (_06117_, _03737_, _02191_);
  and _57556_ (_06119_, _03707_, _02203_);
  nor _57557_ (_06120_, _06119_, _06117_);
  and _57558_ (_06122_, _06120_, _06116_);
  and _57559_ (_06123_, _03730_, _02198_);
  and _57560_ (_06125_, _03726_, _02213_);
  nor _57561_ (_06126_, _06125_, _06123_);
  and _57562_ (_06127_, _03724_, _02172_);
  and _57563_ (_06128_, _03700_, _02183_);
  nor _57564_ (_06129_, _06128_, _06127_);
  and _57565_ (_06130_, _06129_, _06126_);
  and _57566_ (_06131_, _06130_, _06122_);
  and _57567_ (_06132_, _06131_, _06111_);
  and _57568_ (_06133_, _06132_, _06087_);
  and _57569_ (_06134_, _03689_, _02120_);
  and _57570_ (_06135_, _03721_, _02147_);
  nor _57571_ (_06136_, _06135_, _06134_);
  and _57572_ (_06137_, _03698_, _02114_);
  and _57573_ (_06138_, _03693_, _02134_);
  nor _57574_ (_06139_, _06138_, _06137_);
  and _57575_ (_06140_, _06139_, _06136_);
  and _57576_ (_06141_, _03704_, _02154_);
  and _57577_ (_06142_, _03707_, _02145_);
  nor _57578_ (_06143_, _06142_, _06141_);
  and _57579_ (_06144_, _03711_, _02151_);
  and _57580_ (_06145_, _03713_, _02131_);
  nor _57581_ (_06146_, _06145_, _06144_);
  and _57582_ (_06147_, _06146_, _06143_);
  and _57583_ (_06148_, _06147_, _06140_);
  and _57584_ (_06149_, _03700_, _02128_);
  and _57585_ (_06150_, _03719_, _02126_);
  nor _57586_ (_06151_, _06150_, _06149_);
  and _57587_ (_06152_, _03724_, _02109_);
  and _57588_ (_06153_, _03726_, _02157_);
  nor _57589_ (_06154_, _06153_, _06152_);
  and _57590_ (_06155_, _06154_, _06151_);
  and _57591_ (_06156_, _03730_, _02142_);
  and _57592_ (_06157_, _03732_, _02122_);
  nor _57593_ (_06158_, _06157_, _06156_);
  and _57594_ (_06159_, _03735_, _02112_);
  and _57595_ (_06160_, _03737_, _02136_);
  nor _57596_ (_06161_, _06160_, _06159_);
  and _57597_ (_06162_, _06161_, _06158_);
  and _57598_ (_06163_, _06162_, _06155_);
  and _57599_ (_06164_, _06163_, _06148_);
  and _57600_ (_06165_, _03721_, _02088_);
  and _57601_ (_06166_, _03707_, _02091_);
  nor _57602_ (_06167_, _06166_, _06165_);
  and _57603_ (_06168_, _03730_, _02086_);
  and _57604_ (_06169_, _03737_, _02081_);
  nor _57605_ (_06170_, _06169_, _06168_);
  and _57606_ (_06171_, _06170_, _06167_);
  and _57607_ (_06172_, _03698_, _02053_);
  and _57608_ (_06173_, _03704_, _02098_);
  nor _57609_ (_06174_, _06173_, _06172_);
  and _57610_ (_06175_, _03719_, _02075_);
  and _57611_ (_06176_, _03693_, _02079_);
  nor _57612_ (_06177_, _06176_, _06175_);
  and _57613_ (_06178_, _06177_, _06174_);
  and _57614_ (_06179_, _06178_, _06171_);
  and _57615_ (_06180_, _03689_, _02066_);
  and _57616_ (_06181_, _03724_, _02060_);
  nor _57617_ (_06182_, _06181_, _06180_);
  and _57618_ (_06183_, _03735_, _02056_);
  and _57619_ (_06184_, _03732_, _02064_);
  nor _57620_ (_06185_, _06184_, _06183_);
  and _57621_ (_06186_, _06185_, _06182_);
  and _57622_ (_06187_, _03726_, _02101_);
  and _57623_ (_06188_, _03700_, _02073_);
  nor _57624_ (_06189_, _06188_, _06187_);
  and _57625_ (_06190_, _03711_, _02095_);
  and _57626_ (_06191_, _03713_, _02071_);
  nor _57627_ (_06192_, _06191_, _06190_);
  and _57628_ (_06193_, _06192_, _06189_);
  and _57629_ (_06194_, _06193_, _06186_);
  and _57630_ (_06195_, _06194_, _06179_);
  and _57631_ (_06196_, _06195_, _06164_);
  and _57632_ (_06197_, _06196_, _06133_);
  nor _57633_ (_06198_, _04317_, _04109_);
  and _57634_ (_06199_, _06198_, _06197_);
  and _57635_ (_06200_, _06199_, _06089_);
  and _57636_ (_06201_, _06200_, \oc8051_golden_model_1.DPH [7]);
  not _57637_ (_06202_, _04109_);
  and _57638_ (_06203_, _04317_, _06202_);
  nor _57639_ (_06204_, _03920_, _03742_);
  and _57640_ (_06205_, _06204_, _06197_);
  and _57641_ (_06206_, _06205_, _06203_);
  and _57642_ (_06207_, _06206_, \oc8051_golden_model_1.TH1 [7]);
  nor _57643_ (_06208_, _06207_, _06201_);
  and _57644_ (_06209_, _04317_, _04109_);
  and _57645_ (_06210_, _06209_, _06089_);
  not _57646_ (_06211_, _06164_);
  and _57647_ (_06212_, _06195_, _06211_);
  and _57648_ (_06213_, _06212_, _06133_);
  and _57649_ (_06214_, _06213_, _06210_);
  and _57650_ (_06215_, _06214_, \oc8051_golden_model_1.P2INREG [7]);
  not _57651_ (_06216_, _06215_);
  not _57652_ (_06217_, _03742_);
  and _57653_ (_06218_, _03920_, _06217_);
  and _57654_ (_06219_, _06218_, _06203_);
  and _57655_ (_06220_, _06219_, _06197_);
  and _57656_ (_06221_, _06220_, \oc8051_golden_model_1.TMOD [7]);
  not _57657_ (_06222_, _04317_);
  and _57658_ (_06223_, _06222_, _04109_);
  and _57659_ (_06224_, _06218_, _06197_);
  and _57660_ (_06225_, _06224_, _06223_);
  and _57661_ (_06226_, _06225_, \oc8051_golden_model_1.TL0 [7]);
  nor _57662_ (_06227_, _06226_, _06221_);
  and _57663_ (_06228_, _06227_, _06216_);
  and _57664_ (_06229_, _06218_, _06209_);
  and _57665_ (_06230_, _06229_, _06213_);
  and _57666_ (_06231_, _06230_, \oc8051_golden_model_1.IE [7]);
  not _57667_ (_06232_, _06231_);
  not _57668_ (_06233_, _06195_);
  and _57669_ (_06234_, _06233_, _06164_);
  and _57670_ (_06235_, _06234_, _06133_);
  and _57671_ (_06236_, _06235_, _06229_);
  and _57672_ (_06237_, _06236_, \oc8051_golden_model_1.SCON [7]);
  and _57673_ (_06238_, _06235_, _06219_);
  and _57674_ (_06239_, _06238_, \oc8051_golden_model_1.SBUF [7]);
  nor _57675_ (_06240_, _06239_, _06237_);
  and _57676_ (_06241_, _06240_, _06232_);
  and _57677_ (_06242_, _06210_, _06197_);
  and _57678_ (_06243_, _06242_, \oc8051_golden_model_1.P0INREG [7]);
  not _57679_ (_06244_, _06243_);
  and _57680_ (_06245_, _06235_, _06210_);
  and _57681_ (_06246_, _06245_, \oc8051_golden_model_1.P1INREG [7]);
  nor _57682_ (_06247_, _06195_, _06164_);
  and _57683_ (_06248_, _06247_, _06133_);
  and _57684_ (_06249_, _06248_, _06210_);
  and _57685_ (_06250_, _06249_, \oc8051_golden_model_1.P3INREG [7]);
  nor _57686_ (_06251_, _06250_, _06246_);
  and _57687_ (_06252_, _06251_, _06244_);
  and _57688_ (_06253_, _06252_, _06241_);
  and _57689_ (_06254_, _06253_, _06228_);
  and _57690_ (_06255_, _06254_, _06208_);
  and _57691_ (_06256_, _06209_, _06205_);
  and _57692_ (_06257_, _06256_, \oc8051_golden_model_1.TH0 [7]);
  and _57693_ (_06258_, _06218_, _06199_);
  and _57694_ (_06259_, _06258_, \oc8051_golden_model_1.TL1 [7]);
  nor _57695_ (_06260_, _06259_, _06257_);
  not _57696_ (_06261_, _03920_);
  and _57697_ (_06262_, _06261_, _03742_);
  and _57698_ (_06263_, _06262_, _06199_);
  and _57699_ (_06264_, _06263_, \oc8051_golden_model_1.PCON [7]);
  and _57700_ (_06265_, _06224_, _06209_);
  and _57701_ (_06266_, _06265_, \oc8051_golden_model_1.TCON [7]);
  nor _57702_ (_06267_, _06266_, _06264_);
  and _57703_ (_06268_, _06267_, _06260_);
  and _57704_ (_06269_, _06248_, _06229_);
  and _57705_ (_06270_, _06269_, \oc8051_golden_model_1.IP [7]);
  nor _57706_ (_06271_, _06132_, _06086_);
  and _57707_ (_06272_, _06271_, _06210_);
  and _57708_ (_06273_, _06272_, _06247_);
  and _57709_ (_06274_, _06273_, \oc8051_golden_model_1.B [7]);
  nor _57710_ (_06275_, _06274_, _06270_);
  and _57711_ (_06276_, _06272_, _06234_);
  and _57712_ (_06277_, _06276_, \oc8051_golden_model_1.PSW [7]);
  and _57713_ (_06278_, _06272_, _06212_);
  and _57714_ (_06279_, _06278_, \oc8051_golden_model_1.ACC [7]);
  nor _57715_ (_06280_, _06279_, _06277_);
  and _57716_ (_06281_, _06280_, _06275_);
  and _57717_ (_06282_, _06197_, _06089_);
  and _57718_ (_06283_, _06282_, _06203_);
  and _57719_ (_06284_, _06283_, \oc8051_golden_model_1.SP [7]);
  and _57720_ (_06285_, _06282_, _06223_);
  and _57721_ (_06286_, _06285_, \oc8051_golden_model_1.DPL [7]);
  nor _57722_ (_06287_, _06286_, _06284_);
  and _57723_ (_06288_, _06287_, _06281_);
  and _57724_ (_06289_, _06288_, _06268_);
  and _57725_ (_06290_, _06289_, _06255_);
  not _57726_ (_06291_, _06290_);
  nor _57727_ (_06292_, _06291_, _06088_);
  nor _57728_ (_06293_, _06292_, _06050_);
  or _57729_ (_06294_, _06293_, _06055_);
  or _57730_ (_06295_, _06294_, _06054_);
  and _57731_ (_06296_, _06295_, _05777_);
  and _57732_ (_06297_, _06087_, _03439_);
  or _57733_ (_06298_, _06297_, _03189_);
  or _57734_ (_06299_, _06298_, _06296_);
  and _57735_ (_06300_, _05994_, _03189_);
  nor _57736_ (_06301_, _06300_, _04500_);
  and _57737_ (_06302_, _06301_, _06299_);
  nor _57738_ (_06303_, _06086_, _05281_);
  and _57739_ (_06304_, _06086_, _05281_);
  nor _57740_ (_06305_, _06304_, _06303_);
  and _57741_ (_06306_, _06305_, _04500_);
  or _57742_ (_06307_, _06306_, _06302_);
  and _57743_ (_06308_, _06307_, _05772_);
  nor _57744_ (_06309_, _05281_, _05834_);
  and _57745_ (_06310_, _05281_, _05834_);
  nor _57746_ (_06311_, _06310_, _06309_);
  and _57747_ (_06312_, _06311_, _04502_);
  or _57748_ (_06313_, _06312_, _06308_);
  and _57749_ (_06314_, _06313_, _05771_);
  and _57750_ (_06315_, _06303_, _04506_);
  or _57751_ (_06316_, _06315_, _04497_);
  or _57752_ (_06317_, _06316_, _06314_);
  or _57753_ (_06318_, _06309_, _04498_);
  and _57754_ (_06319_, _06318_, _06317_);
  or _57755_ (_06320_, _06319_, _03192_);
  and _57756_ (_06321_, _05994_, _03192_);
  nor _57757_ (_06322_, _06321_, _04516_);
  and _57758_ (_06323_, _06322_, _06320_);
  not _57759_ (_06324_, _04518_);
  and _57760_ (_06325_, _06304_, _06324_);
  nor _57761_ (_06326_, _06325_, _04519_);
  or _57762_ (_06327_, _06326_, _06323_);
  not _57763_ (_06328_, _03179_);
  nand _57764_ (_06329_, _06310_, _04518_);
  and _57765_ (_06330_, _06329_, _06328_);
  and _57766_ (_06331_, _06330_, _06327_);
  nand _57767_ (_06332_, _05841_, _03179_);
  nand _57768_ (_06333_, _06332_, _04709_);
  or _57769_ (_06334_, _06333_, _06331_);
  not _57770_ (_06335_, _04681_);
  or _57771_ (_06336_, _05830_, _04709_);
  and _57772_ (_06337_, _06336_, _06335_);
  and _57773_ (_06338_, _06337_, _06334_);
  and _57774_ (_06339_, _05830_, _04681_);
  or _57775_ (_06340_, _06339_, _04527_);
  or _57776_ (_06341_, _06340_, _06338_);
  not _57777_ (_06342_, _04526_);
  not _57778_ (_06343_, _04527_);
  or _57779_ (_06344_, _05880_, \oc8051_golden_model_1.IRAM[1] [6]);
  or _57780_ (_06345_, _05889_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _57781_ (_06346_, _06345_, _05888_);
  and _57782_ (_06347_, _06346_, _06344_);
  or _57783_ (_06348_, _05889_, \oc8051_golden_model_1.IRAM[2] [6]);
  or _57784_ (_06349_, _05880_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _57785_ (_06350_, _06349_, _05894_);
  and _57786_ (_06351_, _06350_, _06348_);
  nor _57787_ (_06352_, _06351_, _06347_);
  nand _57788_ (_06353_, _06352_, _05873_);
  or _57789_ (_06354_, _05880_, \oc8051_golden_model_1.IRAM[5] [6]);
  or _57790_ (_06355_, _05889_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _57791_ (_06356_, _06355_, _05888_);
  and _57792_ (_06357_, _06356_, _06354_);
  or _57793_ (_06358_, _05889_, \oc8051_golden_model_1.IRAM[6] [6]);
  or _57794_ (_06359_, _05880_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _57795_ (_06360_, _06359_, _05894_);
  and _57796_ (_06361_, _06360_, _06358_);
  nor _57797_ (_06362_, _06361_, _06357_);
  nand _57798_ (_06363_, _06362_, _05900_);
  nand _57799_ (_06364_, _06363_, _06353_);
  nand _57800_ (_06365_, _06364_, _05863_);
  or _57801_ (_06366_, _05889_, \oc8051_golden_model_1.IRAM[8] [6]);
  or _57802_ (_06367_, _05880_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand _57803_ (_06368_, _06367_, _06366_);
  nand _57804_ (_06369_, _06368_, _05888_);
  or _57805_ (_06370_, _05889_, \oc8051_golden_model_1.IRAM[10] [6]);
  or _57806_ (_06371_, _05880_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _57807_ (_06372_, _06371_, _06370_);
  nand _57808_ (_06373_, _06372_, _05894_);
  nand _57809_ (_06374_, _06373_, _06369_);
  nand _57810_ (_06375_, _06374_, _05873_);
  or _57811_ (_06376_, _05889_, \oc8051_golden_model_1.IRAM[12] [6]);
  or _57812_ (_06377_, _05880_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand _57813_ (_06378_, _06377_, _06376_);
  nand _57814_ (_06379_, _06378_, _05888_);
  or _57815_ (_06380_, _05889_, \oc8051_golden_model_1.IRAM[14] [6]);
  or _57816_ (_06381_, _05880_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _57817_ (_06382_, _06381_, _06380_);
  nand _57818_ (_06383_, _06382_, _05894_);
  nand _57819_ (_06384_, _06383_, _06379_);
  nand _57820_ (_06385_, _06384_, _05900_);
  nand _57821_ (_06386_, _06385_, _06375_);
  nand _57822_ (_06387_, _06386_, _05864_);
  nand _57823_ (_06388_, _06387_, _06365_);
  or _57824_ (_06389_, _05880_, \oc8051_golden_model_1.IRAM[1] [1]);
  or _57825_ (_06390_, _05889_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _57826_ (_06391_, _06390_, _05888_);
  and _57827_ (_06392_, _06391_, _06389_);
  or _57828_ (_06393_, _05889_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _57829_ (_06394_, _05880_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _57830_ (_06395_, _06394_, _05894_);
  and _57831_ (_06396_, _06395_, _06393_);
  nor _57832_ (_06397_, _06396_, _06392_);
  nand _57833_ (_06398_, _06397_, _05873_);
  or _57834_ (_06399_, _05880_, \oc8051_golden_model_1.IRAM[5] [1]);
  or _57835_ (_06400_, _05889_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _57836_ (_06401_, _06400_, _05888_);
  and _57837_ (_06402_, _06401_, _06399_);
  or _57838_ (_06403_, _05889_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _57839_ (_06404_, _05880_, \oc8051_golden_model_1.IRAM[7] [1]);
  and _57840_ (_06405_, _06404_, _05894_);
  and _57841_ (_06406_, _06405_, _06403_);
  nor _57842_ (_06407_, _06406_, _06402_);
  nand _57843_ (_06408_, _06407_, _05900_);
  nand _57844_ (_06409_, _06408_, _06398_);
  nand _57845_ (_06410_, _06409_, _05863_);
  or _57846_ (_06411_, _05889_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _57847_ (_06412_, _05880_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand _57848_ (_06413_, _06412_, _06411_);
  nand _57849_ (_06414_, _06413_, _05888_);
  or _57850_ (_06415_, _05889_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _57851_ (_06416_, _05880_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _57852_ (_06417_, _06416_, _06415_);
  nand _57853_ (_06418_, _06417_, _05894_);
  nand _57854_ (_06419_, _06418_, _06414_);
  nand _57855_ (_06420_, _06419_, _05873_);
  or _57856_ (_06421_, _05889_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _57857_ (_06422_, _05880_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand _57858_ (_06423_, _06422_, _06421_);
  nand _57859_ (_06424_, _06423_, _05888_);
  or _57860_ (_06425_, _05889_, \oc8051_golden_model_1.IRAM[14] [1]);
  or _57861_ (_06426_, _05880_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _57862_ (_06427_, _06426_, _06425_);
  nand _57863_ (_06428_, _06427_, _05894_);
  nand _57864_ (_06429_, _06428_, _06424_);
  nand _57865_ (_06430_, _06429_, _05900_);
  nand _57866_ (_06431_, _06430_, _06420_);
  nand _57867_ (_06432_, _06431_, _05864_);
  nand _57868_ (_06433_, _06432_, _06410_);
  or _57869_ (_06434_, _05880_, \oc8051_golden_model_1.IRAM[1] [0]);
  or _57870_ (_06435_, _05889_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _57871_ (_06436_, _06435_, _05888_);
  and _57872_ (_06437_, _06436_, _06434_);
  or _57873_ (_06438_, _05889_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _57874_ (_06439_, _05880_, \oc8051_golden_model_1.IRAM[3] [0]);
  and _57875_ (_06440_, _06439_, _05894_);
  and _57876_ (_06441_, _06440_, _06438_);
  nor _57877_ (_06442_, _06441_, _06437_);
  nand _57878_ (_06443_, _06442_, _05873_);
  or _57879_ (_06444_, _05880_, \oc8051_golden_model_1.IRAM[5] [0]);
  or _57880_ (_06445_, _05889_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _57881_ (_06446_, _06445_, _05888_);
  and _57882_ (_06447_, _06446_, _06444_);
  or _57883_ (_06448_, _05889_, \oc8051_golden_model_1.IRAM[6] [0]);
  or _57884_ (_06449_, _05880_, \oc8051_golden_model_1.IRAM[7] [0]);
  and _57885_ (_06450_, _06449_, _05894_);
  and _57886_ (_06451_, _06450_, _06448_);
  nor _57887_ (_06452_, _06451_, _06447_);
  nand _57888_ (_06453_, _06452_, _05900_);
  nand _57889_ (_06454_, _06453_, _06443_);
  nand _57890_ (_06455_, _06454_, _05863_);
  or _57891_ (_06456_, _05889_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _57892_ (_06457_, _05880_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _57893_ (_06458_, _06457_, _06456_);
  nand _57894_ (_06459_, _06458_, _05888_);
  or _57895_ (_06460_, _05889_, \oc8051_golden_model_1.IRAM[10] [0]);
  or _57896_ (_06461_, _05880_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _57897_ (_06462_, _06461_, _06460_);
  nand _57898_ (_06463_, _06462_, _05894_);
  nand _57899_ (_06464_, _06463_, _06459_);
  nand _57900_ (_06465_, _06464_, _05873_);
  or _57901_ (_06466_, _05889_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _57902_ (_06467_, _05880_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand _57903_ (_06468_, _06467_, _06466_);
  nand _57904_ (_06469_, _06468_, _05888_);
  or _57905_ (_06470_, _05889_, \oc8051_golden_model_1.IRAM[14] [0]);
  or _57906_ (_06471_, _05880_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _57907_ (_06472_, _06471_, _06470_);
  nand _57908_ (_06473_, _06472_, _05894_);
  nand _57909_ (_06474_, _06473_, _06469_);
  nand _57910_ (_06475_, _06474_, _05900_);
  nand _57911_ (_06476_, _06475_, _06465_);
  nand _57912_ (_06477_, _06476_, _05864_);
  nand _57913_ (_06478_, _06477_, _06455_);
  and _57914_ (_06479_, _06478_, _06433_);
  or _57915_ (_06480_, _05880_, \oc8051_golden_model_1.IRAM[1] [3]);
  or _57916_ (_06481_, _05889_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _57917_ (_06482_, _06481_, _05888_);
  and _57918_ (_06483_, _06482_, _06480_);
  or _57919_ (_06484_, _05889_, \oc8051_golden_model_1.IRAM[2] [3]);
  or _57920_ (_06485_, _05880_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _57921_ (_06486_, _06485_, _05894_);
  and _57922_ (_06487_, _06486_, _06484_);
  nor _57923_ (_06488_, _06487_, _06483_);
  nand _57924_ (_06489_, _06488_, _05873_);
  or _57925_ (_06490_, _05880_, \oc8051_golden_model_1.IRAM[5] [3]);
  or _57926_ (_06491_, _05889_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _57927_ (_06492_, _06491_, _05888_);
  and _57928_ (_06493_, _06492_, _06490_);
  or _57929_ (_06494_, _05889_, \oc8051_golden_model_1.IRAM[6] [3]);
  or _57930_ (_06495_, _05880_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _57931_ (_06496_, _06495_, _05894_);
  and _57932_ (_06497_, _06496_, _06494_);
  nor _57933_ (_06498_, _06497_, _06493_);
  nand _57934_ (_06499_, _06498_, _05900_);
  nand _57935_ (_06500_, _06499_, _06489_);
  nand _57936_ (_06501_, _06500_, _05863_);
  or _57937_ (_06502_, _05889_, \oc8051_golden_model_1.IRAM[8] [3]);
  or _57938_ (_06503_, _05880_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand _57939_ (_06504_, _06503_, _06502_);
  nand _57940_ (_06505_, _06504_, _05888_);
  or _57941_ (_06506_, _05889_, \oc8051_golden_model_1.IRAM[10] [3]);
  or _57942_ (_06507_, _05880_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _57943_ (_06508_, _06507_, _06506_);
  nand _57944_ (_06509_, _06508_, _05894_);
  nand _57945_ (_06510_, _06509_, _06505_);
  nand _57946_ (_06511_, _06510_, _05873_);
  or _57947_ (_06512_, _05889_, \oc8051_golden_model_1.IRAM[12] [3]);
  or _57948_ (_06513_, _05880_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand _57949_ (_06514_, _06513_, _06512_);
  nand _57950_ (_06515_, _06514_, _05888_);
  or _57951_ (_06516_, _05889_, \oc8051_golden_model_1.IRAM[14] [3]);
  or _57952_ (_06517_, _05880_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _57953_ (_06518_, _06517_, _06516_);
  nand _57954_ (_06519_, _06518_, _05894_);
  nand _57955_ (_06520_, _06519_, _06515_);
  nand _57956_ (_06521_, _06520_, _05900_);
  nand _57957_ (_06522_, _06521_, _06511_);
  nand _57958_ (_06523_, _06522_, _05864_);
  nand _57959_ (_06524_, _06523_, _06501_);
  or _57960_ (_06525_, _05880_, \oc8051_golden_model_1.IRAM[1] [2]);
  or _57961_ (_06526_, _05889_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _57962_ (_06527_, _06526_, _05888_);
  and _57963_ (_06528_, _06527_, _06525_);
  or _57964_ (_06529_, _05889_, \oc8051_golden_model_1.IRAM[2] [2]);
  or _57965_ (_06530_, _05880_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _57966_ (_06531_, _06530_, _05894_);
  and _57967_ (_06532_, _06531_, _06529_);
  nor _57968_ (_06533_, _06532_, _06528_);
  nand _57969_ (_06534_, _06533_, _05873_);
  or _57970_ (_06535_, _05880_, \oc8051_golden_model_1.IRAM[5] [2]);
  or _57971_ (_06536_, _05889_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _57972_ (_06537_, _06536_, _05888_);
  and _57973_ (_06538_, _06537_, _06535_);
  or _57974_ (_06539_, _05889_, \oc8051_golden_model_1.IRAM[6] [2]);
  or _57975_ (_06540_, _05880_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _57976_ (_06541_, _06540_, _05894_);
  and _57977_ (_06542_, _06541_, _06539_);
  nor _57978_ (_06543_, _06542_, _06538_);
  nand _57979_ (_06544_, _06543_, _05900_);
  nand _57980_ (_06545_, _06544_, _06534_);
  nand _57981_ (_06546_, _06545_, _05863_);
  or _57982_ (_06547_, _05889_, \oc8051_golden_model_1.IRAM[8] [2]);
  or _57983_ (_06548_, _05880_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand _57984_ (_06549_, _06548_, _06547_);
  nand _57985_ (_06550_, _06549_, _05888_);
  or _57986_ (_06551_, _05889_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _57987_ (_06552_, _05880_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _57988_ (_06553_, _06552_, _06551_);
  nand _57989_ (_06554_, _06553_, _05894_);
  nand _57990_ (_06555_, _06554_, _06550_);
  nand _57991_ (_06556_, _06555_, _05873_);
  or _57992_ (_06557_, _05889_, \oc8051_golden_model_1.IRAM[12] [2]);
  or _57993_ (_06558_, _05880_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand _57994_ (_06559_, _06558_, _06557_);
  nand _57995_ (_06560_, _06559_, _05888_);
  or _57996_ (_06561_, _05889_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _57997_ (_06562_, _05880_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _57998_ (_06563_, _06562_, _06561_);
  nand _57999_ (_06564_, _06563_, _05894_);
  nand _58000_ (_06565_, _06564_, _06560_);
  nand _58001_ (_06566_, _06565_, _05900_);
  nand _58002_ (_06567_, _06566_, _06556_);
  nand _58003_ (_06568_, _06567_, _05864_);
  nand _58004_ (_06569_, _06568_, _06546_);
  and _58005_ (_06570_, _06569_, _06524_);
  and _58006_ (_06571_, _06570_, _06479_);
  or _58007_ (_06572_, _05880_, \oc8051_golden_model_1.IRAM[1] [5]);
  or _58008_ (_06573_, _05889_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _58009_ (_06574_, _06573_, _05888_);
  and _58010_ (_06575_, _06574_, _06572_);
  or _58011_ (_06576_, _05889_, \oc8051_golden_model_1.IRAM[2] [5]);
  or _58012_ (_06577_, _05880_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _58013_ (_06578_, _06577_, _05894_);
  and _58014_ (_06579_, _06578_, _06576_);
  nor _58015_ (_06580_, _06579_, _06575_);
  nand _58016_ (_06581_, _06580_, _05873_);
  or _58017_ (_06582_, _05880_, \oc8051_golden_model_1.IRAM[5] [5]);
  or _58018_ (_06583_, _05889_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _58019_ (_06584_, _06583_, _05888_);
  and _58020_ (_06585_, _06584_, _06582_);
  or _58021_ (_06586_, _05889_, \oc8051_golden_model_1.IRAM[6] [5]);
  or _58022_ (_06587_, _05880_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _58023_ (_06588_, _06587_, _05894_);
  and _58024_ (_06589_, _06588_, _06586_);
  nor _58025_ (_06590_, _06589_, _06585_);
  nand _58026_ (_06591_, _06590_, _05900_);
  nand _58027_ (_06592_, _06591_, _06581_);
  nand _58028_ (_06593_, _06592_, _05863_);
  or _58029_ (_06594_, _05889_, \oc8051_golden_model_1.IRAM[8] [5]);
  or _58030_ (_06595_, _05880_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand _58031_ (_06596_, _06595_, _06594_);
  nand _58032_ (_06597_, _06596_, _05888_);
  or _58033_ (_06598_, _05889_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _58034_ (_06599_, _05880_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _58035_ (_06600_, _06599_, _06598_);
  nand _58036_ (_06601_, _06600_, _05894_);
  nand _58037_ (_06602_, _06601_, _06597_);
  nand _58038_ (_06603_, _06602_, _05873_);
  or _58039_ (_06604_, _05889_, \oc8051_golden_model_1.IRAM[12] [5]);
  or _58040_ (_06605_, _05880_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand _58041_ (_06606_, _06605_, _06604_);
  nand _58042_ (_06607_, _06606_, _05888_);
  or _58043_ (_06608_, _05889_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _58044_ (_06609_, _05880_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _58045_ (_06610_, _06609_, _06608_);
  nand _58046_ (_06611_, _06610_, _05894_);
  nand _58047_ (_06612_, _06611_, _06607_);
  nand _58048_ (_06613_, _06612_, _05900_);
  nand _58049_ (_06614_, _06613_, _06603_);
  nand _58050_ (_06615_, _06614_, _05864_);
  nand _58051_ (_06616_, _06615_, _06593_);
  or _58052_ (_06617_, _05880_, \oc8051_golden_model_1.IRAM[1] [4]);
  or _58053_ (_06618_, _05889_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _58054_ (_06619_, _06618_, _05888_);
  and _58055_ (_06620_, _06619_, _06617_);
  or _58056_ (_06621_, _05889_, \oc8051_golden_model_1.IRAM[2] [4]);
  or _58057_ (_06622_, _05880_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _58058_ (_06623_, _06622_, _05894_);
  and _58059_ (_06624_, _06623_, _06621_);
  nor _58060_ (_06625_, _06624_, _06620_);
  nand _58061_ (_06626_, _06625_, _05873_);
  or _58062_ (_06627_, _05880_, \oc8051_golden_model_1.IRAM[5] [4]);
  or _58063_ (_06628_, _05889_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _58064_ (_06629_, _06628_, _05888_);
  and _58065_ (_06630_, _06629_, _06627_);
  or _58066_ (_06631_, _05889_, \oc8051_golden_model_1.IRAM[6] [4]);
  or _58067_ (_06632_, _05880_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _58068_ (_06633_, _06632_, _05894_);
  and _58069_ (_06634_, _06633_, _06631_);
  nor _58070_ (_06635_, _06634_, _06630_);
  nand _58071_ (_06636_, _06635_, _05900_);
  nand _58072_ (_06637_, _06636_, _06626_);
  nand _58073_ (_06638_, _06637_, _05863_);
  or _58074_ (_06639_, _05889_, \oc8051_golden_model_1.IRAM[8] [4]);
  or _58075_ (_06640_, _05880_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand _58076_ (_06641_, _06640_, _06639_);
  nand _58077_ (_06642_, _06641_, _05888_);
  or _58078_ (_06643_, _05889_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _58079_ (_06644_, _05880_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _58080_ (_06645_, _06644_, _06643_);
  nand _58081_ (_06646_, _06645_, _05894_);
  nand _58082_ (_06647_, _06646_, _06642_);
  nand _58083_ (_06648_, _06647_, _05873_);
  or _58084_ (_06649_, _05889_, \oc8051_golden_model_1.IRAM[12] [4]);
  or _58085_ (_06650_, _05880_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand _58086_ (_06651_, _06650_, _06649_);
  nand _58087_ (_06652_, _06651_, _05888_);
  or _58088_ (_06653_, _05889_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _58089_ (_06654_, _05880_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _58090_ (_06655_, _06654_, _06653_);
  nand _58091_ (_06656_, _06655_, _05894_);
  nand _58092_ (_06657_, _06656_, _06652_);
  nand _58093_ (_06658_, _06657_, _05900_);
  nand _58094_ (_06659_, _06658_, _06648_);
  nand _58095_ (_06660_, _06659_, _05864_);
  nand _58096_ (_06661_, _06660_, _06638_);
  and _58097_ (_06662_, _06661_, _06616_);
  and _58098_ (_06663_, _06662_, _06571_);
  and _58099_ (_06664_, _06663_, _06388_);
  nor _58100_ (_06665_, _06664_, _06004_);
  and _58101_ (_06666_, _06664_, _06004_);
  or _58102_ (_06667_, _06666_, _06665_);
  or _58103_ (_06668_, _06667_, _06343_);
  and _58104_ (_06669_, _06668_, _06342_);
  and _58105_ (_06670_, _06669_, _06341_);
  and _58106_ (_06671_, _05949_, _04526_);
  or _58107_ (_06672_, _06671_, _03641_);
  or _58108_ (_06673_, _06672_, _06670_);
  and _58109_ (_06674_, _02891_, \oc8051_golden_model_1.PC [2]);
  and _58110_ (_06675_, _06674_, \oc8051_golden_model_1.PC [3]);
  and _58111_ (_06676_, _06675_, _05837_);
  and _58112_ (_06677_, _06676_, \oc8051_golden_model_1.PC [7]);
  nor _58113_ (_06678_, _06676_, \oc8051_golden_model_1.PC [7]);
  nor _58114_ (_06679_, _06678_, _06677_);
  not _58115_ (_06680_, _06679_);
  nand _58116_ (_06681_, _06680_, _03641_);
  and _58117_ (_06682_, _06681_, _06673_);
  or _58118_ (_06683_, _06682_, _03160_);
  and _58119_ (_06684_, _05994_, _03160_);
  nor _58120_ (_06685_, _06684_, _03435_);
  and _58121_ (_06686_, _06685_, _06683_);
  nand _58122_ (_06687_, _06031_, _03435_);
  nor _58123_ (_06688_, _04205_, _04766_);
  nand _58124_ (_06689_, _06688_, _06687_);
  or _58125_ (_06690_, _06689_, _06686_);
  not _58126_ (_06691_, _04693_);
  nor _58127_ (_06692_, _04603_, _04439_);
  nor _58128_ (_06693_, _05026_, _04843_);
  and _58129_ (_06694_, _06693_, _06692_);
  nor _58130_ (_06695_, _05712_, _05422_);
  and _58131_ (_06697_, _06695_, _06694_);
  or _58132_ (_06698_, _06697_, _05821_);
  and _58133_ (_06699_, _05327_, _05176_);
  nor _58134_ (_06700_, _05327_, _05176_);
  nor _58135_ (_06701_, _06700_, _06699_);
  not _58136_ (_06702_, _06701_);
  nand _58137_ (_06703_, _06702_, _06697_);
  and _58138_ (_06704_, _06703_, _06698_);
  or _58139_ (_06705_, _06704_, _06688_);
  and _58140_ (_06706_, _06705_, _06691_);
  and _58141_ (_06707_, _06706_, _06690_);
  and _58142_ (_06708_, _06704_, _04693_);
  or _58143_ (_06709_, _06708_, _04540_);
  or _58144_ (_06710_, _06709_, _06707_);
  not _58145_ (_06711_, _04544_);
  not _58146_ (_06712_, _04540_);
  and _58147_ (_06713_, _06387_, _06365_);
  and _58148_ (_06714_, _06432_, _06410_);
  and _58149_ (_06715_, _06477_, _06455_);
  and _58150_ (_06716_, _06715_, _06714_);
  and _58151_ (_06717_, _06523_, _06501_);
  and _58152_ (_06718_, _06568_, _06546_);
  and _58153_ (_06719_, _06718_, _06717_);
  and _58154_ (_06720_, _06719_, _06716_);
  and _58155_ (_06721_, _06615_, _06593_);
  and _58156_ (_06722_, _06660_, _06638_);
  and _58157_ (_06723_, _06722_, _06721_);
  and _58158_ (_06724_, _06723_, _06720_);
  and _58159_ (_06725_, _06724_, _06713_);
  nor _58160_ (_06726_, _06725_, _06004_);
  and _58161_ (_06727_, _06725_, _06004_);
  or _58162_ (_06728_, _06727_, _06726_);
  or _58163_ (_06729_, _06728_, _06712_);
  and _58164_ (_06730_, _06729_, _06711_);
  and _58165_ (_06731_, _06730_, _06710_);
  or _58166_ (_06732_, _06731_, _05768_);
  and _58167_ (_06733_, _06732_, _04794_);
  or _58168_ (_06734_, _06733_, _05123_);
  and _58169_ (_06735_, _06734_, _05122_);
  not _58170_ (_06736_, \oc8051_golden_model_1.PC [15]);
  and _58171_ (_06737_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and _58172_ (_06738_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and _58173_ (_06739_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and _58174_ (_06740_, _06739_, _06738_);
  and _58175_ (_06741_, _06740_, _05839_);
  and _58176_ (_06742_, _06741_, _06737_);
  and _58177_ (_06743_, _06742_, \oc8051_golden_model_1.PC [14]);
  and _58178_ (_06744_, _06743_, _06736_);
  nor _58179_ (_06745_, _06743_, _06736_);
  or _58180_ (_06746_, _06745_, _06744_);
  not _58181_ (_06747_, _06746_);
  nor _58182_ (_06748_, _06747_, _03641_);
  and _58183_ (_06749_, _06740_, _06677_);
  and _58184_ (_06750_, _06749_, _06737_);
  and _58185_ (_06751_, _06750_, \oc8051_golden_model_1.PC [14]);
  and _58186_ (_06752_, _06751_, _06736_);
  nor _58187_ (_06753_, _06751_, _06736_);
  or _58188_ (_06754_, _06753_, _06752_);
  and _58189_ (_06755_, _06754_, _03641_);
  or _58190_ (_06756_, _06755_, _06748_);
  and _58191_ (_06757_, _06756_, _05117_);
  and _58192_ (_06758_, _06757_, _05120_);
  or _58193_ (_40514_, _06758_, _06735_);
  not _58194_ (_06759_, \oc8051_golden_model_1.B [7]);
  nor _58195_ (_06760_, _42963_, _06759_);
  nor _58196_ (_06761_, _05221_, _06759_);
  not _58197_ (_06762_, _05221_);
  nor _58198_ (_06763_, _06762_, _05176_);
  or _58199_ (_06764_, _06763_, _06761_);
  or _58200_ (_06765_, _06764_, _06039_);
  nor _58201_ (_06766_, _05785_, _06759_);
  and _58202_ (_06767_, _05818_, _05785_);
  or _58203_ (_06768_, _06767_, _06766_);
  and _58204_ (_06769_, _06768_, _03512_);
  and _58205_ (_06770_, _05949_, _05221_);
  or _58206_ (_06771_, _06770_, _06761_);
  or _58207_ (_06772_, _06771_, _04444_);
  and _58208_ (_06773_, _05221_, \oc8051_golden_model_1.ACC [7]);
  or _58209_ (_06774_, _06773_, _06761_);
  and _58210_ (_06775_, _06774_, _04426_);
  nor _58211_ (_06776_, _04426_, _06759_);
  or _58212_ (_06777_, _06776_, _03570_);
  or _58213_ (_06778_, _06777_, _06775_);
  and _58214_ (_06779_, _06778_, _03517_);
  and _58215_ (_06780_, _06779_, _06772_);
  and _58216_ (_06781_, _05954_, _05785_);
  or _58217_ (_06782_, _06781_, _06766_);
  and _58218_ (_06783_, _06782_, _03516_);
  or _58219_ (_06784_, _06783_, _03568_);
  or _58220_ (_06785_, _06784_, _06780_);
  or _58221_ (_06786_, _06764_, _03983_);
  and _58222_ (_06787_, _06786_, _06785_);
  or _58223_ (_06788_, _06787_, _03575_);
  or _58224_ (_06789_, _06774_, _03583_);
  and _58225_ (_06790_, _06789_, _03513_);
  and _58226_ (_06791_, _06790_, _06788_);
  or _58227_ (_06792_, _06791_, _06769_);
  and _58228_ (_06793_, _06792_, _03506_);
  and _58229_ (_06794_, _03637_, _03596_);
  or _58230_ (_06795_, _06766_, _05989_);
  and _58231_ (_06796_, _06795_, _03505_);
  and _58232_ (_06797_, _06796_, _06782_);
  or _58233_ (_06798_, _06797_, _06794_);
  or _58234_ (_06799_, _06798_, _06793_);
  not _58235_ (_06800_, _06794_);
  and _58236_ (_06801_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and _58237_ (_06802_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and _58238_ (_06803_, _06802_, _06801_);
  and _58239_ (_06804_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and _58240_ (_06805_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor _58241_ (_06806_, _06805_, _06804_);
  nor _58242_ (_06807_, _06806_, _06803_);
  and _58243_ (_06808_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and _58244_ (_06809_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and _58245_ (_06810_, _06809_, _06808_);
  and _58246_ (_06811_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and _58247_ (_06812_, _06811_, _06802_);
  and _58248_ (_06813_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  nor _58249_ (_06814_, _06811_, _06802_);
  nor _58250_ (_06815_, _06814_, _06812_);
  and _58251_ (_06816_, _06815_, _06813_);
  nor _58252_ (_06817_, _06816_, _06812_);
  and _58253_ (_06818_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and _58254_ (_06819_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and _58255_ (_06820_, _06819_, _06818_);
  nor _58256_ (_06821_, _06819_, _06818_);
  nor _58257_ (_06822_, _06821_, _06820_);
  not _58258_ (_06823_, _06822_);
  nor _58259_ (_06824_, _06823_, _06817_);
  and _58260_ (_06825_, _06823_, _06817_);
  nor _58261_ (_06826_, _06825_, _06824_);
  and _58262_ (_06827_, _06826_, _06810_);
  nor _58263_ (_06828_, _06826_, _06810_);
  nor _58264_ (_06829_, _06828_, _06827_);
  and _58265_ (_06830_, _06829_, _06807_);
  and _58266_ (_06831_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and _58267_ (_06832_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and _58268_ (_06833_, _06832_, _06831_);
  nor _58269_ (_06834_, _06832_, _06831_);
  nor _58270_ (_06835_, _06834_, _06833_);
  and _58271_ (_06836_, _06835_, _06803_);
  nor _58272_ (_06837_, _06835_, _06803_);
  nor _58273_ (_06838_, _06837_, _06836_);
  and _58274_ (_06839_, _06838_, _06820_);
  nor _58275_ (_06840_, _06838_, _06820_);
  nor _58276_ (_06841_, _06840_, _06839_);
  and _58277_ (_06842_, _06841_, _06801_);
  nor _58278_ (_06843_, _06841_, _06801_);
  nor _58279_ (_06844_, _06843_, _06842_);
  and _58280_ (_06845_, _06844_, _06830_);
  nor _58281_ (_06846_, _06827_, _06824_);
  not _58282_ (_06847_, _06846_);
  nor _58283_ (_06848_, _06844_, _06830_);
  nor _58284_ (_06849_, _06848_, _06845_);
  and _58285_ (_06850_, _06849_, _06847_);
  nor _58286_ (_06851_, _06850_, _06845_);
  nor _58287_ (_06852_, _06839_, _06836_);
  not _58288_ (_06853_, _06852_);
  and _58289_ (_06854_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and _58290_ (_06855_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and _58291_ (_06856_, _06855_, _06854_);
  nor _58292_ (_06857_, _06855_, _06854_);
  nor _58293_ (_06858_, _06857_, _06856_);
  and _58294_ (_06859_, _06858_, _06833_);
  nor _58295_ (_06860_, _06858_, _06833_);
  nor _58296_ (_06861_, _06860_, _06859_);
  and _58297_ (_06862_, _06861_, _06842_);
  nor _58298_ (_06863_, _06861_, _06842_);
  nor _58299_ (_06864_, _06863_, _06862_);
  and _58300_ (_06865_, _06864_, _06853_);
  nor _58301_ (_06866_, _06864_, _06853_);
  nor _58302_ (_06867_, _06866_, _06865_);
  not _58303_ (_06868_, _06867_);
  nor _58304_ (_06869_, _06868_, _06851_);
  and _58305_ (_06870_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not _58306_ (_06871_, _06870_);
  nor _58307_ (_06872_, _06871_, _06832_);
  nor _58308_ (_06873_, _06872_, _06859_);
  nor _58309_ (_06874_, _06865_, _06862_);
  nor _58310_ (_06875_, _06874_, _06873_);
  and _58311_ (_06876_, _06874_, _06873_);
  nor _58312_ (_06877_, _06876_, _06875_);
  and _58313_ (_06878_, _06877_, _06869_);
  or _58314_ (_06879_, _06875_, _06856_);
  or _58315_ (_06880_, _06879_, _06878_);
  and _58316_ (_06881_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  and _58317_ (_06882_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and _58318_ (_06883_, _06882_, _06881_);
  not _58319_ (_06884_, _06881_);
  and _58320_ (_06885_, _06882_, _06884_);
  and _58321_ (_06886_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and _58322_ (_06887_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and _58323_ (_06888_, _06887_, _06802_);
  and _58324_ (_06889_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  and _58325_ (_06890_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  nor _58326_ (_06891_, _06890_, _06889_);
  nor _58327_ (_06892_, _06891_, _06888_);
  and _58328_ (_06893_, _06892_, _06886_);
  nor _58329_ (_06894_, _06892_, _06886_);
  nor _58330_ (_06895_, _06894_, _06893_);
  and _58331_ (_06896_, _06895_, _06885_);
  nor _58332_ (_06897_, _06896_, _06883_);
  nor _58333_ (_06898_, _06815_, _06813_);
  nor _58334_ (_06899_, _06898_, _06816_);
  not _58335_ (_06900_, _06899_);
  nor _58336_ (_06901_, _06900_, _06897_);
  and _58337_ (_06902_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and _58338_ (_06903_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and _58339_ (_06904_, _06903_, _06902_);
  nor _58340_ (_06905_, _06893_, _06888_);
  nor _58341_ (_06906_, _06809_, _06808_);
  nor _58342_ (_06907_, _06906_, _06810_);
  not _58343_ (_06908_, _06907_);
  nor _58344_ (_06909_, _06908_, _06905_);
  and _58345_ (_06910_, _06908_, _06905_);
  nor _58346_ (_06911_, _06910_, _06909_);
  and _58347_ (_06912_, _06911_, _06904_);
  nor _58348_ (_06913_, _06911_, _06904_);
  nor _58349_ (_06914_, _06913_, _06912_);
  and _58350_ (_06915_, _06900_, _06897_);
  nor _58351_ (_06916_, _06915_, _06901_);
  and _58352_ (_06917_, _06916_, _06914_);
  nor _58353_ (_06918_, _06917_, _06901_);
  not _58354_ (_06919_, _06918_);
  nor _58355_ (_06920_, _06829_, _06807_);
  nor _58356_ (_06921_, _06920_, _06830_);
  and _58357_ (_06922_, _06921_, _06919_);
  nor _58358_ (_06923_, _06912_, _06909_);
  not _58359_ (_06924_, _06923_);
  nor _58360_ (_06925_, _06921_, _06919_);
  nor _58361_ (_06926_, _06925_, _06922_);
  and _58362_ (_06927_, _06926_, _06924_);
  nor _58363_ (_06928_, _06927_, _06922_);
  nor _58364_ (_06929_, _06849_, _06847_);
  nor _58365_ (_06930_, _06929_, _06850_);
  not _58366_ (_06931_, _06930_);
  nor _58367_ (_06932_, _06931_, _06928_);
  and _58368_ (_06933_, _06868_, _06851_);
  nor _58369_ (_06934_, _06933_, _06869_);
  and _58370_ (_06935_, _06934_, _06932_);
  and _58371_ (_06936_, _06935_, _06877_);
  and _58372_ (_06937_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and _58373_ (_06938_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and _58374_ (_06939_, _06938_, _06937_);
  and _58375_ (_06940_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and _58376_ (_06941_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor _58377_ (_06942_, _06941_, _06881_);
  nor _58378_ (_06943_, _06942_, _06939_);
  and _58379_ (_06944_, _06943_, _06940_);
  nor _58380_ (_06945_, _06944_, _06939_);
  and _58381_ (_06946_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor _58382_ (_06947_, _06946_, _06937_);
  nor _58383_ (_06948_, _06947_, _06883_);
  not _58384_ (_06949_, _06948_);
  nor _58385_ (_06950_, _06949_, _06945_);
  and _58386_ (_06951_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and _58387_ (_06952_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and _58388_ (_06953_, _06952_, _06887_);
  nor _58389_ (_06954_, _06952_, _06887_);
  nor _58390_ (_06955_, _06954_, _06953_);
  and _58391_ (_06956_, _06955_, _06951_);
  nor _58392_ (_06957_, _06955_, _06951_);
  nor _58393_ (_06958_, _06957_, _06956_);
  and _58394_ (_06959_, _06949_, _06945_);
  nor _58395_ (_06960_, _06959_, _06950_);
  and _58396_ (_06961_, _06960_, _06958_);
  nor _58397_ (_06962_, _06961_, _06950_);
  nor _58398_ (_06963_, _06895_, _06885_);
  nor _58399_ (_06964_, _06963_, _06896_);
  not _58400_ (_06965_, _06964_);
  nor _58401_ (_06966_, _06965_, _06962_);
  and _58402_ (_06967_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and _58403_ (_06968_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and _58404_ (_06969_, _06968_, _06967_);
  nor _58405_ (_06970_, _06956_, _06953_);
  nor _58406_ (_06971_, _06903_, _06902_);
  nor _58407_ (_06972_, _06971_, _06904_);
  not _58408_ (_06973_, _06972_);
  nor _58409_ (_06974_, _06973_, _06970_);
  and _58410_ (_06975_, _06973_, _06970_);
  nor _58411_ (_06976_, _06975_, _06974_);
  and _58412_ (_06977_, _06976_, _06969_);
  nor _58413_ (_06978_, _06976_, _06969_);
  nor _58414_ (_06979_, _06978_, _06977_);
  and _58415_ (_06980_, _06965_, _06962_);
  nor _58416_ (_06981_, _06980_, _06966_);
  and _58417_ (_06982_, _06981_, _06979_);
  nor _58418_ (_06983_, _06982_, _06966_);
  nor _58419_ (_06984_, _06916_, _06914_);
  nor _58420_ (_06985_, _06984_, _06917_);
  not _58421_ (_06986_, _06985_);
  nor _58422_ (_06987_, _06986_, _06983_);
  nor _58423_ (_06988_, _06977_, _06974_);
  not _58424_ (_06989_, _06988_);
  and _58425_ (_06990_, _06986_, _06983_);
  nor _58426_ (_06991_, _06990_, _06987_);
  and _58427_ (_06992_, _06991_, _06989_);
  nor _58428_ (_06993_, _06992_, _06987_);
  nor _58429_ (_06994_, _06926_, _06924_);
  nor _58430_ (_06995_, _06994_, _06927_);
  not _58431_ (_06996_, _06995_);
  nor _58432_ (_06997_, _06996_, _06993_);
  and _58433_ (_06998_, _06931_, _06928_);
  nor _58434_ (_06999_, _06998_, _06932_);
  and _58435_ (_07000_, _06999_, _06997_);
  nor _58436_ (_07001_, _06934_, _06932_);
  nor _58437_ (_07002_, _07001_, _06935_);
  and _58438_ (_07003_, _07002_, _07000_);
  nor _58439_ (_07004_, _07002_, _07000_);
  and _58440_ (_07005_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and _58441_ (_07006_, _07005_, _06881_);
  and _58442_ (_07007_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and _58443_ (_07008_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor _58444_ (_07009_, _07008_, _06938_);
  nor _58445_ (_07010_, _07009_, _07006_);
  and _58446_ (_07011_, _07010_, _07007_);
  nor _58447_ (_07012_, _07011_, _07006_);
  not _58448_ (_07013_, _07012_);
  nor _58449_ (_07014_, _06943_, _06940_);
  nor _58450_ (_07015_, _07014_, _06944_);
  and _58451_ (_07016_, _07015_, _07013_);
  and _58452_ (_07017_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and _58453_ (_07018_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and _58454_ (_07019_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and _58455_ (_07020_, _07019_, _07018_);
  nor _58456_ (_07021_, _07019_, _07018_);
  nor _58457_ (_07022_, _07021_, _07020_);
  and _58458_ (_07023_, _07022_, _07017_);
  nor _58459_ (_07024_, _07022_, _07017_);
  nor _58460_ (_07025_, _07024_, _07023_);
  nor _58461_ (_07026_, _07015_, _07013_);
  nor _58462_ (_07027_, _07026_, _07016_);
  and _58463_ (_07028_, _07027_, _07025_);
  nor _58464_ (_07029_, _07028_, _07016_);
  nor _58465_ (_07030_, _06960_, _06958_);
  nor _58466_ (_07031_, _07030_, _06961_);
  not _58467_ (_07032_, _07031_);
  nor _58468_ (_07033_, _07032_, _07029_);
  and _58469_ (_07034_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and _58470_ (_07035_, _07034_, _06968_);
  nor _58471_ (_07036_, _07023_, _07020_);
  nor _58472_ (_07037_, _06968_, _06967_);
  nor _58473_ (_07038_, _07037_, _06969_);
  not _58474_ (_07039_, _07038_);
  nor _58475_ (_07040_, _07039_, _07036_);
  and _58476_ (_07041_, _07039_, _07036_);
  nor _58477_ (_07042_, _07041_, _07040_);
  and _58478_ (_07043_, _07042_, _07035_);
  nor _58479_ (_07044_, _07042_, _07035_);
  nor _58480_ (_07045_, _07044_, _07043_);
  and _58481_ (_07046_, _07032_, _07029_);
  nor _58482_ (_07047_, _07046_, _07033_);
  and _58483_ (_07048_, _07047_, _07045_);
  nor _58484_ (_07049_, _07048_, _07033_);
  nor _58485_ (_07050_, _06981_, _06979_);
  nor _58486_ (_07051_, _07050_, _06982_);
  not _58487_ (_07052_, _07051_);
  nor _58488_ (_07053_, _07052_, _07049_);
  nor _58489_ (_07054_, _07043_, _07040_);
  not _58490_ (_07055_, _07054_);
  and _58491_ (_07056_, _07052_, _07049_);
  nor _58492_ (_07057_, _07056_, _07053_);
  and _58493_ (_07058_, _07057_, _07055_);
  nor _58494_ (_07059_, _07058_, _07053_);
  nor _58495_ (_07060_, _06991_, _06989_);
  nor _58496_ (_07061_, _07060_, _06992_);
  not _58497_ (_07062_, _07061_);
  nor _58498_ (_07063_, _07062_, _07059_);
  and _58499_ (_07064_, _06996_, _06993_);
  nor _58500_ (_07065_, _07064_, _06997_);
  and _58501_ (_07066_, _07065_, _07063_);
  nor _58502_ (_07067_, _06999_, _06997_);
  nor _58503_ (_07068_, _07067_, _07000_);
  nand _58504_ (_07069_, _07068_, _07066_);
  and _58505_ (_07070_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and _58506_ (_07071_, _07070_, _07005_);
  and _58507_ (_07072_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor _58508_ (_07073_, _07070_, _07005_);
  nor _58509_ (_07074_, _07073_, _07071_);
  and _58510_ (_07075_, _07074_, _07072_);
  nor _58511_ (_07076_, _07075_, _07071_);
  not _58512_ (_07077_, _07076_);
  nor _58513_ (_07078_, _07010_, _07007_);
  nor _58514_ (_07079_, _07078_, _07011_);
  and _58515_ (_07080_, _07079_, _07077_);
  and _58516_ (_07081_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and _58517_ (_07082_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and _58518_ (_07083_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and _58519_ (_07084_, _07083_, _07082_);
  nor _58520_ (_07085_, _07083_, _07082_);
  nor _58521_ (_07086_, _07085_, _07084_);
  and _58522_ (_07087_, _07086_, _07081_);
  nor _58523_ (_07088_, _07086_, _07081_);
  nor _58524_ (_07089_, _07088_, _07087_);
  nor _58525_ (_07090_, _07079_, _07077_);
  nor _58526_ (_07091_, _07090_, _07080_);
  and _58527_ (_07092_, _07091_, _07089_);
  nor _58528_ (_07093_, _07092_, _07080_);
  not _58529_ (_07094_, _07093_);
  nor _58530_ (_07095_, _07027_, _07025_);
  nor _58531_ (_07096_, _07095_, _07028_);
  and _58532_ (_07097_, _07096_, _07094_);
  nor _58533_ (_07098_, _07087_, _07084_);
  and _58534_ (_07099_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and _58535_ (_07100_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor _58536_ (_07101_, _07100_, _07099_);
  nor _58537_ (_07102_, _07101_, _07035_);
  not _58538_ (_07103_, _07102_);
  nor _58539_ (_07104_, _07103_, _07098_);
  and _58540_ (_07105_, _07103_, _07098_);
  nor _58541_ (_07106_, _07105_, _07104_);
  nor _58542_ (_07107_, _07096_, _07094_);
  nor _58543_ (_07108_, _07107_, _07097_);
  and _58544_ (_07109_, _07108_, _07106_);
  nor _58545_ (_07110_, _07109_, _07097_);
  nor _58546_ (_07111_, _07047_, _07045_);
  nor _58547_ (_07112_, _07111_, _07048_);
  not _58548_ (_07113_, _07112_);
  nor _58549_ (_07114_, _07113_, _07110_);
  and _58550_ (_07115_, _07113_, _07110_);
  nor _58551_ (_07116_, _07115_, _07114_);
  and _58552_ (_07117_, _07116_, _07104_);
  nor _58553_ (_07118_, _07117_, _07114_);
  nor _58554_ (_07119_, _07057_, _07055_);
  nor _58555_ (_07120_, _07119_, _07058_);
  not _58556_ (_07121_, _07120_);
  nor _58557_ (_07122_, _07121_, _07118_);
  and _58558_ (_07123_, _07062_, _07059_);
  nor _58559_ (_07124_, _07123_, _07063_);
  and _58560_ (_07125_, _07124_, _07122_);
  nor _58561_ (_07126_, _07065_, _07063_);
  nor _58562_ (_07127_, _07126_, _07066_);
  and _58563_ (_07128_, _07127_, _07125_);
  nor _58564_ (_07129_, _07127_, _07125_);
  nor _58565_ (_07130_, _07129_, _07128_);
  and _58566_ (_07131_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and _58567_ (_07132_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and _58568_ (_07133_, _07132_, _07131_);
  and _58569_ (_07134_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor _58570_ (_07135_, _07132_, _07131_);
  nor _58571_ (_07136_, _07135_, _07133_);
  and _58572_ (_07137_, _07136_, _07134_);
  nor _58573_ (_07138_, _07137_, _07133_);
  not _58574_ (_07139_, _07138_);
  nor _58575_ (_07140_, _07074_, _07072_);
  nor _58576_ (_07141_, _07140_, _07075_);
  and _58577_ (_07142_, _07141_, _07139_);
  and _58578_ (_07143_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and _58579_ (_07144_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and _58580_ (_07145_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and _58581_ (_07146_, _07145_, _07144_);
  nor _58582_ (_07147_, _07145_, _07144_);
  nor _58583_ (_07148_, _07147_, _07146_);
  and _58584_ (_07149_, _07148_, _07143_);
  nor _58585_ (_07150_, _07148_, _07143_);
  nor _58586_ (_07151_, _07150_, _07149_);
  nor _58587_ (_07152_, _07141_, _07139_);
  nor _58588_ (_07153_, _07152_, _07142_);
  and _58589_ (_07154_, _07153_, _07151_);
  nor _58590_ (_07155_, _07154_, _07142_);
  not _58591_ (_07156_, _07155_);
  nor _58592_ (_07157_, _07091_, _07089_);
  nor _58593_ (_07158_, _07157_, _07092_);
  and _58594_ (_07159_, _07158_, _07156_);
  not _58595_ (_07160_, _07034_);
  nor _58596_ (_07161_, _07149_, _07146_);
  nor _58597_ (_07162_, _07161_, _07160_);
  and _58598_ (_07163_, _07161_, _07160_);
  nor _58599_ (_07164_, _07163_, _07162_);
  nor _58600_ (_07165_, _07158_, _07156_);
  nor _58601_ (_07166_, _07165_, _07159_);
  and _58602_ (_07167_, _07166_, _07164_);
  nor _58603_ (_07168_, _07167_, _07159_);
  not _58604_ (_07169_, _07168_);
  nor _58605_ (_07170_, _07108_, _07106_);
  nor _58606_ (_07171_, _07170_, _07109_);
  and _58607_ (_07172_, _07171_, _07169_);
  nor _58608_ (_07173_, _07171_, _07169_);
  nor _58609_ (_07174_, _07173_, _07172_);
  and _58610_ (_07175_, _07174_, _07162_);
  nor _58611_ (_07176_, _07175_, _07172_);
  nor _58612_ (_07177_, _07116_, _07104_);
  nor _58613_ (_07178_, _07177_, _07117_);
  not _58614_ (_07179_, _07178_);
  nor _58615_ (_07180_, _07179_, _07176_);
  and _58616_ (_07181_, _07121_, _07118_);
  nor _58617_ (_07182_, _07181_, _07122_);
  and _58618_ (_07183_, _07182_, _07180_);
  nor _58619_ (_07184_, _07124_, _07122_);
  nor _58620_ (_07185_, _07184_, _07125_);
  nand _58621_ (_07186_, _07185_, _07183_);
  or _58622_ (_07187_, _07185_, _07183_);
  and _58623_ (_07188_, _07187_, _07186_);
  and _58624_ (_07189_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and _58625_ (_07190_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and _58626_ (_07191_, _07190_, _07189_);
  and _58627_ (_07192_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor _58628_ (_07193_, _07190_, _07189_);
  nor _58629_ (_07194_, _07193_, _07191_);
  and _58630_ (_07195_, _07194_, _07192_);
  nor _58631_ (_07196_, _07195_, _07191_);
  not _58632_ (_07197_, _07196_);
  nor _58633_ (_07198_, _07136_, _07134_);
  nor _58634_ (_07199_, _07198_, _07137_);
  and _58635_ (_07200_, _07199_, _07197_);
  and _58636_ (_07201_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and _58637_ (_07202_, _07201_, _07145_);
  and _58638_ (_07203_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and _58639_ (_07204_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor _58640_ (_07205_, _07204_, _07203_);
  nor _58641_ (_07206_, _07205_, _07202_);
  nor _58642_ (_07207_, _07199_, _07197_);
  nor _58643_ (_07208_, _07207_, _07200_);
  and _58644_ (_07209_, _07208_, _07206_);
  nor _58645_ (_07210_, _07209_, _07200_);
  not _58646_ (_07211_, _07210_);
  nor _58647_ (_07212_, _07153_, _07151_);
  nor _58648_ (_07213_, _07212_, _07154_);
  and _58649_ (_07214_, _07213_, _07211_);
  nor _58650_ (_07215_, _07213_, _07211_);
  nor _58651_ (_07216_, _07215_, _07214_);
  and _58652_ (_07217_, _07216_, _07202_);
  nor _58653_ (_07218_, _07217_, _07214_);
  not _58654_ (_07219_, _07218_);
  nor _58655_ (_07220_, _07166_, _07164_);
  nor _58656_ (_07221_, _07220_, _07167_);
  and _58657_ (_07222_, _07221_, _07219_);
  nor _58658_ (_07223_, _07174_, _07162_);
  nor _58659_ (_07224_, _07223_, _07175_);
  and _58660_ (_07225_, _07224_, _07222_);
  and _58661_ (_07226_, _07179_, _07176_);
  nor _58662_ (_07227_, _07226_, _07180_);
  and _58663_ (_07228_, _07227_, _07225_);
  nor _58664_ (_07229_, _07182_, _07180_);
  nor _58665_ (_07230_, _07229_, _07183_);
  and _58666_ (_07231_, _07230_, _07228_);
  nor _58667_ (_07232_, _07230_, _07228_);
  nor _58668_ (_07233_, _07232_, _07231_);
  and _58669_ (_07234_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and _58670_ (_07235_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and _58671_ (_07236_, _07235_, _07234_);
  and _58672_ (_07237_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor _58673_ (_07238_, _07235_, _07234_);
  nor _58674_ (_07239_, _07238_, _07236_);
  and _58675_ (_07240_, _07239_, _07237_);
  nor _58676_ (_07241_, _07240_, _07236_);
  not _58677_ (_07242_, _07241_);
  nor _58678_ (_07243_, _07194_, _07192_);
  nor _58679_ (_07244_, _07243_, _07195_);
  and _58680_ (_07245_, _07244_, _07242_);
  nor _58681_ (_07246_, _07244_, _07242_);
  nor _58682_ (_07247_, _07246_, _07245_);
  and _58683_ (_07248_, _07247_, _07201_);
  nor _58684_ (_07249_, _07248_, _07245_);
  not _58685_ (_07250_, _07249_);
  nor _58686_ (_07251_, _07208_, _07206_);
  nor _58687_ (_07252_, _07251_, _07209_);
  and _58688_ (_07253_, _07252_, _07250_);
  nor _58689_ (_07254_, _07216_, _07202_);
  nor _58690_ (_07255_, _07254_, _07217_);
  and _58691_ (_07256_, _07255_, _07253_);
  nor _58692_ (_07257_, _07221_, _07219_);
  nor _58693_ (_07258_, _07257_, _07222_);
  and _58694_ (_07259_, _07258_, _07256_);
  nor _58695_ (_07260_, _07224_, _07222_);
  nor _58696_ (_07261_, _07260_, _07225_);
  and _58697_ (_07262_, _07261_, _07259_);
  nor _58698_ (_07263_, _07227_, _07225_);
  nor _58699_ (_07264_, _07263_, _07228_);
  and _58700_ (_07265_, _07264_, _07262_);
  and _58701_ (_07266_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and _58702_ (_07267_, _07266_, _07235_);
  nor _58703_ (_07268_, _07239_, _07237_);
  nor _58704_ (_07269_, _07268_, _07240_);
  and _58705_ (_07270_, _07269_, _07267_);
  nor _58706_ (_07271_, _07247_, _07201_);
  nor _58707_ (_07272_, _07271_, _07248_);
  and _58708_ (_07273_, _07272_, _07270_);
  nor _58709_ (_07274_, _07252_, _07250_);
  nor _58710_ (_07275_, _07274_, _07253_);
  and _58711_ (_07276_, _07275_, _07273_);
  nor _58712_ (_07277_, _07255_, _07253_);
  nor _58713_ (_07278_, _07277_, _07256_);
  and _58714_ (_07279_, _07278_, _07276_);
  nor _58715_ (_07280_, _07258_, _07256_);
  nor _58716_ (_07281_, _07280_, _07259_);
  and _58717_ (_07282_, _07281_, _07279_);
  nor _58718_ (_07283_, _07261_, _07259_);
  nor _58719_ (_07284_, _07283_, _07262_);
  and _58720_ (_07285_, _07284_, _07282_);
  nor _58721_ (_07286_, _07264_, _07262_);
  nor _58722_ (_07287_, _07286_, _07265_);
  and _58723_ (_07288_, _07287_, _07285_);
  nor _58724_ (_07289_, _07288_, _07265_);
  not _58725_ (_07290_, _07289_);
  and _58726_ (_07291_, _07290_, _07233_);
  or _58727_ (_07292_, _07291_, _07231_);
  nand _58728_ (_07293_, _07292_, _07188_);
  and _58729_ (_07294_, _07293_, _07186_);
  not _58730_ (_07295_, _07294_);
  and _58731_ (_07296_, _07295_, _07130_);
  or _58732_ (_07297_, _07296_, _07128_);
  or _58733_ (_07298_, _07068_, _07066_);
  and _58734_ (_07299_, _07298_, _07069_);
  nand _58735_ (_07300_, _07299_, _07297_);
  and _58736_ (_07301_, _07300_, _07069_);
  nor _58737_ (_07302_, _07301_, _07004_);
  or _58738_ (_07303_, _07302_, _07003_);
  nor _58739_ (_07304_, _06935_, _06869_);
  and _58740_ (_07305_, _07304_, _06877_);
  nor _58741_ (_07306_, _07304_, _06877_);
  or _58742_ (_07307_, _07306_, _07305_);
  and _58743_ (_07308_, _07307_, _07303_);
  or _58744_ (_07309_, _07308_, _06936_);
  or _58745_ (_07310_, _07309_, _06880_);
  or _58746_ (_07311_, _07310_, _06800_);
  and _58747_ (_07312_, _07311_, _03500_);
  and _58748_ (_07313_, _07312_, _06799_);
  not _58749_ (_07314_, _06039_);
  not _58750_ (_07315_, _05785_);
  nor _58751_ (_07316_, _06034_, _07315_);
  or _58752_ (_07317_, _07316_, _06766_);
  and _58753_ (_07318_, _07317_, _03499_);
  or _58754_ (_07319_, _07318_, _07314_);
  or _58755_ (_07320_, _07319_, _07313_);
  and _58756_ (_07321_, _07320_, _06765_);
  or _58757_ (_07322_, _07321_, _03479_);
  and _58758_ (_07323_, _05935_, _05221_);
  or _58759_ (_07324_, _06761_, _06044_);
  or _58760_ (_07325_, _07324_, _07323_);
  and _58761_ (_07326_, _07325_, _03474_);
  and _58762_ (_07327_, _07326_, _07322_);
  and _58763_ (_07328_, _03637_, _03186_);
  nor _58764_ (_07329_, _06292_, _06762_);
  or _58765_ (_07330_, _07329_, _06761_);
  and _58766_ (_07331_, _07330_, _03221_);
  or _58767_ (_07332_, _07331_, _07328_);
  or _58768_ (_07333_, _07332_, _07327_);
  not _58769_ (_07334_, \oc8051_golden_model_1.B [1]);
  nor _58770_ (_07335_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.B [4]);
  nor _58771_ (_07336_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [3]);
  and _58772_ (_07337_, _07336_, _07335_);
  and _58773_ (_07338_, _07337_, _07334_);
  nor _58774_ (_07339_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not _58775_ (_07340_, \oc8051_golden_model_1.B [0]);
  and _58776_ (_07341_, _07340_, \oc8051_golden_model_1.ACC [7]);
  and _58777_ (_07342_, _07341_, _07339_);
  and _58778_ (_07343_, _07342_, _07338_);
  and _58779_ (_07344_, _07339_, _07338_);
  or _58780_ (_07345_, _07344_, _05834_);
  not _58781_ (_07346_, \oc8051_golden_model_1.ACC [6]);
  and _58782_ (_07347_, \oc8051_golden_model_1.B [0], _07346_);
  nor _58783_ (_07348_, _07347_, _05834_);
  nor _58784_ (_07349_, _07348_, _07334_);
  and _58785_ (_07350_, _07339_, _07337_);
  not _58786_ (_07351_, _07350_);
  nor _58787_ (_07352_, _07351_, _07349_);
  nor _58788_ (_07353_, _07352_, _07345_);
  nor _58789_ (_07354_, _07353_, _07343_);
  and _58790_ (_07355_, _07352_, \oc8051_golden_model_1.B [0]);
  nor _58791_ (_07356_, _07355_, _07346_);
  and _58792_ (_07357_, _07356_, _07334_);
  nor _58793_ (_07358_, _07356_, _07334_);
  nor _58794_ (_07359_, _07358_, _07357_);
  nor _58795_ (_07360_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor _58796_ (_07361_, _07360_, _07005_);
  nor _58797_ (_07362_, _07361_, \oc8051_golden_model_1.ACC [4]);
  nor _58798_ (_07363_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and _58799_ (_07364_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor _58800_ (_07365_, _07364_, _07340_);
  nor _58801_ (_07366_, _07365_, _07363_);
  nor _58802_ (_07367_, _07366_, _07362_);
  not _58803_ (_07368_, _07367_);
  and _58804_ (_07369_, _07368_, _07359_);
  nor _58805_ (_07370_, _07354_, \oc8051_golden_model_1.B [2]);
  nor _58806_ (_07371_, _07370_, _07357_);
  not _58807_ (_07372_, _07371_);
  nor _58808_ (_07373_, _07372_, _07369_);
  not _58809_ (_07374_, \oc8051_golden_model_1.B [3]);
  nor _58810_ (_07375_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and _58811_ (_07376_, _07375_, _07335_);
  and _58812_ (_07377_, _07376_, _07374_);
  and _58813_ (_07378_, \oc8051_golden_model_1.B [2], _05834_);
  not _58814_ (_07379_, _07378_);
  and _58815_ (_07380_, _07379_, _07377_);
  not _58816_ (_07381_, _07380_);
  nor _58817_ (_07382_, _07381_, _07373_);
  nor _58818_ (_07383_, _07382_, _07354_);
  nor _58819_ (_07384_, _07383_, _07343_);
  and _58820_ (_07385_, _07376_, \oc8051_golden_model_1.ACC [7]);
  nor _58821_ (_07386_, _07385_, _07377_);
  nor _58822_ (_07387_, _07384_, \oc8051_golden_model_1.B [3]);
  not _58823_ (_07388_, \oc8051_golden_model_1.B [2]);
  nor _58824_ (_07389_, _07368_, _07359_);
  nor _58825_ (_07390_, _07389_, _07369_);
  not _58826_ (_07391_, _07390_);
  and _58827_ (_07392_, _07391_, _07382_);
  nor _58828_ (_07393_, _07382_, _07356_);
  nor _58829_ (_07394_, _07393_, _07392_);
  and _58830_ (_07395_, _07394_, _07388_);
  nor _58831_ (_07396_, _07394_, _07388_);
  nor _58832_ (_07397_, _07396_, _07395_);
  not _58833_ (_07398_, _07397_);
  not _58834_ (_07399_, \oc8051_golden_model_1.ACC [5]);
  nor _58835_ (_07400_, _07382_, _07399_);
  and _58836_ (_07401_, _07382_, _07361_);
  or _58837_ (_07402_, _07401_, _07400_);
  and _58838_ (_07403_, _07402_, _07334_);
  nor _58839_ (_07404_, _07402_, _07334_);
  not _58840_ (_07405_, \oc8051_golden_model_1.ACC [4]);
  and _58841_ (_07406_, \oc8051_golden_model_1.B [0], _07405_);
  nor _58842_ (_07407_, _07406_, _07404_);
  nor _58843_ (_07408_, _07407_, _07403_);
  nor _58844_ (_07409_, _07408_, _07398_);
  or _58845_ (_07410_, _07409_, _07395_);
  nor _58846_ (_07411_, _07410_, _07387_);
  nor _58847_ (_07412_, _07411_, _07386_);
  nor _58848_ (_07413_, _07412_, _07384_);
  nor _58849_ (_07414_, _07413_, _07343_);
  not _58850_ (_07415_, _07412_);
  and _58851_ (_07416_, _07408_, _07398_);
  nor _58852_ (_07417_, _07416_, _07409_);
  nor _58853_ (_07418_, _07417_, _07415_);
  nor _58854_ (_07419_, _07412_, _07394_);
  nor _58855_ (_07420_, _07419_, _07418_);
  and _58856_ (_07421_, _07420_, _07374_);
  nor _58857_ (_07422_, _07420_, _07374_);
  nor _58858_ (_07423_, _07422_, _07421_);
  not _58859_ (_07424_, _07423_);
  nor _58860_ (_07425_, _07412_, _07402_);
  nor _58861_ (_07426_, _07404_, _07403_);
  and _58862_ (_07427_, _07426_, _07406_);
  nor _58863_ (_07428_, _07426_, _07406_);
  nor _58864_ (_07429_, _07428_, _07427_);
  and _58865_ (_07430_, _07429_, _07412_);
  or _58866_ (_07431_, _07430_, _07425_);
  nor _58867_ (_07432_, _07431_, \oc8051_golden_model_1.B [2]);
  and _58868_ (_07433_, _07431_, \oc8051_golden_model_1.B [2]);
  nor _58869_ (_07434_, _07412_, _07405_);
  nor _58870_ (_07435_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor _58871_ (_07436_, _07435_, _07131_);
  and _58872_ (_07437_, _07412_, _07436_);
  or _58873_ (_07438_, _07437_, _07434_);
  and _58874_ (_07439_, _07438_, _07334_);
  nor _58875_ (_07440_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor _58876_ (_07441_, _07440_, _07189_);
  nor _58877_ (_07442_, _07441_, \oc8051_golden_model_1.ACC [2]);
  nor _58878_ (_07443_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and _58879_ (_07444_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor _58880_ (_07445_, _07444_, _07340_);
  nor _58881_ (_07446_, _07445_, _07443_);
  nor _58882_ (_07447_, _07446_, _07442_);
  not _58883_ (_07448_, _07447_);
  nor _58884_ (_07449_, _07438_, _07334_);
  nor _58885_ (_07450_, _07449_, _07439_);
  and _58886_ (_07451_, _07450_, _07448_);
  nor _58887_ (_07452_, _07451_, _07439_);
  nor _58888_ (_07453_, _07452_, _07433_);
  nor _58889_ (_07454_, _07453_, _07432_);
  nor _58890_ (_07455_, _07454_, _07424_);
  nor _58891_ (_07456_, _07414_, \oc8051_golden_model_1.B [4]);
  nor _58892_ (_07457_, _07456_, _07421_);
  not _58893_ (_07458_, _07457_);
  nor _58894_ (_07459_, _07458_, _07455_);
  not _58895_ (_07460_, \oc8051_golden_model_1.B [5]);
  and _58896_ (_07461_, _07375_, _07460_);
  not _58897_ (_07462_, _07461_);
  and _58898_ (_07463_, \oc8051_golden_model_1.B [4], _05834_);
  nor _58899_ (_07464_, _07463_, _07462_);
  not _58900_ (_07465_, _07464_);
  nor _58901_ (_07466_, _07465_, _07459_);
  nor _58902_ (_07467_, _07466_, _07414_);
  nor _58903_ (_07468_, _07467_, _07343_);
  and _58904_ (_07469_, _07375_, \oc8051_golden_model_1.ACC [7]);
  nor _58905_ (_07470_, _07469_, _07461_);
  nor _58906_ (_07471_, _07468_, \oc8051_golden_model_1.B [5]);
  not _58907_ (_07472_, \oc8051_golden_model_1.B [4]);
  and _58908_ (_07473_, _07454_, _07424_);
  nor _58909_ (_07474_, _07473_, _07455_);
  not _58910_ (_07475_, _07474_);
  and _58911_ (_07476_, _07475_, _07466_);
  nor _58912_ (_07477_, _07466_, _07420_);
  nor _58913_ (_07478_, _07477_, _07476_);
  and _58914_ (_07479_, _07478_, _07472_);
  nor _58915_ (_07480_, _07478_, _07472_);
  nor _58916_ (_07481_, _07480_, _07479_);
  not _58917_ (_07482_, _07481_);
  nor _58918_ (_07483_, _07466_, _07431_);
  nor _58919_ (_07484_, _07433_, _07432_);
  and _58920_ (_07485_, _07484_, _07452_);
  nor _58921_ (_07486_, _07484_, _07452_);
  nor _58922_ (_07487_, _07486_, _07485_);
  not _58923_ (_07488_, _07487_);
  and _58924_ (_07489_, _07488_, _07466_);
  nor _58925_ (_07490_, _07489_, _07483_);
  nor _58926_ (_07491_, _07490_, \oc8051_golden_model_1.B [3]);
  and _58927_ (_07492_, _07490_, \oc8051_golden_model_1.B [3]);
  nor _58928_ (_07493_, _07450_, _07448_);
  nor _58929_ (_07494_, _07493_, _07451_);
  not _58930_ (_07495_, _07494_);
  and _58931_ (_07496_, _07495_, _07466_);
  nor _58932_ (_07497_, _07466_, _07438_);
  nor _58933_ (_07498_, _07497_, _07496_);
  and _58934_ (_07499_, _07498_, _07388_);
  not _58935_ (_07500_, \oc8051_golden_model_1.ACC [3]);
  nor _58936_ (_07501_, _07466_, _07500_);
  and _58937_ (_07502_, _07466_, _07441_);
  or _58938_ (_07503_, _07502_, _07501_);
  and _58939_ (_07504_, _07503_, _07334_);
  nor _58940_ (_07505_, _07503_, _07334_);
  not _58941_ (_07506_, \oc8051_golden_model_1.ACC [2]);
  and _58942_ (_07507_, \oc8051_golden_model_1.B [0], _07506_);
  nor _58943_ (_07508_, _07507_, _07505_);
  nor _58944_ (_07509_, _07508_, _07504_);
  nor _58945_ (_07510_, _07498_, _07388_);
  nor _58946_ (_07511_, _07510_, _07499_);
  not _58947_ (_07512_, _07511_);
  nor _58948_ (_07513_, _07512_, _07509_);
  nor _58949_ (_07514_, _07513_, _07499_);
  nor _58950_ (_07515_, _07514_, _07492_);
  nor _58951_ (_07516_, _07515_, _07491_);
  nor _58952_ (_07517_, _07516_, _07482_);
  or _58953_ (_07518_, _07517_, _07479_);
  nor _58954_ (_07519_, _07518_, _07471_);
  nor _58955_ (_07520_, _07519_, _07470_);
  nor _58956_ (_07521_, _07520_, _07468_);
  not _58957_ (_07522_, _07520_);
  and _58958_ (_07523_, _07516_, _07482_);
  nor _58959_ (_07524_, _07523_, _07517_);
  nor _58960_ (_07525_, _07524_, _07522_);
  nor _58961_ (_07526_, _07520_, _07478_);
  nor _58962_ (_07527_, _07526_, _07525_);
  and _58963_ (_07528_, _07527_, _07460_);
  nor _58964_ (_07529_, _07527_, _07460_);
  nor _58965_ (_07530_, _07529_, _07528_);
  not _58966_ (_07531_, _07530_);
  nor _58967_ (_07532_, _07520_, _07490_);
  nor _58968_ (_07533_, _07492_, _07491_);
  nor _58969_ (_07534_, _07533_, _07514_);
  and _58970_ (_07535_, _07533_, _07514_);
  or _58971_ (_07536_, _07535_, _07534_);
  and _58972_ (_07537_, _07536_, _07520_);
  or _58973_ (_07538_, _07537_, _07532_);
  and _58974_ (_07539_, _07538_, _07472_);
  nor _58975_ (_07540_, _07538_, _07472_);
  and _58976_ (_07541_, _07512_, _07509_);
  nor _58977_ (_07542_, _07541_, _07513_);
  nor _58978_ (_07543_, _07542_, _07522_);
  nor _58979_ (_07544_, _07520_, _07498_);
  nor _58980_ (_07545_, _07544_, _07543_);
  and _58981_ (_07546_, _07545_, _07374_);
  nor _58982_ (_07547_, _07505_, _07504_);
  nor _58983_ (_07548_, _07547_, _07507_);
  and _58984_ (_07549_, _07547_, _07507_);
  or _58985_ (_07550_, _07549_, _07548_);
  nor _58986_ (_07551_, _07550_, _07522_);
  nor _58987_ (_07552_, _07520_, _07503_);
  nor _58988_ (_07553_, _07552_, _07551_);
  and _58989_ (_07554_, _07553_, _07388_);
  nor _58990_ (_07555_, _07553_, _07388_);
  nor _58991_ (_07556_, _07520_, _07506_);
  nor _58992_ (_07557_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor _58993_ (_07558_, _07557_, _07234_);
  and _58994_ (_07559_, _07520_, _07558_);
  or _58995_ (_07560_, _07559_, _07556_);
  and _58996_ (_07561_, _07560_, _07334_);
  and _58997_ (_07562_, \oc8051_golden_model_1.B [0], _03233_);
  not _58998_ (_07563_, _07562_);
  nor _58999_ (_07564_, _07560_, _07334_);
  nor _59000_ (_07565_, _07564_, _07561_);
  and _59001_ (_07566_, _07565_, _07563_);
  nor _59002_ (_07567_, _07566_, _07561_);
  nor _59003_ (_07568_, _07567_, _07555_);
  nor _59004_ (_07569_, _07568_, _07554_);
  nor _59005_ (_07570_, _07545_, _07374_);
  nor _59006_ (_07571_, _07570_, _07546_);
  not _59007_ (_07572_, _07571_);
  nor _59008_ (_07573_, _07572_, _07569_);
  nor _59009_ (_07574_, _07573_, _07546_);
  nor _59010_ (_07575_, _07574_, _07540_);
  nor _59011_ (_07576_, _07575_, _07539_);
  nor _59012_ (_07577_, _07576_, _07531_);
  nor _59013_ (_07578_, _07577_, _07528_);
  and _59014_ (_07579_, _06759_, \oc8051_golden_model_1.ACC [7]);
  nor _59015_ (_07580_, _07579_, _07375_);
  nor _59016_ (_07581_, _07580_, _07578_);
  not _59017_ (_07582_, _07375_);
  nor _59018_ (_07583_, _07521_, _07343_);
  nor _59019_ (_07584_, _07583_, _07582_);
  nor _59020_ (_07585_, _07584_, _07581_);
  and _59021_ (_07586_, _07585_, _07521_);
  nor _59022_ (_07587_, _07586_, _07343_);
  and _59023_ (_07588_, _07587_, \oc8051_golden_model_1.B [7]);
  and _59024_ (_07589_, _07587_, _06759_);
  nor _59025_ (_07590_, _07589_, _06870_);
  not _59026_ (_07591_, _07590_);
  not _59027_ (_07592_, \oc8051_golden_model_1.B [6]);
  and _59028_ (_07593_, _07576_, _07531_);
  nor _59029_ (_07594_, _07593_, _07577_);
  nor _59030_ (_07595_, _07594_, _07585_);
  not _59031_ (_07596_, _07585_);
  nor _59032_ (_07597_, _07596_, _07527_);
  nor _59033_ (_07598_, _07597_, _07595_);
  nor _59034_ (_07599_, _07598_, _07592_);
  and _59035_ (_07600_, _07598_, _07592_);
  nor _59036_ (_07601_, _07540_, _07539_);
  nor _59037_ (_07602_, _07601_, _07574_);
  and _59038_ (_07603_, _07601_, _07574_);
  or _59039_ (_07604_, _07603_, _07602_);
  nor _59040_ (_07605_, _07604_, _07585_);
  nor _59041_ (_07606_, _07596_, _07538_);
  nor _59042_ (_07607_, _07606_, _07605_);
  nor _59043_ (_07608_, _07607_, _07460_);
  and _59044_ (_07609_, _07607_, _07460_);
  not _59045_ (_07610_, _07609_);
  and _59046_ (_07611_, _07572_, _07569_);
  nor _59047_ (_07612_, _07611_, _07573_);
  nor _59048_ (_07613_, _07612_, _07585_);
  nor _59049_ (_07614_, _07596_, _07545_);
  nor _59050_ (_07615_, _07614_, _07613_);
  nor _59051_ (_07616_, _07615_, _07472_);
  and _59052_ (_07617_, _07585_, _07553_);
  nor _59053_ (_07618_, _07555_, _07554_);
  and _59054_ (_07619_, _07618_, _07567_);
  nor _59055_ (_07620_, _07618_, _07567_);
  nor _59056_ (_07621_, _07620_, _07619_);
  nor _59057_ (_07622_, _07621_, _07585_);
  or _59058_ (_07623_, _07622_, _07617_);
  and _59059_ (_07624_, _07623_, _07374_);
  nor _59060_ (_07625_, _07623_, _07374_);
  nor _59061_ (_07626_, _07625_, _07624_);
  nor _59062_ (_07627_, _07565_, _07563_);
  nor _59063_ (_07628_, _07627_, _07566_);
  nor _59064_ (_07629_, _07628_, _07585_);
  nor _59065_ (_07630_, _07596_, _07560_);
  nor _59066_ (_07631_, _07630_, _07629_);
  nor _59067_ (_07632_, _07631_, _07388_);
  and _59068_ (_07633_, _07631_, _07388_);
  nor _59069_ (_07634_, _07633_, _07632_);
  and _59070_ (_07635_, _07634_, _07626_);
  and _59071_ (_07636_, _07585_, _03233_);
  and _59072_ (_07637_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor _59073_ (_07638_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor _59074_ (_07639_, _07638_, _07637_);
  nor _59075_ (_07640_, _07585_, _07639_);
  nor _59076_ (_07641_, _07640_, _07636_);
  and _59077_ (_07642_, _07641_, _07334_);
  nor _59078_ (_07643_, _07641_, _07334_);
  and _59079_ (_07644_, _07340_, \oc8051_golden_model_1.ACC [0]);
  not _59080_ (_07645_, _07644_);
  nor _59081_ (_07646_, _07645_, _07643_);
  nor _59082_ (_07647_, _07646_, _07642_);
  and _59083_ (_07648_, _07647_, _07635_);
  and _59084_ (_07649_, _07632_, _07626_);
  nor _59085_ (_07650_, _07649_, _07625_);
  not _59086_ (_07651_, _07650_);
  nor _59087_ (_07652_, _07651_, _07648_);
  and _59088_ (_07653_, _07615_, _07472_);
  nor _59089_ (_07654_, _07653_, _07652_);
  or _59090_ (_07655_, _07654_, _07616_);
  and _59091_ (_07656_, _07655_, _07610_);
  nor _59092_ (_07657_, _07656_, _07608_);
  nor _59093_ (_07658_, _07657_, _07600_);
  or _59094_ (_07659_, _07658_, _07599_);
  and _59095_ (_07660_, _07659_, _07591_);
  nor _59096_ (_07661_, _07660_, _07588_);
  nor _59097_ (_07662_, _07653_, _07616_);
  nor _59098_ (_07663_, _07609_, _07608_);
  and _59099_ (_07664_, _07663_, _07662_);
  nor _59100_ (_07665_, _07600_, _07599_);
  and _59101_ (_07666_, _07665_, _07591_);
  and _59102_ (_07667_, _07666_, _07664_);
  and _59103_ (_07668_, \oc8051_golden_model_1.B [0], _03321_);
  not _59104_ (_07669_, _07668_);
  nor _59105_ (_07670_, _07643_, _07642_);
  and _59106_ (_07671_, _07670_, _07669_);
  and _59107_ (_07672_, _07671_, _07645_);
  and _59108_ (_07673_, _07672_, _07635_);
  and _59109_ (_07674_, _07673_, _07667_);
  nor _59110_ (_07675_, _07674_, _07661_);
  and _59111_ (_07676_, _07675_, _07586_);
  not _59112_ (_07677_, _07328_);
  or _59113_ (_07678_, _07343_, _07677_);
  or _59114_ (_07679_, _07678_, _07676_);
  and _59115_ (_07680_, _07679_, _07333_);
  or _59116_ (_07681_, _07680_, _03437_);
  and _59117_ (_07682_, _06087_, _05221_);
  or _59118_ (_07683_, _07682_, _06761_);
  or _59119_ (_07684_, _07683_, _03438_);
  and _59120_ (_07685_, _07684_, _04499_);
  and _59121_ (_07686_, _07685_, _07681_);
  and _59122_ (_07687_, _06305_, _05221_);
  or _59123_ (_07688_, _07687_, _06761_);
  and _59124_ (_07689_, _07688_, _03636_);
  or _59125_ (_07690_, _07689_, _03769_);
  or _59126_ (_07691_, _07690_, _07686_);
  and _59127_ (_07692_, _06311_, _05221_);
  or _59128_ (_07693_, _07692_, _06761_);
  or _59129_ (_07694_, _07693_, _04501_);
  and _59130_ (_07695_, _07694_, _05769_);
  and _59131_ (_07696_, _07695_, _07691_);
  or _59132_ (_07697_, _06761_, _05282_);
  and _59133_ (_07698_, _07697_, _03754_);
  and _59134_ (_07699_, _07698_, _07683_);
  or _59135_ (_07700_, _07699_, _07696_);
  and _59136_ (_07701_, _07700_, _03753_);
  and _59137_ (_07702_, _06774_, _03752_);
  and _59138_ (_07703_, _07702_, _07697_);
  or _59139_ (_07704_, _07703_, _03758_);
  or _59140_ (_07705_, _07704_, _07701_);
  nor _59141_ (_07706_, _06304_, _06762_);
  or _59142_ (_07707_, _06761_, _03759_);
  or _59143_ (_07708_, _07707_, _07706_);
  and _59144_ (_07709_, _07708_, _04517_);
  and _59145_ (_07710_, _07709_, _07705_);
  nor _59146_ (_07711_, _06310_, _06762_);
  or _59147_ (_07712_, _07711_, _06761_);
  and _59148_ (_07713_, _07712_, _03760_);
  or _59149_ (_07714_, _07713_, _03790_);
  or _59150_ (_07715_, _07714_, _07710_);
  or _59151_ (_07716_, _06771_, _04192_);
  and _59152_ (_07717_, _07716_, _03152_);
  and _59153_ (_07718_, _07717_, _07715_);
  and _59154_ (_07719_, _06768_, _03151_);
  or _59155_ (_07720_, _07719_, _03520_);
  or _59156_ (_07721_, _07720_, _07718_);
  and _59157_ (_07722_, _05767_, _05221_);
  or _59158_ (_07723_, _06761_, _03521_);
  or _59159_ (_07724_, _07723_, _07722_);
  and _59160_ (_07725_, _07724_, _42963_);
  and _59161_ (_07726_, _07725_, _07721_);
  or _59162_ (_07727_, _07726_, _06760_);
  and _59163_ (_40515_, _07727_, _41755_);
  nor _59164_ (_07728_, _42963_, _05834_);
  and _59165_ (_07729_, _03230_, _03171_);
  nand _59166_ (_07730_, _07729_, _07346_);
  and _59167_ (_07731_, _03478_, _03171_);
  not _59168_ (_07732_, _07731_);
  and _59169_ (_07733_, _06004_, _05834_);
  and _59170_ (_07734_, _05935_, \oc8051_golden_model_1.ACC [7]);
  nor _59171_ (_07735_, _07734_, _07733_);
  and _59172_ (_07736_, _06713_, \oc8051_golden_model_1.ACC [6]);
  and _59173_ (_07737_, _06388_, _07346_);
  nor _59174_ (_07738_, _07737_, _07736_);
  and _59175_ (_07739_, _06721_, \oc8051_golden_model_1.ACC [5]);
  and _59176_ (_07740_, _06616_, _07399_);
  nor _59177_ (_07741_, _07740_, _07739_);
  not _59178_ (_07742_, _07741_);
  and _59179_ (_07743_, _06722_, \oc8051_golden_model_1.ACC [4]);
  and _59180_ (_07744_, _06661_, _07405_);
  nor _59181_ (_07745_, _07744_, _07743_);
  and _59182_ (_07746_, _06524_, _07500_);
  not _59183_ (_07747_, _07746_);
  and _59184_ (_07748_, _06717_, \oc8051_golden_model_1.ACC [3]);
  not _59185_ (_07749_, _07748_);
  and _59186_ (_07750_, _06718_, \oc8051_golden_model_1.ACC [2]);
  and _59187_ (_07751_, _06569_, _07506_);
  nor _59188_ (_07752_, _07751_, _07750_);
  not _59189_ (_07753_, _07752_);
  and _59190_ (_07754_, _06714_, \oc8051_golden_model_1.ACC [1]);
  and _59191_ (_07755_, _06433_, _03233_);
  nor _59192_ (_07756_, _07755_, _07754_);
  and _59193_ (_07757_, _06715_, \oc8051_golden_model_1.ACC [0]);
  and _59194_ (_07758_, _07757_, _07756_);
  nor _59195_ (_07759_, _07758_, _07754_);
  nor _59196_ (_07760_, _07759_, _07753_);
  nor _59197_ (_07761_, _07760_, _07750_);
  nand _59198_ (_07762_, _07761_, _07749_);
  and _59199_ (_07763_, _07762_, _07747_);
  and _59200_ (_07764_, _07763_, _07745_);
  nor _59201_ (_07765_, _07764_, _07743_);
  nor _59202_ (_07766_, _07765_, _07742_);
  or _59203_ (_07767_, _07766_, _07739_);
  and _59204_ (_07768_, _07767_, _07738_);
  nor _59205_ (_07769_, _07768_, _07736_);
  nor _59206_ (_07770_, _07769_, _07735_);
  and _59207_ (_07771_, _07769_, _07735_);
  or _59208_ (_07772_, _07771_, _07770_);
  or _59209_ (_07773_, _07772_, _07732_);
  and _59210_ (_07774_, _03476_, _03171_);
  not _59211_ (_07775_, _07774_);
  not _59212_ (_07776_, _03662_);
  nor _59213_ (_07777_, _07776_, _03484_);
  and _59214_ (_07778_, _07777_, _04002_);
  or _59215_ (_07779_, _07778_, _04178_);
  and _59216_ (_07780_, _07779_, _07775_);
  and _59217_ (_07781_, _03650_, _03171_);
  nor _59218_ (_07782_, _05176_, _05834_);
  and _59219_ (_07783_, _05176_, _05834_);
  nor _59220_ (_07784_, _07783_, _07782_);
  nor _59221_ (_07785_, _05327_, _07346_);
  and _59222_ (_07786_, _05327_, _07346_);
  nor _59223_ (_07787_, _07786_, _07785_);
  and _59224_ (_07788_, _05422_, _07399_);
  not _59225_ (_07789_, _07788_);
  nor _59226_ (_07790_, _05422_, _07399_);
  not _59227_ (_07791_, _07790_);
  nor _59228_ (_07792_, _05712_, _07405_);
  and _59229_ (_07793_, _05712_, _07405_);
  nor _59230_ (_07794_, _07793_, _07792_);
  and _59231_ (_07795_, _04843_, _07500_);
  not _59232_ (_07796_, _07795_);
  nor _59233_ (_07797_, _04843_, _07500_);
  not _59234_ (_07798_, _07797_);
  nor _59235_ (_07799_, _05026_, _07506_);
  and _59236_ (_07800_, _05026_, _07506_);
  nor _59237_ (_07801_, _07800_, _07799_);
  not _59238_ (_07802_, _07801_);
  nor _59239_ (_07803_, _04603_, _03233_);
  and _59240_ (_07804_, _04603_, _03233_);
  nor _59241_ (_07805_, _07804_, _07803_);
  and _59242_ (_07806_, _04419_, \oc8051_golden_model_1.ACC [0]);
  and _59243_ (_07807_, _07806_, _07805_);
  nor _59244_ (_07808_, _07807_, _07803_);
  nor _59245_ (_07809_, _07808_, _07802_);
  nor _59246_ (_07810_, _07809_, _07799_);
  nand _59247_ (_07811_, _07810_, _07798_);
  and _59248_ (_07812_, _07811_, _07796_);
  and _59249_ (_07813_, _07812_, _07794_);
  nor _59250_ (_07814_, _07813_, _07792_);
  nand _59251_ (_07815_, _07814_, _07791_);
  and _59252_ (_07816_, _07815_, _07789_);
  and _59253_ (_07817_, _07816_, _07787_);
  nor _59254_ (_07818_, _07817_, _07785_);
  nor _59255_ (_07819_, _07818_, _07784_);
  and _59256_ (_07820_, _07818_, _07784_);
  or _59257_ (_07821_, _07820_, _07819_);
  not _59258_ (_07822_, _07821_);
  nor _59259_ (_07823_, _07822_, _07781_);
  or _59260_ (_07824_, _07823_, _07780_);
  and _59261_ (_07825_, _03478_, _03177_);
  or _59262_ (_07826_, _07777_, _04156_);
  nand _59263_ (_07827_, _03475_, _03228_);
  nor _59264_ (_07828_, _07827_, _04156_);
  not _59265_ (_07829_, _07828_);
  and _59266_ (_07830_, _07829_, _07826_);
  not _59267_ (_07831_, _05327_);
  and _59268_ (_07832_, _06697_, \oc8051_golden_model_1.PSW [7]);
  and _59269_ (_07833_, _07832_, _07831_);
  nor _59270_ (_07834_, _07833_, _05176_);
  and _59271_ (_07835_, _07833_, _05176_);
  nor _59272_ (_07836_, _07835_, _07834_);
  and _59273_ (_07837_, _07836_, \oc8051_golden_model_1.ACC [7]);
  nor _59274_ (_07838_, _07836_, \oc8051_golden_model_1.ACC [7]);
  nor _59275_ (_07839_, _07838_, _07837_);
  nor _59276_ (_07840_, _07832_, _07831_);
  nor _59277_ (_07841_, _07840_, _07833_);
  and _59278_ (_07842_, _07841_, \oc8051_golden_model_1.ACC [6]);
  and _59279_ (_07843_, _07841_, _07346_);
  nor _59280_ (_07844_, _07841_, _07346_);
  nor _59281_ (_07845_, _07844_, _07843_);
  not _59282_ (_07846_, _07845_);
  not _59283_ (_07847_, _05422_);
  not _59284_ (_07848_, _05712_);
  and _59285_ (_07849_, _06692_, \oc8051_golden_model_1.PSW [7]);
  and _59286_ (_07850_, _07849_, _06693_);
  and _59287_ (_07851_, _07850_, _07848_);
  nor _59288_ (_07852_, _07851_, _07847_);
  nor _59289_ (_07853_, _07852_, _07832_);
  and _59290_ (_07854_, _07853_, \oc8051_golden_model_1.ACC [5]);
  and _59291_ (_07855_, _07853_, _07399_);
  nor _59292_ (_07856_, _07853_, _07399_);
  nor _59293_ (_07857_, _07856_, _07855_);
  nor _59294_ (_07858_, _07850_, _07848_);
  nor _59295_ (_07859_, _07858_, _07851_);
  and _59296_ (_07860_, _07859_, \oc8051_golden_model_1.ACC [4]);
  nor _59297_ (_07861_, _07859_, _07405_);
  and _59298_ (_07862_, _07859_, _07405_);
  or _59299_ (_07863_, _07862_, _07861_);
  not _59300_ (_07864_, _04843_);
  not _59301_ (_07865_, _05026_);
  and _59302_ (_07866_, _06692_, _07865_);
  and _59303_ (_07867_, _07866_, \oc8051_golden_model_1.PSW [7]);
  nor _59304_ (_07868_, _07867_, _07864_);
  nor _59305_ (_07869_, _07868_, _07850_);
  and _59306_ (_07870_, _07869_, \oc8051_golden_model_1.ACC [3]);
  nor _59307_ (_07871_, _07869_, _07500_);
  and _59308_ (_07872_, _07869_, _07500_);
  nor _59309_ (_07873_, _07872_, _07871_);
  nor _59310_ (_07874_, _07849_, _07865_);
  nor _59311_ (_07875_, _07874_, _07867_);
  and _59312_ (_07876_, _07875_, \oc8051_golden_model_1.ACC [2]);
  nor _59313_ (_07877_, _07875_, _07506_);
  and _59314_ (_07878_, _07875_, _07506_);
  nor _59315_ (_07879_, _07878_, _07877_);
  not _59316_ (_07880_, _04603_);
  and _59317_ (_07881_, _04419_, \oc8051_golden_model_1.PSW [7]);
  nor _59318_ (_07882_, _07881_, _07880_);
  nor _59319_ (_07883_, _07882_, _07849_);
  and _59320_ (_07884_, _07883_, \oc8051_golden_model_1.ACC [1]);
  nor _59321_ (_07885_, _07883_, _03233_);
  and _59322_ (_07886_, _07883_, _03233_);
  nor _59323_ (_07887_, _07886_, _07885_);
  not _59324_ (_07888_, \oc8051_golden_model_1.PSW [7]);
  and _59325_ (_07889_, _04439_, _07888_);
  nor _59326_ (_07890_, _07889_, _07881_);
  and _59327_ (_07891_, _07890_, \oc8051_golden_model_1.ACC [0]);
  not _59328_ (_07892_, _07891_);
  nor _59329_ (_07893_, _07892_, _07887_);
  nor _59330_ (_07894_, _07893_, _07884_);
  nor _59331_ (_07895_, _07894_, _07879_);
  nor _59332_ (_07896_, _07895_, _07876_);
  nor _59333_ (_07897_, _07896_, _07873_);
  or _59334_ (_07898_, _07897_, _07870_);
  and _59335_ (_07899_, _07898_, _07863_);
  nor _59336_ (_07900_, _07899_, _07860_);
  nor _59337_ (_07901_, _07900_, _07857_);
  or _59338_ (_07902_, _07901_, _07854_);
  and _59339_ (_07903_, _07902_, _07846_);
  nor _59340_ (_07904_, _07903_, _07842_);
  nor _59341_ (_07905_, _07904_, _07839_);
  and _59342_ (_07906_, _07904_, _07839_);
  nor _59343_ (_07907_, _07906_, _07905_);
  or _59344_ (_07908_, _07907_, _07830_);
  and _59345_ (_07909_, _03637_, _03191_);
  not _59346_ (_07910_, _07909_);
  not _59347_ (_07911_, _03755_);
  or _59348_ (_07912_, _06309_, _07911_);
  and _59349_ (_07913_, _07912_, _07910_);
  and _59350_ (_07914_, _07782_, _04135_);
  nor _59351_ (_07915_, _05227_, _05834_);
  and _59352_ (_07916_, _07915_, _03769_);
  or _59353_ (_07917_, _03401_, _03232_);
  not _59354_ (_07918_, _05227_);
  nor _59355_ (_07919_, _07918_, _05176_);
  nor _59356_ (_07920_, _07919_, _07915_);
  nand _59357_ (_07921_, _07920_, _07314_);
  nand _59358_ (_07922_, _03222_, _03147_);
  not _59359_ (_07923_, _07922_);
  not _59360_ (_07924_, _03978_);
  and _59361_ (_07925_, _04711_, _03944_);
  and _59362_ (_07926_, _07925_, _07924_);
  and _59363_ (_07927_, _07926_, _04750_);
  not _59364_ (_07928_, _07927_);
  nand _59365_ (_07929_, _07928_, _05176_);
  or _59366_ (_07930_, _03478_, _03650_);
  nor _59367_ (_07931_, _07930_, _03220_);
  and _59368_ (_07932_, _07931_, _03666_);
  nor _59369_ (_07933_, _07932_, _03207_);
  nand _59370_ (_07934_, _07933_, _05176_);
  and _59371_ (_07935_, _03637_, _03571_);
  not _59372_ (_07936_, _07935_);
  nor _59373_ (_07937_, _04012_, _05834_);
  and _59374_ (_07938_, _04012_, _05834_);
  or _59375_ (_07939_, _07938_, _07937_);
  or _59376_ (_07940_, _07939_, _07933_);
  and _59377_ (_07941_, _07940_, _07936_);
  and _59378_ (_07942_, _07941_, _07934_);
  and _59379_ (_07943_, _07935_, _05935_);
  or _59380_ (_07944_, _07943_, _07942_);
  not _59381_ (_07945_, _03208_);
  nor _59382_ (_07946_, _03570_, _07945_);
  and _59383_ (_07947_, _07946_, _07944_);
  and _59384_ (_07948_, _03637_, _03515_);
  and _59385_ (_07949_, _05949_, _05227_);
  nor _59386_ (_07950_, _07949_, _07915_);
  nor _59387_ (_07951_, _07950_, _04444_);
  or _59388_ (_07952_, _07951_, _07948_);
  or _59389_ (_07953_, _07952_, _07947_);
  nor _59390_ (_07954_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor _59391_ (_07955_, _07954_, _07500_);
  and _59392_ (_07956_, _07955_, _07364_);
  and _59393_ (_07957_, _07956_, \oc8051_golden_model_1.ACC [6]);
  and _59394_ (_07958_, _07957_, \oc8051_golden_model_1.ACC [7]);
  nor _59395_ (_07959_, _07957_, \oc8051_golden_model_1.ACC [7]);
  nor _59396_ (_07960_, _07959_, _07958_);
  and _59397_ (_07961_, _07955_, \oc8051_golden_model_1.ACC [4]);
  nor _59398_ (_07962_, _07961_, \oc8051_golden_model_1.ACC [5]);
  nor _59399_ (_07963_, _07962_, _07956_);
  nor _59400_ (_07964_, _07956_, \oc8051_golden_model_1.ACC [6]);
  nor _59401_ (_07965_, _07964_, _07957_);
  nor _59402_ (_07966_, _07965_, _07963_);
  not _59403_ (_07967_, _07966_);
  and _59404_ (_07968_, _07967_, _07960_);
  nor _59405_ (_07969_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor _59406_ (_07970_, _07969_, _07966_);
  nor _59407_ (_07971_, _07970_, _07960_);
  nor _59408_ (_07972_, _07971_, _07968_);
  not _59409_ (_07973_, _07972_);
  nand _59410_ (_07974_, _07973_, _07948_);
  and _59411_ (_07975_, _07974_, _03576_);
  and _59412_ (_07976_, _07975_, _07953_);
  nor _59413_ (_07977_, _05792_, _05834_);
  and _59414_ (_07978_, _05954_, _05792_);
  nor _59415_ (_07979_, _07978_, _07977_);
  nor _59416_ (_07980_, _07979_, _03517_);
  nor _59417_ (_07981_, _07920_, _03983_);
  or _59418_ (_07982_, _07981_, _07928_);
  or _59419_ (_07983_, _07982_, _07980_);
  or _59420_ (_07984_, _07983_, _07976_);
  and _59421_ (_07985_, _07984_, _07929_);
  or _59422_ (_07986_, _07985_, _04458_);
  not _59423_ (_07987_, _04458_);
  or _59424_ (_07988_, _05935_, _07987_);
  and _59425_ (_07989_, _07988_, _03583_);
  and _59426_ (_07990_, _07989_, _07986_);
  and _59427_ (_07991_, _03637_, _03510_);
  nor _59428_ (_07992_, _05984_, _03583_);
  or _59429_ (_07993_, _07992_, _07991_);
  or _59430_ (_07994_, _07993_, _07990_);
  nand _59431_ (_07995_, _07991_, _07500_);
  and _59432_ (_07996_, _07995_, _07994_);
  or _59433_ (_07997_, _07996_, _03512_);
  and _59434_ (_07998_, _05818_, _05792_);
  nor _59435_ (_07999_, _07998_, _07977_);
  nand _59436_ (_08000_, _07999_, _03512_);
  and _59437_ (_08001_, _08000_, _03506_);
  and _59438_ (_08002_, _08001_, _07997_);
  and _59439_ (_08003_, _07978_, _05989_);
  nor _59440_ (_08004_, _08003_, _07977_);
  nor _59441_ (_08005_, _08004_, _03506_);
  or _59442_ (_08006_, _08005_, _06794_);
  or _59443_ (_08007_, _08006_, _08002_);
  nor _59444_ (_08008_, _07284_, _07282_);
  nor _59445_ (_08009_, _08008_, _07285_);
  or _59446_ (_08010_, _08009_, _06800_);
  and _59447_ (_08011_, _08010_, _08007_);
  or _59448_ (_08012_, _08011_, _07923_);
  not _59449_ (_08013_, _07857_);
  or _59450_ (_08014_, _07863_, _08013_);
  and _59451_ (_08015_, _07879_, _07873_);
  and _59452_ (_08016_, _07890_, _03321_);
  nor _59453_ (_08017_, _08016_, _07886_);
  or _59454_ (_08018_, _08017_, _07885_);
  and _59455_ (_08019_, _08018_, _08015_);
  and _59456_ (_08020_, _07877_, _07873_);
  or _59457_ (_08021_, _08020_, _07871_);
  nor _59458_ (_08022_, _08021_, _08019_);
  nor _59459_ (_08023_, _08022_, _08014_);
  and _59460_ (_08024_, _07861_, _07857_);
  nor _59461_ (_08025_, _08024_, _07856_);
  not _59462_ (_08026_, _08025_);
  nor _59463_ (_08027_, _08026_, _08023_);
  nor _59464_ (_08028_, _07846_, _08027_);
  or _59465_ (_08029_, _08028_, _07844_);
  or _59466_ (_08030_, _08029_, _07839_);
  nand _59467_ (_08031_, _08029_, _07839_);
  and _59468_ (_08032_, _08031_, _08030_);
  or _59469_ (_08033_, _08032_, _07922_);
  and _59470_ (_08034_, _08033_, _08012_);
  and _59471_ (_08035_, _03478_, _03222_);
  or _59472_ (_08036_, _08035_, _08034_);
  not _59473_ (_08037_, _08035_);
  and _59474_ (_08038_, _06725_, \oc8051_golden_model_1.PSW [7]);
  nor _59475_ (_08039_, _08038_, _06004_);
  and _59476_ (_08040_, _08038_, _06004_);
  nor _59477_ (_08041_, _08040_, _08039_);
  and _59478_ (_08042_, _08041_, \oc8051_golden_model_1.ACC [7]);
  nor _59479_ (_08043_, _08041_, \oc8051_golden_model_1.ACC [7]);
  nor _59480_ (_08044_, _08043_, _08042_);
  not _59481_ (_08045_, _08044_);
  and _59482_ (_08046_, _06720_, _06722_);
  and _59483_ (_08047_, _08046_, \oc8051_golden_model_1.PSW [7]);
  and _59484_ (_08048_, _08047_, _06721_);
  nor _59485_ (_08049_, _08048_, _06713_);
  nor _59486_ (_08050_, _08049_, _08038_);
  nor _59487_ (_08051_, _08050_, _07346_);
  nor _59488_ (_08052_, _08047_, _06721_);
  nor _59489_ (_08053_, _08052_, _08048_);
  and _59490_ (_08054_, _08053_, _07399_);
  nor _59491_ (_08055_, _08053_, _07399_);
  and _59492_ (_08056_, _06716_, \oc8051_golden_model_1.PSW [7]);
  and _59493_ (_08057_, _08056_, _06719_);
  nor _59494_ (_08058_, _08057_, _06722_);
  nor _59495_ (_08059_, _08058_, _08047_);
  nor _59496_ (_08060_, _08059_, _07405_);
  nor _59497_ (_08061_, _08060_, _08055_);
  nor _59498_ (_08062_, _08061_, _08054_);
  nor _59499_ (_08063_, _08055_, _08054_);
  not _59500_ (_08064_, _08063_);
  and _59501_ (_08065_, _08059_, _07405_);
  or _59502_ (_08066_, _08065_, _08060_);
  or _59503_ (_08067_, _08066_, _08064_);
  and _59504_ (_08068_, _06716_, _06718_);
  and _59505_ (_08069_, _08068_, \oc8051_golden_model_1.PSW [7]);
  nor _59506_ (_08070_, _08069_, _06717_);
  nor _59507_ (_08071_, _08070_, _08057_);
  nor _59508_ (_08072_, _08071_, _07500_);
  and _59509_ (_08073_, _08071_, _07500_);
  nor _59510_ (_08074_, _08073_, _08072_);
  nor _59511_ (_08075_, _08056_, _06718_);
  nor _59512_ (_08076_, _08075_, _08069_);
  nor _59513_ (_08077_, _08076_, _07506_);
  and _59514_ (_08078_, _08076_, _07506_);
  nor _59515_ (_08079_, _08078_, _08077_);
  and _59516_ (_08080_, _08079_, _08074_);
  and _59517_ (_08081_, _06715_, \oc8051_golden_model_1.PSW [7]);
  nor _59518_ (_08082_, _08081_, _06714_);
  nor _59519_ (_08083_, _08082_, _08056_);
  nor _59520_ (_08084_, _08083_, _03233_);
  and _59521_ (_08085_, _08083_, _03233_);
  and _59522_ (_08086_, _06478_, _07888_);
  nor _59523_ (_08087_, _08086_, _08081_);
  and _59524_ (_08088_, _08087_, _03321_);
  nor _59525_ (_08089_, _08088_, _08085_);
  or _59526_ (_08090_, _08089_, _08084_);
  nand _59527_ (_08091_, _08090_, _08080_);
  and _59528_ (_08092_, _08077_, _08074_);
  nor _59529_ (_08093_, _08092_, _08072_);
  and _59530_ (_08094_, _08093_, _08091_);
  nor _59531_ (_08095_, _08094_, _08067_);
  nor _59532_ (_08096_, _08095_, _08062_);
  and _59533_ (_08097_, _08050_, _07346_);
  nor _59534_ (_08098_, _08051_, _08097_);
  not _59535_ (_08099_, _08098_);
  nor _59536_ (_08100_, _08099_, _08096_);
  or _59537_ (_08101_, _08100_, _08051_);
  and _59538_ (_08102_, _08101_, _08045_);
  nor _59539_ (_08103_, _08101_, _08045_);
  or _59540_ (_08104_, _08103_, _08102_);
  or _59541_ (_08105_, _08104_, _08037_);
  and _59542_ (_08106_, _08105_, _08036_);
  or _59543_ (_08107_, _08106_, _03614_);
  and _59544_ (_08108_, _03637_, _03222_);
  not _59545_ (_08109_, _08108_);
  and _59546_ (_08110_, _05276_, \oc8051_golden_model_1.P0INREG [6]);
  not _59547_ (_08111_, _08110_);
  not _59548_ (_08112_, _05350_);
  and _59549_ (_08113_, _05359_, _08112_);
  and _59550_ (_08114_, _08113_, _08111_);
  and _59551_ (_08115_, _05244_, \oc8051_golden_model_1.P1INREG [6]);
  not _59552_ (_08116_, _08115_);
  and _59553_ (_08117_, _05210_, \oc8051_golden_model_1.P2INREG [6]);
  and _59554_ (_08118_, _05200_, \oc8051_golden_model_1.P3INREG [6]);
  nor _59555_ (_08119_, _08118_, _08117_);
  and _59556_ (_08120_, _08119_, _05366_);
  and _59557_ (_08121_, _08120_, _08116_);
  and _59558_ (_08122_, _08121_, _05364_);
  and _59559_ (_08123_, _08122_, _08114_);
  and _59560_ (_08124_, _08123_, _05348_);
  and _59561_ (_08125_, _08124_, _05328_);
  not _59562_ (_08126_, _08125_);
  not _59563_ (_08127_, _05493_);
  and _59564_ (_08128_, _05517_, _08127_);
  nor _59565_ (_08129_, _05497_, _05494_);
  and _59566_ (_08130_, _08129_, _05505_);
  and _59567_ (_08131_, _05210_, \oc8051_golden_model_1.P2INREG [3]);
  and _59568_ (_08132_, _05200_, \oc8051_golden_model_1.P3INREG [3]);
  nor _59569_ (_08133_, _08132_, _08131_);
  and _59570_ (_08134_, _05244_, \oc8051_golden_model_1.P1INREG [3]);
  and _59571_ (_08135_, _05276_, \oc8051_golden_model_1.P0INREG [3]);
  nor _59572_ (_08136_, _08135_, _08134_);
  and _59573_ (_08137_, _08136_, _08133_);
  and _59574_ (_08138_, _08137_, _08130_);
  and _59575_ (_08139_, _08138_, _08128_);
  and _59576_ (_08140_, _05502_, _05479_);
  and _59577_ (_08141_, _08140_, _05492_);
  and _59578_ (_08142_, _08141_, _08139_);
  and _59579_ (_08143_, _08142_, _05473_);
  not _59580_ (_08144_, _08143_);
  not _59581_ (_08145_, _05623_);
  not _59582_ (_08146_, _05659_);
  and _59583_ (_08147_, _08146_, _05622_);
  and _59584_ (_08148_, _08147_, _08145_);
  nor _59585_ (_08149_, _05627_, _05624_);
  and _59586_ (_08150_, _08149_, _05635_);
  and _59587_ (_08151_, _05210_, \oc8051_golden_model_1.P2INREG [2]);
  and _59588_ (_08152_, _05200_, \oc8051_golden_model_1.P3INREG [2]);
  nor _59589_ (_08153_, _08152_, _08151_);
  and _59590_ (_08154_, _05276_, \oc8051_golden_model_1.P0INREG [2]);
  and _59591_ (_08155_, _05244_, \oc8051_golden_model_1.P1INREG [2]);
  nor _59592_ (_08156_, _08155_, _08154_);
  and _59593_ (_08157_, _08156_, _08153_);
  and _59594_ (_08158_, _08157_, _08150_);
  and _59595_ (_08159_, _08158_, _08148_);
  and _59596_ (_08160_, _05632_, _05647_);
  and _59597_ (_08161_, _08160_, _05657_);
  and _59598_ (_08162_, _08161_, _08159_);
  and _59599_ (_08163_, _08162_, _05619_);
  not _59600_ (_08164_, _08163_);
  and _59601_ (_08165_, _05244_, \oc8051_golden_model_1.P1INREG [1]);
  not _59602_ (_08166_, _08165_);
  and _59603_ (_08167_, _05210_, \oc8051_golden_model_1.P2INREG [1]);
  and _59604_ (_08168_, _05200_, \oc8051_golden_model_1.P3INREG [1]);
  nor _59605_ (_08169_, _08168_, _08167_);
  and _59606_ (_08170_, _08169_, _08166_);
  and _59607_ (_08171_, _08170_, _05555_);
  and _59608_ (_08172_, _05276_, \oc8051_golden_model_1.P0INREG [1]);
  nor _59609_ (_08173_, _08172_, _05564_);
  and _59610_ (_08174_, _08173_, _08171_);
  and _59611_ (_08175_, _08174_, _05548_);
  and _59612_ (_08176_, _08175_, _05542_);
  and _59613_ (_08177_, _08176_, _05522_);
  not _59614_ (_08178_, _08177_);
  and _59615_ (_08179_, _05276_, \oc8051_golden_model_1.P0INREG [0]);
  not _59616_ (_08180_, _08179_);
  and _59617_ (_08181_, _05244_, \oc8051_golden_model_1.P1INREG [0]);
  not _59618_ (_08182_, _08181_);
  and _59619_ (_08183_, _05210_, \oc8051_golden_model_1.P2INREG [0]);
  and _59620_ (_08184_, _05200_, \oc8051_golden_model_1.P3INREG [0]);
  nor _59621_ (_08185_, _08184_, _08183_);
  and _59622_ (_08186_, _08185_, _08182_);
  and _59623_ (_08187_, _08186_, _05577_);
  and _59624_ (_08188_, _08187_, _08180_);
  and _59625_ (_08189_, _08188_, _05597_);
  and _59626_ (_08190_, _08189_, _05615_);
  and _59627_ (_08191_, _08190_, _05570_);
  nor _59628_ (_08192_, _08191_, _07888_);
  and _59629_ (_08193_, _08192_, _08178_);
  and _59630_ (_08194_, _08193_, _08164_);
  and _59631_ (_08195_, _08194_, _08144_);
  and _59632_ (_08196_, _05210_, \oc8051_golden_model_1.P2INREG [5]);
  and _59633_ (_08197_, _05200_, \oc8051_golden_model_1.P3INREG [5]);
  nor _59634_ (_08198_, _08197_, _08196_);
  and _59635_ (_08199_, _05276_, \oc8051_golden_model_1.P0INREG [5]);
  and _59636_ (_08200_, _05244_, \oc8051_golden_model_1.P1INREG [5]);
  nor _59637_ (_08201_, _08200_, _08199_);
  and _59638_ (_08202_, _08201_, _08198_);
  and _59639_ (_08203_, _08202_, _05459_);
  and _59640_ (_08204_, _08203_, _05449_);
  and _59641_ (_08205_, _08204_, _05423_);
  not _59642_ (_08206_, _05723_);
  and _59643_ (_08207_, _05755_, _08206_);
  nor _59644_ (_08208_, _05727_, _05724_);
  and _59645_ (_08209_, _08208_, _05735_);
  and _59646_ (_08210_, _05210_, \oc8051_golden_model_1.P2INREG [4]);
  and _59647_ (_08211_, _05200_, \oc8051_golden_model_1.P3INREG [4]);
  nor _59648_ (_08212_, _08211_, _08210_);
  and _59649_ (_08213_, _05276_, \oc8051_golden_model_1.P0INREG [4]);
  and _59650_ (_08214_, _05244_, \oc8051_golden_model_1.P1INREG [4]);
  nor _59651_ (_08215_, _08214_, _08213_);
  and _59652_ (_08216_, _08215_, _08212_);
  and _59653_ (_08217_, _08216_, _08209_);
  and _59654_ (_08218_, _08217_, _08207_);
  and _59655_ (_08219_, _05732_, _05743_);
  and _59656_ (_08220_, _08219_, _05722_);
  and _59657_ (_08221_, _08220_, _08218_);
  and _59658_ (_08222_, _08221_, _05713_);
  nor _59659_ (_08223_, _08222_, _08205_);
  and _59660_ (_08224_, _08223_, _08195_);
  and _59661_ (_08225_, _08224_, _08126_);
  nor _59662_ (_08226_, _08225_, _05984_);
  and _59663_ (_08227_, _08225_, _05984_);
  nor _59664_ (_08228_, _08227_, _08226_);
  and _59665_ (_08229_, _08228_, \oc8051_golden_model_1.ACC [7]);
  nor _59666_ (_08230_, _08228_, \oc8051_golden_model_1.ACC [7]);
  nor _59667_ (_08231_, _08230_, _08229_);
  nor _59668_ (_08232_, _08224_, _08126_);
  nor _59669_ (_08233_, _08232_, _08225_);
  nor _59670_ (_08234_, _08233_, _07346_);
  not _59671_ (_08235_, _08205_);
  not _59672_ (_08236_, _08222_);
  and _59673_ (_08237_, _08195_, _08236_);
  nor _59674_ (_08238_, _08237_, _08235_);
  nor _59675_ (_08239_, _08238_, _08224_);
  and _59676_ (_08240_, _08239_, _07399_);
  nor _59677_ (_08241_, _08239_, _07399_);
  nor _59678_ (_08242_, _08195_, _08236_);
  nor _59679_ (_08243_, _08242_, _08237_);
  nor _59680_ (_08244_, _08243_, _07405_);
  nor _59681_ (_08245_, _08244_, _08241_);
  nor _59682_ (_08246_, _08245_, _08240_);
  nor _59683_ (_08247_, _08241_, _08240_);
  and _59684_ (_08248_, _08243_, _07405_);
  nor _59685_ (_08249_, _08248_, _08244_);
  and _59686_ (_08250_, _08249_, _08247_);
  not _59687_ (_08251_, _08250_);
  nor _59688_ (_08252_, _08194_, _08144_);
  nor _59689_ (_08253_, _08252_, _08195_);
  nor _59690_ (_08254_, _08253_, _07500_);
  and _59691_ (_08255_, _08253_, _07500_);
  nor _59692_ (_08256_, _08255_, _08254_);
  nor _59693_ (_08257_, _08193_, _08164_);
  nor _59694_ (_08258_, _08257_, _08194_);
  nor _59695_ (_08259_, _08258_, _07506_);
  and _59696_ (_08260_, _08258_, _07506_);
  nor _59697_ (_08261_, _08260_, _08259_);
  and _59698_ (_08262_, _08261_, _08256_);
  nor _59699_ (_08263_, _08192_, _08178_);
  nor _59700_ (_08264_, _08263_, _08193_);
  nor _59701_ (_08265_, _08264_, _03233_);
  and _59702_ (_08266_, _08264_, _03233_);
  and _59703_ (_08267_, _08191_, _07888_);
  nor _59704_ (_08268_, _08267_, _08192_);
  and _59705_ (_08269_, _08268_, _03321_);
  nor _59706_ (_08270_, _08269_, _08266_);
  or _59707_ (_08271_, _08270_, _08265_);
  nand _59708_ (_08272_, _08271_, _08262_);
  nor _59709_ (_08273_, _08259_, _08254_);
  or _59710_ (_08274_, _08273_, _08255_);
  and _59711_ (_08275_, _08274_, _08272_);
  nor _59712_ (_08276_, _08275_, _08251_);
  or _59713_ (_08277_, _08276_, _08246_);
  and _59714_ (_08278_, _08233_, _07346_);
  nor _59715_ (_08279_, _08234_, _08278_);
  and _59716_ (_08280_, _08279_, _08277_);
  nor _59717_ (_08281_, _08280_, _08234_);
  or _59718_ (_08282_, _08281_, _08231_);
  nand _59719_ (_08283_, _08281_, _08231_);
  and _59720_ (_08284_, _08283_, _08282_);
  nand _59721_ (_08285_, _08284_, _03614_);
  and _59722_ (_08286_, _08285_, _08109_);
  and _59723_ (_08287_, _08286_, _08107_);
  and _59724_ (_08288_, _05206_, \oc8051_golden_model_1.PSW [7]);
  and _59725_ (_08289_, _08288_, _05232_);
  and _59726_ (_08290_, _08289_, _05198_);
  and _59727_ (_08291_, _08290_, _04956_);
  nor _59728_ (_08292_, _08291_, _05215_);
  and _59729_ (_08293_, _08291_, _05215_);
  nor _59730_ (_08294_, _08293_, _08292_);
  and _59731_ (_08295_, _08294_, \oc8051_golden_model_1.ACC [7]);
  nor _59732_ (_08296_, _08294_, \oc8051_golden_model_1.ACC [7]);
  nor _59733_ (_08297_, _08296_, _08295_);
  not _59734_ (_08298_, _08297_);
  nor _59735_ (_08299_, _08290_, _04956_);
  nor _59736_ (_08300_, _08299_, _08291_);
  nor _59737_ (_08301_, _08300_, _07346_);
  and _59738_ (_08302_, _08289_, _05182_);
  nor _59739_ (_08303_, _08302_, _05190_);
  nor _59740_ (_08304_, _08303_, _08290_);
  and _59741_ (_08305_, _08304_, _07399_);
  nor _59742_ (_08306_, _08304_, _07399_);
  nor _59743_ (_08307_, _08289_, _05182_);
  nor _59744_ (_08308_, _08307_, _08302_);
  nor _59745_ (_08309_, _08308_, _07405_);
  nor _59746_ (_08310_, _08309_, _08306_);
  nor _59747_ (_08311_, _08310_, _08305_);
  nor _59748_ (_08312_, _08306_, _08305_);
  not _59749_ (_08313_, _08312_);
  and _59750_ (_08314_, _08308_, _07405_);
  or _59751_ (_08315_, _08314_, _08309_);
  or _59752_ (_08316_, _08315_, _08313_);
  nor _59753_ (_08317_, _06032_, _03563_);
  nor _59754_ (_08318_, _08317_, _08289_);
  nor _59755_ (_08319_, _08318_, _07500_);
  and _59756_ (_08320_, _08318_, _07500_);
  nor _59757_ (_08321_, _08320_, _08319_);
  nor _59758_ (_08322_, _08288_, _04965_);
  nor _59759_ (_08323_, _08322_, _06032_);
  nor _59760_ (_08324_, _08323_, _07506_);
  and _59761_ (_08325_, _08323_, _07506_);
  nor _59762_ (_08326_, _08325_, _08324_);
  and _59763_ (_08327_, _08326_, _08321_);
  nor _59764_ (_08328_, _03471_, _07888_);
  nor _59765_ (_08329_, _08328_, _04548_);
  nor _59766_ (_08330_, _08329_, _08288_);
  nor _59767_ (_08331_, _08330_, _03233_);
  and _59768_ (_08332_, _08330_, _03233_);
  and _59769_ (_08333_, _03471_, _07888_);
  nor _59770_ (_08334_, _08333_, _08328_);
  and _59771_ (_08335_, _08334_, _03321_);
  nor _59772_ (_08336_, _08335_, _08332_);
  or _59773_ (_08337_, _08336_, _08331_);
  nand _59774_ (_08338_, _08337_, _08327_);
  and _59775_ (_08339_, _08324_, _08321_);
  nor _59776_ (_08340_, _08339_, _08319_);
  and _59777_ (_08341_, _08340_, _08338_);
  nor _59778_ (_08342_, _08341_, _08316_);
  nor _59779_ (_08343_, _08342_, _08311_);
  and _59780_ (_08344_, _08300_, _07346_);
  nor _59781_ (_08345_, _08301_, _08344_);
  not _59782_ (_08346_, _08345_);
  nor _59783_ (_08347_, _08346_, _08343_);
  or _59784_ (_08348_, _08347_, _08301_);
  and _59785_ (_08349_, _08348_, _08298_);
  nor _59786_ (_08350_, _08348_, _08298_);
  or _59787_ (_08351_, _08350_, _08349_);
  and _59788_ (_08352_, _08351_, _08108_);
  or _59789_ (_08353_, _08352_, _03311_);
  or _59790_ (_08354_, _08353_, _08287_);
  or _59791_ (_08355_, _03401_, _03254_);
  and _59792_ (_08356_, _08355_, _03500_);
  and _59793_ (_08357_, _08356_, _08354_);
  not _59794_ (_08358_, _05792_);
  nor _59795_ (_08359_, _06034_, _08358_);
  nor _59796_ (_08360_, _08359_, _07977_);
  nor _59797_ (_08361_, _08360_, _03500_);
  or _59798_ (_08362_, _08361_, _07314_);
  or _59799_ (_08363_, _08362_, _08357_);
  and _59800_ (_08364_, _08363_, _07921_);
  or _59801_ (_08365_, _08364_, _03479_);
  and _59802_ (_08366_, _05935_, _05227_);
  nor _59803_ (_08367_, _08366_, _07915_);
  nand _59804_ (_08368_, _08367_, _03479_);
  and _59805_ (_08369_, _08368_, _03474_);
  and _59806_ (_08370_, _08369_, _08365_);
  nor _59807_ (_08371_, _06292_, _07918_);
  nor _59808_ (_08372_, _08371_, _07915_);
  nor _59809_ (_08373_, _08372_, _03474_);
  or _59810_ (_08374_, _08373_, _07328_);
  or _59811_ (_08375_, _08374_, _08370_);
  and _59812_ (_08376_, \oc8051_golden_model_1.B [0], _05834_);
  not _59813_ (_08377_, _08376_);
  and _59814_ (_08378_, _08377_, _07344_);
  not _59815_ (_08379_, _08378_);
  nand _59816_ (_08380_, _08379_, _07328_);
  and _59817_ (_08381_, _08380_, _08375_);
  or _59818_ (_08382_, _08381_, _03231_);
  and _59819_ (_08383_, _08382_, _07917_);
  or _59820_ (_08384_, _08383_, _03437_);
  and _59821_ (_08385_, _03637_, _03188_);
  not _59822_ (_08386_, _08385_);
  and _59823_ (_08387_, _06087_, _05227_);
  nor _59824_ (_08388_, _08387_, _07915_);
  nand _59825_ (_08389_, _08388_, _03437_);
  and _59826_ (_08390_, _08389_, _08386_);
  and _59827_ (_08391_, _08390_, _08384_);
  not _59828_ (_08392_, _03936_);
  and _59829_ (_08393_, _08385_, _03401_);
  or _59830_ (_08394_, _08393_, _08392_);
  or _59831_ (_08395_, _08394_, _08391_);
  nor _59832_ (_08396_, _04325_, _04123_);
  and _59833_ (_08397_, _08396_, _03936_);
  and _59834_ (_08398_, _08396_, _07784_);
  or _59835_ (_08399_, _08398_, _08397_);
  and _59836_ (_08400_, _08399_, _08395_);
  not _59837_ (_08401_, _08396_);
  and _59838_ (_08402_, _08401_, _07784_);
  or _59839_ (_08403_, _08402_, _04128_);
  or _59840_ (_08404_, _08403_, _08400_);
  and _59841_ (_08405_, _03478_, _03193_);
  not _59842_ (_08406_, _08405_);
  and _59843_ (_08407_, _08406_, _07784_);
  or _59844_ (_08408_, _08405_, _04128_);
  not _59845_ (_08409_, _08408_);
  or _59846_ (_08410_, _08409_, _08407_);
  and _59847_ (_08411_, _08410_, _08404_);
  and _59848_ (_08412_, _08405_, _07735_);
  or _59849_ (_08413_, _08412_, _03767_);
  or _59850_ (_08414_, _08413_, _08411_);
  and _59851_ (_08415_, _03637_, _03193_);
  not _59852_ (_08416_, _08415_);
  or _59853_ (_08417_, _06311_, _03768_);
  and _59854_ (_08418_, _08417_, _08416_);
  and _59855_ (_08419_, _08418_, _08414_);
  nor _59856_ (_08420_, _03401_, \oc8051_golden_model_1.ACC [7]);
  and _59857_ (_08421_, _03401_, \oc8051_golden_model_1.ACC [7]);
  nor _59858_ (_08422_, _08421_, _08420_);
  and _59859_ (_08423_, _08415_, _08422_);
  or _59860_ (_08424_, _08423_, _03636_);
  or _59861_ (_08425_, _08424_, _08419_);
  and _59862_ (_08426_, _06305_, _05227_);
  nor _59863_ (_08427_, _08426_, _07915_);
  nand _59864_ (_08428_, _08427_, _03636_);
  and _59865_ (_08429_, _08428_, _04501_);
  and _59866_ (_08430_, _08429_, _08425_);
  or _59867_ (_08431_, _08430_, _07916_);
  nand _59868_ (_08432_, _03481_, _03191_);
  and _59869_ (_08433_, _08432_, _08431_);
  not _59870_ (_08434_, _04345_);
  and _59871_ (_08435_, _08432_, _08434_);
  not _59872_ (_08436_, _08435_);
  or _59873_ (_08437_, _07782_, _04345_);
  and _59874_ (_08438_, _08437_, _08436_);
  or _59875_ (_08439_, _08438_, _08433_);
  not _59876_ (_08440_, _04135_);
  or _59877_ (_08441_, _07782_, _08434_);
  and _59878_ (_08442_, _08441_, _08440_);
  and _59879_ (_08443_, _08442_, _08439_);
  or _59880_ (_08444_, _08443_, _07914_);
  and _59881_ (_08445_, _03478_, _03191_);
  not _59882_ (_08446_, _08445_);
  and _59883_ (_08447_, _08446_, _08444_);
  and _59884_ (_08448_, _08445_, _07734_);
  or _59885_ (_08449_, _08448_, _03755_);
  or _59886_ (_08450_, _08449_, _08447_);
  and _59887_ (_08451_, _08450_, _07913_);
  and _59888_ (_08452_, _08421_, _07909_);
  or _59889_ (_08453_, _08452_, _08451_);
  and _59890_ (_08454_, _08453_, _05769_);
  and _59891_ (_08455_, _03661_, _03182_);
  and _59892_ (_08456_, _03481_, _03182_);
  nor _59893_ (_08457_, _08456_, _08455_);
  not _59894_ (_08458_, _08457_);
  or _59895_ (_08459_, _08388_, _06310_);
  nor _59896_ (_08460_, _08459_, _04505_);
  or _59897_ (_08461_, _08460_, _08458_);
  or _59898_ (_08462_, _08461_, _08454_);
  nand _59899_ (_08463_, _08458_, _07783_);
  not _59900_ (_08464_, _03182_);
  nor _59901_ (_08465_, _03665_, _08464_);
  nor _59902_ (_08466_, _08465_, _04161_);
  and _59903_ (_08467_, _08466_, _08463_);
  and _59904_ (_08468_, _08467_, _08462_);
  and _59905_ (_08469_, _03478_, _03182_);
  nor _59906_ (_08470_, _08466_, _07783_);
  or _59907_ (_08471_, _08470_, _08469_);
  or _59908_ (_08472_, _08471_, _08468_);
  not _59909_ (_08473_, _03761_);
  nand _59910_ (_08474_, _08469_, _07733_);
  and _59911_ (_08475_, _08474_, _08473_);
  and _59912_ (_08476_, _08475_, _08472_);
  and _59913_ (_08477_, _03637_, _03182_);
  nor _59914_ (_08478_, _08477_, _03761_);
  not _59915_ (_08479_, _08478_);
  not _59916_ (_08480_, _08477_);
  nand _59917_ (_08481_, _08480_, _06310_);
  and _59918_ (_08482_, _08481_, _08479_);
  or _59919_ (_08483_, _08482_, _08476_);
  nand _59920_ (_08484_, _08477_, _08420_);
  and _59921_ (_08485_, _08484_, _03759_);
  and _59922_ (_08486_, _08485_, _08483_);
  nor _59923_ (_08487_, _06304_, _07918_);
  nor _59924_ (_08488_, _08487_, _07915_);
  nor _59925_ (_08489_, _08488_, _03759_);
  not _59926_ (_08490_, _07830_);
  or _59927_ (_08491_, _08490_, _08489_);
  or _59928_ (_08492_, _08491_, _08486_);
  and _59929_ (_08493_, _08492_, _07908_);
  or _59930_ (_08494_, _08493_, _07825_);
  not _59931_ (_08495_, _07825_);
  and _59932_ (_08496_, _08050_, \oc8051_golden_model_1.ACC [6]);
  and _59933_ (_08497_, _08053_, \oc8051_golden_model_1.ACC [5]);
  and _59934_ (_08498_, _08059_, \oc8051_golden_model_1.ACC [4]);
  and _59935_ (_08499_, _08071_, \oc8051_golden_model_1.ACC [3]);
  and _59936_ (_08500_, _08076_, \oc8051_golden_model_1.ACC [2]);
  and _59937_ (_08501_, _08083_, \oc8051_golden_model_1.ACC [1]);
  nor _59938_ (_08502_, _08085_, _08084_);
  and _59939_ (_08503_, _08087_, \oc8051_golden_model_1.ACC [0]);
  not _59940_ (_08504_, _08503_);
  nor _59941_ (_08505_, _08504_, _08502_);
  nor _59942_ (_08506_, _08505_, _08501_);
  nor _59943_ (_08507_, _08506_, _08079_);
  nor _59944_ (_08508_, _08507_, _08500_);
  nor _59945_ (_08509_, _08508_, _08074_);
  or _59946_ (_08510_, _08509_, _08499_);
  and _59947_ (_08511_, _08510_, _08066_);
  nor _59948_ (_08512_, _08511_, _08498_);
  nor _59949_ (_08513_, _08512_, _08063_);
  or _59950_ (_08514_, _08513_, _08497_);
  and _59951_ (_08515_, _08514_, _08099_);
  nor _59952_ (_08516_, _08515_, _08496_);
  nor _59953_ (_08517_, _08516_, _08044_);
  and _59954_ (_08518_, _08516_, _08044_);
  nor _59955_ (_08519_, _08518_, _08517_);
  or _59956_ (_08520_, _08519_, _08495_);
  and _59957_ (_08521_, _08520_, _03766_);
  and _59958_ (_08522_, _08521_, _08494_);
  and _59959_ (_08523_, _03637_, _03177_);
  nor _59960_ (_08524_, _08523_, _03765_);
  not _59961_ (_08525_, _08524_);
  and _59962_ (_08526_, _08233_, \oc8051_golden_model_1.ACC [6]);
  not _59963_ (_08527_, _08279_);
  and _59964_ (_08528_, _08239_, \oc8051_golden_model_1.ACC [5]);
  and _59965_ (_08529_, _08243_, \oc8051_golden_model_1.ACC [4]);
  not _59966_ (_08530_, _08249_);
  and _59967_ (_08531_, _08253_, \oc8051_golden_model_1.ACC [3]);
  and _59968_ (_08532_, _08258_, \oc8051_golden_model_1.ACC [2]);
  and _59969_ (_08533_, _08264_, \oc8051_golden_model_1.ACC [1]);
  nor _59970_ (_08534_, _08265_, _08266_);
  and _59971_ (_08535_, _08268_, \oc8051_golden_model_1.ACC [0]);
  not _59972_ (_08536_, _08535_);
  nor _59973_ (_08537_, _08536_, _08534_);
  nor _59974_ (_08538_, _08537_, _08533_);
  nor _59975_ (_08539_, _08538_, _08261_);
  nor _59976_ (_08540_, _08539_, _08532_);
  nor _59977_ (_08541_, _08540_, _08256_);
  or _59978_ (_08542_, _08541_, _08531_);
  and _59979_ (_08543_, _08542_, _08530_);
  nor _59980_ (_08544_, _08543_, _08529_);
  nor _59981_ (_08545_, _08544_, _08247_);
  or _59982_ (_08546_, _08545_, _08528_);
  and _59983_ (_08547_, _08546_, _08527_);
  nor _59984_ (_08548_, _08547_, _08526_);
  nor _59985_ (_08549_, _08548_, _08231_);
  and _59986_ (_08550_, _08548_, _08231_);
  nor _59987_ (_08551_, _08550_, _08549_);
  or _59988_ (_08552_, _08551_, _08523_);
  and _59989_ (_08553_, _08552_, _08525_);
  or _59990_ (_08554_, _08553_, _08522_);
  and _59991_ (_08555_, _03230_, _03177_);
  not _59992_ (_08556_, _08555_);
  not _59993_ (_08557_, _08523_);
  and _59994_ (_08558_, _08300_, \oc8051_golden_model_1.ACC [6]);
  and _59995_ (_08559_, _08304_, \oc8051_golden_model_1.ACC [5]);
  and _59996_ (_08560_, _08308_, \oc8051_golden_model_1.ACC [4]);
  and _59997_ (_08561_, _08318_, \oc8051_golden_model_1.ACC [3]);
  and _59998_ (_08562_, _08323_, \oc8051_golden_model_1.ACC [2]);
  and _59999_ (_08563_, _08330_, \oc8051_golden_model_1.ACC [1]);
  nor _60000_ (_08564_, _08332_, _08331_);
  and _60001_ (_08565_, _08334_, \oc8051_golden_model_1.ACC [0]);
  not _60002_ (_08566_, _08565_);
  nor _60003_ (_08567_, _08566_, _08564_);
  nor _60004_ (_08568_, _08567_, _08563_);
  nor _60005_ (_08569_, _08568_, _08326_);
  nor _60006_ (_08570_, _08569_, _08562_);
  nor _60007_ (_08571_, _08570_, _08321_);
  or _60008_ (_08572_, _08571_, _08561_);
  and _60009_ (_08573_, _08572_, _08315_);
  nor _60010_ (_08574_, _08573_, _08560_);
  nor _60011_ (_08575_, _08574_, _08312_);
  or _60012_ (_08576_, _08575_, _08559_);
  and _60013_ (_08577_, _08576_, _08346_);
  nor _60014_ (_08578_, _08577_, _08558_);
  nor _60015_ (_08579_, _08578_, _08297_);
  and _60016_ (_08580_, _08578_, _08297_);
  nor _60017_ (_08581_, _08580_, _08579_);
  or _60018_ (_08582_, _08581_, _08557_);
  and _60019_ (_08583_, _08582_, _08556_);
  and _60020_ (_08584_, _08583_, _08554_);
  nor _60021_ (_08585_, _07777_, _04178_);
  and _60022_ (_08586_, _08555_, \oc8051_golden_model_1.ACC [6]);
  nor _60023_ (_08587_, _03665_, _04178_);
  or _60024_ (_08588_, _08587_, _08586_);
  or _60025_ (_08589_, _08588_, _08585_);
  or _60026_ (_08590_, _08589_, _08584_);
  and _60027_ (_08591_, _08590_, _07824_);
  and _60028_ (_08592_, _07821_, _07781_);
  or _60029_ (_08593_, _08592_, _07731_);
  or _60030_ (_08594_, _08593_, _08591_);
  and _60031_ (_08595_, _08594_, _07773_);
  or _60032_ (_08596_, _08595_, _03524_);
  and _60033_ (_08597_, _03637_, _03171_);
  not _60034_ (_08598_, _08597_);
  and _60035_ (_08599_, _05984_, _05834_);
  nor _60036_ (_08600_, _05984_, _05834_);
  nor _60037_ (_08601_, _08600_, _08599_);
  nor _60038_ (_08602_, _08125_, _07346_);
  and _60039_ (_08603_, _08125_, \oc8051_golden_model_1.ACC [6]);
  nor _60040_ (_08604_, _08125_, \oc8051_golden_model_1.ACC [6]);
  nor _60041_ (_08605_, _08604_, _08603_);
  not _60042_ (_08606_, _08605_);
  nor _60043_ (_08607_, _08205_, _07399_);
  nor _60044_ (_08608_, _08205_, \oc8051_golden_model_1.ACC [5]);
  and _60045_ (_08609_, _08205_, \oc8051_golden_model_1.ACC [5]);
  nor _60046_ (_08610_, _08609_, _08608_);
  nor _60047_ (_08611_, _08222_, _07405_);
  and _60048_ (_08612_, _08222_, \oc8051_golden_model_1.ACC [4]);
  nor _60049_ (_08613_, _08222_, \oc8051_golden_model_1.ACC [4]);
  nor _60050_ (_08614_, _08613_, _08612_);
  not _60051_ (_08615_, _08614_);
  nand _60052_ (_08616_, _08143_, _07500_);
  or _60053_ (_08617_, _08143_, _07500_);
  nor _60054_ (_08618_, _08163_, _07506_);
  and _60055_ (_08619_, _08163_, \oc8051_golden_model_1.ACC [2]);
  nor _60056_ (_08620_, _08163_, \oc8051_golden_model_1.ACC [2]);
  nor _60057_ (_08621_, _08620_, _08619_);
  nor _60058_ (_08622_, _08177_, _03233_);
  nor _60059_ (_08623_, _08177_, \oc8051_golden_model_1.ACC [1]);
  and _60060_ (_08624_, _08177_, \oc8051_golden_model_1.ACC [1]);
  nor _60061_ (_08625_, _08624_, _08623_);
  nor _60062_ (_08626_, _08191_, _03321_);
  not _60063_ (_08627_, _08626_);
  nor _60064_ (_08628_, _08627_, _08625_);
  nor _60065_ (_08629_, _08628_, _08622_);
  nor _60066_ (_08630_, _08629_, _08621_);
  nor _60067_ (_08631_, _08630_, _08618_);
  nand _60068_ (_08632_, _08631_, _08617_);
  and _60069_ (_08633_, _08632_, _08616_);
  and _60070_ (_08634_, _08633_, _08615_);
  nor _60071_ (_08635_, _08634_, _08611_);
  nor _60072_ (_08636_, _08635_, _08610_);
  or _60073_ (_08637_, _08636_, _08607_);
  and _60074_ (_08638_, _08637_, _08606_);
  nor _60075_ (_08639_, _08638_, _08602_);
  nor _60076_ (_08640_, _08639_, _08601_);
  and _60077_ (_08641_, _08639_, _08601_);
  or _60078_ (_08642_, _08641_, _08640_);
  or _60079_ (_08643_, _08642_, _03526_);
  and _60080_ (_08644_, _08643_, _08598_);
  and _60081_ (_08645_, _08644_, _08596_);
  nor _60082_ (_08646_, _03561_, _07346_);
  and _60083_ (_08647_, _03561_, _07346_);
  or _60084_ (_08648_, _08647_, _08646_);
  not _60085_ (_08649_, _08648_);
  nor _60086_ (_08650_, _03834_, _07399_);
  and _60087_ (_08651_, _03834_, _07399_);
  nor _60088_ (_08652_, _08650_, _08651_);
  not _60089_ (_08653_, _08652_);
  nor _60090_ (_08654_, _04249_, _07405_);
  and _60091_ (_08655_, _04249_, _07405_);
  nor _60092_ (_08656_, _08654_, _08655_);
  nor _60093_ (_08657_, _03432_, _07500_);
  and _60094_ (_08658_, _03432_, _07500_);
  nor _60095_ (_08659_, _03877_, _07506_);
  and _60096_ (_08660_, _03877_, _07506_);
  nor _60097_ (_08661_, _08659_, _08660_);
  not _60098_ (_08662_, _08661_);
  nor _60099_ (_08663_, _04284_, _03233_);
  and _60100_ (_08664_, _04284_, _03233_);
  nor _60101_ (_08665_, _08663_, _08664_);
  nor _60102_ (_08666_, _03471_, _03321_);
  and _60103_ (_08667_, _08666_, _08665_);
  nor _60104_ (_08668_, _08667_, _08663_);
  nor _60105_ (_08669_, _08668_, _08662_);
  nor _60106_ (_08670_, _08669_, _08659_);
  nor _60107_ (_08671_, _08670_, _08658_);
  or _60108_ (_08672_, _08671_, _08657_);
  and _60109_ (_08673_, _08672_, _08656_);
  nor _60110_ (_08674_, _08673_, _08654_);
  nor _60111_ (_08675_, _08674_, _08653_);
  or _60112_ (_08676_, _08675_, _08650_);
  and _60113_ (_08677_, _08676_, _08649_);
  nor _60114_ (_08678_, _08677_, _08646_);
  nor _60115_ (_08679_, _08678_, _08422_);
  and _60116_ (_08680_, _08678_, _08422_);
  nor _60117_ (_08681_, _08680_, _08679_);
  nor _60118_ (_08682_, _08681_, _08598_);
  or _60119_ (_08683_, _08682_, _07729_);
  or _60120_ (_08684_, _08683_, _08645_);
  and _60121_ (_08685_, _08684_, _07730_);
  or _60122_ (_08686_, _08685_, _03790_);
  and _60123_ (_08687_, _03637_, _03010_);
  not _60124_ (_08688_, _08687_);
  nand _60125_ (_08689_, _07950_, _03790_);
  and _60126_ (_08690_, _08689_, _08688_);
  and _60127_ (_08691_, _08690_, _08686_);
  and _60128_ (_08692_, _03230_, _03010_);
  nor _60129_ (_08693_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and _60130_ (_08694_, _08693_, _07443_);
  and _60131_ (_08695_, _08694_, _07363_);
  and _60132_ (_08696_, _08695_, _07346_);
  nor _60133_ (_08697_, _08696_, _05834_);
  and _60134_ (_08698_, _08696_, _05834_);
  nor _60135_ (_08699_, _08698_, _08697_);
  nor _60136_ (_08700_, _08699_, _08688_);
  or _60137_ (_08701_, _08700_, _08692_);
  or _60138_ (_08702_, _08701_, _08691_);
  nand _60139_ (_08703_, _08692_, _07888_);
  and _60140_ (_08704_, _08703_, _03152_);
  and _60141_ (_08705_, _08704_, _08702_);
  nor _60142_ (_08706_, _07999_, _03152_);
  or _60143_ (_08707_, _08706_, _03520_);
  or _60144_ (_08708_, _08707_, _08705_);
  and _60145_ (_08709_, _03637_, _03165_);
  not _60146_ (_08710_, _08709_);
  and _60147_ (_08711_, _05767_, _05227_);
  nor _60148_ (_08712_, _08711_, _07915_);
  nand _60149_ (_08713_, _08712_, _03520_);
  and _60150_ (_08714_, _08713_, _08710_);
  and _60151_ (_08715_, _08714_, _08708_);
  and _60152_ (_08716_, _03230_, _03165_);
  and _60153_ (_08717_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand _60154_ (_08718_, _08717_, _07444_);
  nor _60155_ (_08719_, _08718_, _07405_);
  and _60156_ (_08720_, _08719_, \oc8051_golden_model_1.ACC [5]);
  and _60157_ (_08721_, _08720_, \oc8051_golden_model_1.ACC [6]);
  nor _60158_ (_08722_, _08721_, \oc8051_golden_model_1.ACC [7]);
  and _60159_ (_08723_, _08721_, \oc8051_golden_model_1.ACC [7]);
  nor _60160_ (_08724_, _08723_, _08722_);
  and _60161_ (_08725_, _08724_, _08709_);
  or _60162_ (_08726_, _08725_, _08716_);
  or _60163_ (_08727_, _08726_, _08715_);
  nand _60164_ (_08728_, _08716_, _03321_);
  and _60165_ (_08729_, _08728_, _42963_);
  and _60166_ (_08730_, _08729_, _08727_);
  or _60167_ (_08731_, _08730_, _07728_);
  and _60168_ (_40516_, _08731_, _41755_);
  not _60169_ (_08732_, \oc8051_golden_model_1.SBUF [7]);
  nor _60170_ (_08733_, _05185_, _08732_);
  and _60171_ (_08734_, _06311_, _05185_);
  nor _60172_ (_08735_, _08734_, _08733_);
  nor _60173_ (_08736_, _08735_, _04501_);
  not _60174_ (_08737_, _05185_);
  nor _60175_ (_08738_, _08737_, _05176_);
  nor _60176_ (_08739_, _08738_, _08733_);
  and _60177_ (_08740_, _08739_, _07314_);
  and _60178_ (_08741_, _05185_, \oc8051_golden_model_1.ACC [7]);
  nor _60179_ (_08742_, _08741_, _08733_);
  nor _60180_ (_08743_, _08742_, _03583_);
  nor _60181_ (_08744_, _08742_, _04427_);
  nor _60182_ (_08745_, _04426_, _08732_);
  or _60183_ (_08746_, _08745_, _08744_);
  and _60184_ (_08747_, _08746_, _04444_);
  and _60185_ (_08748_, _05949_, _05185_);
  nor _60186_ (_08749_, _08748_, _08733_);
  nor _60187_ (_08750_, _08749_, _04444_);
  or _60188_ (_08751_, _08750_, _08747_);
  and _60189_ (_08752_, _08751_, _03983_);
  nor _60190_ (_08753_, _08739_, _03983_);
  nor _60191_ (_08754_, _08753_, _08752_);
  nor _60192_ (_08755_, _08754_, _03575_);
  or _60193_ (_08756_, _08755_, _07314_);
  nor _60194_ (_08757_, _08756_, _08743_);
  nor _60195_ (_08758_, _08757_, _08740_);
  nor _60196_ (_08759_, _08758_, _03479_);
  and _60197_ (_08760_, _05935_, _05185_);
  nor _60198_ (_08761_, _08733_, _06044_);
  not _60199_ (_08762_, _08761_);
  nor _60200_ (_08763_, _08762_, _08760_);
  or _60201_ (_08764_, _08763_, _03221_);
  nor _60202_ (_08765_, _08764_, _08759_);
  nor _60203_ (_08766_, _06292_, _08737_);
  nor _60204_ (_08767_, _08766_, _08733_);
  nor _60205_ (_08768_, _08767_, _03474_);
  or _60206_ (_08769_, _08768_, _03437_);
  or _60207_ (_08770_, _08769_, _08765_);
  and _60208_ (_08771_, _06087_, _05185_);
  nor _60209_ (_08772_, _08771_, _08733_);
  nand _60210_ (_08773_, _08772_, _03437_);
  and _60211_ (_08774_, _08773_, _08770_);
  nor _60212_ (_08775_, _08774_, _03636_);
  and _60213_ (_08776_, _06305_, _05185_);
  or _60214_ (_08777_, _08733_, _04499_);
  nor _60215_ (_08778_, _08777_, _08776_);
  or _60216_ (_08779_, _08778_, _03769_);
  nor _60217_ (_08780_, _08779_, _08775_);
  nor _60218_ (_08781_, _08780_, _08736_);
  nor _60219_ (_08782_, _08781_, _04504_);
  not _60220_ (_08783_, _08733_);
  and _60221_ (_08784_, _08783_, _05281_);
  or _60222_ (_08785_, _08772_, _04505_);
  nor _60223_ (_08786_, _08785_, _08784_);
  nor _60224_ (_08787_, _08786_, _08782_);
  nor _60225_ (_08788_, _08787_, _03752_);
  or _60226_ (_08789_, _08784_, _03753_);
  nor _60227_ (_08790_, _08789_, _08742_);
  or _60228_ (_08791_, _08790_, _08788_);
  and _60229_ (_08792_, _08791_, _03759_);
  nor _60230_ (_08793_, _06304_, _08737_);
  nor _60231_ (_08794_, _08793_, _08733_);
  nor _60232_ (_08795_, _08794_, _03759_);
  or _60233_ (_08796_, _08795_, _08792_);
  and _60234_ (_08797_, _08796_, _04517_);
  nor _60235_ (_08798_, _06310_, _08737_);
  nor _60236_ (_08799_, _08798_, _08733_);
  nor _60237_ (_08800_, _08799_, _04517_);
  or _60238_ (_08801_, _08800_, _03790_);
  nor _60239_ (_08802_, _08801_, _08797_);
  and _60240_ (_08803_, _08749_, _03790_);
  or _60241_ (_08804_, _08803_, _03520_);
  nor _60242_ (_08805_, _08804_, _08802_);
  and _60243_ (_08806_, _05767_, _05185_);
  nor _60244_ (_08807_, _08806_, _08733_);
  nor _60245_ (_08808_, _08807_, _03521_);
  or _60246_ (_08809_, _08808_, _08805_);
  or _60247_ (_08810_, _08809_, _42967_);
  or _60248_ (_08811_, _42963_, \oc8051_golden_model_1.SBUF [7]);
  and _60249_ (_08812_, _08811_, _41755_);
  and _60250_ (_40517_, _08812_, _08810_);
  not _60251_ (_08813_, \oc8051_golden_model_1.SCON [7]);
  nor _60252_ (_08814_, _05248_, _08813_);
  and _60253_ (_08815_, _06311_, _05248_);
  nor _60254_ (_08816_, _08815_, _08814_);
  nor _60255_ (_08817_, _08816_, _04501_);
  not _60256_ (_08818_, _05248_);
  nor _60257_ (_08819_, _08818_, _05176_);
  nor _60258_ (_08820_, _08819_, _08814_);
  and _60259_ (_08821_, _08820_, _07314_);
  nor _60260_ (_08822_, _05805_, _08813_);
  and _60261_ (_08823_, _05818_, _05805_);
  nor _60262_ (_08824_, _08823_, _08822_);
  nor _60263_ (_08825_, _08824_, _03513_);
  and _60264_ (_08826_, _05248_, \oc8051_golden_model_1.ACC [7]);
  nor _60265_ (_08827_, _08826_, _08814_);
  nor _60266_ (_08828_, _08827_, _04427_);
  nor _60267_ (_08829_, _04426_, _08813_);
  or _60268_ (_08830_, _08829_, _08828_);
  and _60269_ (_08831_, _08830_, _04444_);
  and _60270_ (_08832_, _05949_, _05248_);
  nor _60271_ (_08833_, _08832_, _08814_);
  nor _60272_ (_08834_, _08833_, _04444_);
  or _60273_ (_08835_, _08834_, _08831_);
  and _60274_ (_08836_, _08835_, _03517_);
  and _60275_ (_08837_, _05954_, _05805_);
  nor _60276_ (_08838_, _08837_, _08822_);
  nor _60277_ (_08839_, _08838_, _03517_);
  or _60278_ (_08840_, _08839_, _03568_);
  or _60279_ (_08841_, _08840_, _08836_);
  nand _60280_ (_08842_, _08820_, _03568_);
  and _60281_ (_08843_, _08842_, _08841_);
  and _60282_ (_08844_, _08843_, _03583_);
  nor _60283_ (_08845_, _08827_, _03583_);
  or _60284_ (_08846_, _08845_, _08844_);
  and _60285_ (_08847_, _08846_, _03513_);
  nor _60286_ (_08848_, _08847_, _08825_);
  nor _60287_ (_08849_, _08848_, _03505_);
  nor _60288_ (_08850_, _08822_, _05989_);
  or _60289_ (_08851_, _08838_, _03506_);
  nor _60290_ (_08852_, _08851_, _08850_);
  nor _60291_ (_08853_, _08852_, _08849_);
  nor _60292_ (_08854_, _08853_, _03499_);
  not _60293_ (_08855_, _05805_);
  nor _60294_ (_08856_, _06034_, _08855_);
  nor _60295_ (_08857_, _08856_, _08822_);
  nor _60296_ (_08858_, _08857_, _03500_);
  nor _60297_ (_08859_, _08858_, _07314_);
  not _60298_ (_08860_, _08859_);
  nor _60299_ (_08861_, _08860_, _08854_);
  nor _60300_ (_08862_, _08861_, _08821_);
  nor _60301_ (_08863_, _08862_, _03479_);
  and _60302_ (_08864_, _05935_, _05248_);
  nor _60303_ (_08865_, _08814_, _06044_);
  not _60304_ (_08866_, _08865_);
  nor _60305_ (_08867_, _08866_, _08864_);
  nor _60306_ (_08868_, _08867_, _03221_);
  not _60307_ (_08869_, _08868_);
  nor _60308_ (_08870_, _08869_, _08863_);
  nor _60309_ (_08871_, _06292_, _08818_);
  nor _60310_ (_08872_, _08871_, _08814_);
  nor _60311_ (_08873_, _08872_, _03474_);
  or _60312_ (_08874_, _08873_, _03437_);
  or _60313_ (_08875_, _08874_, _08870_);
  and _60314_ (_08876_, _06087_, _05248_);
  nor _60315_ (_08877_, _08876_, _08814_);
  nand _60316_ (_08878_, _08877_, _03437_);
  and _60317_ (_08879_, _08878_, _08875_);
  nor _60318_ (_08880_, _08879_, _03636_);
  and _60319_ (_08881_, _06305_, _05248_);
  or _60320_ (_08882_, _08814_, _04499_);
  nor _60321_ (_08883_, _08882_, _08881_);
  or _60322_ (_08884_, _08883_, _03769_);
  nor _60323_ (_08885_, _08884_, _08880_);
  nor _60324_ (_08886_, _08885_, _08817_);
  nor _60325_ (_08887_, _08886_, _04504_);
  not _60326_ (_08888_, _08814_);
  and _60327_ (_08889_, _08888_, _05281_);
  or _60328_ (_08890_, _08877_, _04505_);
  nor _60329_ (_08891_, _08890_, _08889_);
  nor _60330_ (_08892_, _08891_, _08887_);
  nor _60331_ (_08893_, _08892_, _03752_);
  or _60332_ (_08894_, _08889_, _03753_);
  or _60333_ (_08895_, _08894_, _08827_);
  and _60334_ (_08896_, _08895_, _03759_);
  not _60335_ (_08897_, _08896_);
  nor _60336_ (_08898_, _08897_, _08893_);
  nor _60337_ (_08899_, _06304_, _08818_);
  or _60338_ (_08900_, _08814_, _03759_);
  nor _60339_ (_08901_, _08900_, _08899_);
  or _60340_ (_08902_, _08901_, _03760_);
  nor _60341_ (_08903_, _08902_, _08898_);
  nor _60342_ (_08904_, _06310_, _08818_);
  nor _60343_ (_08905_, _08904_, _08814_);
  nor _60344_ (_08906_, _08905_, _04517_);
  or _60345_ (_08907_, _08906_, _08903_);
  and _60346_ (_08908_, _08907_, _04192_);
  nor _60347_ (_08909_, _08833_, _04192_);
  or _60348_ (_08910_, _08909_, _08908_);
  and _60349_ (_08911_, _08910_, _03152_);
  nor _60350_ (_08912_, _08824_, _03152_);
  or _60351_ (_08913_, _08912_, _08911_);
  and _60352_ (_08914_, _08913_, _03521_);
  and _60353_ (_08915_, _05767_, _05248_);
  nor _60354_ (_08916_, _08915_, _08814_);
  nor _60355_ (_08917_, _08916_, _03521_);
  or _60356_ (_08918_, _08917_, _08914_);
  or _60357_ (_08919_, _08918_, _42967_);
  or _60358_ (_08920_, _42963_, \oc8051_golden_model_1.SCON [7]);
  and _60359_ (_08921_, _08920_, _41755_);
  and _60360_ (_40518_, _08921_, _08919_);
  not _60361_ (_08922_, \oc8051_golden_model_1.PCON [7]);
  nor _60362_ (_08923_, _05208_, _08922_);
  and _60363_ (_08924_, _06311_, _05208_);
  nor _60364_ (_08925_, _08924_, _08923_);
  nor _60365_ (_08926_, _08925_, _04501_);
  and _60366_ (_08927_, _05208_, \oc8051_golden_model_1.ACC [7]);
  nor _60367_ (_08928_, _08927_, _08923_);
  nor _60368_ (_08929_, _08928_, _03583_);
  nor _60369_ (_08930_, _08928_, _04427_);
  nor _60370_ (_08931_, _04426_, _08922_);
  or _60371_ (_08933_, _08931_, _08930_);
  and _60372_ (_08934_, _08933_, _04444_);
  and _60373_ (_08935_, _05949_, _05208_);
  nor _60374_ (_08936_, _08935_, _08923_);
  nor _60375_ (_08937_, _08936_, _04444_);
  or _60376_ (_08938_, _08937_, _08934_);
  and _60377_ (_08939_, _08938_, _03983_);
  not _60378_ (_08940_, _05208_);
  nor _60379_ (_08941_, _08940_, _05176_);
  nor _60380_ (_08942_, _08941_, _08923_);
  nor _60381_ (_08944_, _08942_, _03983_);
  nor _60382_ (_08945_, _08944_, _08939_);
  nor _60383_ (_08946_, _08945_, _03575_);
  or _60384_ (_08947_, _08946_, _07314_);
  nor _60385_ (_08948_, _08947_, _08929_);
  and _60386_ (_08949_, _08942_, _07314_);
  nor _60387_ (_08950_, _08949_, _08948_);
  nor _60388_ (_08951_, _08950_, _03479_);
  and _60389_ (_08952_, _05935_, _05208_);
  nor _60390_ (_08953_, _08923_, _06044_);
  not _60391_ (_08955_, _08953_);
  nor _60392_ (_08956_, _08955_, _08952_);
  or _60393_ (_08957_, _08956_, _03221_);
  nor _60394_ (_08958_, _08957_, _08951_);
  nor _60395_ (_08959_, _06292_, _08940_);
  nor _60396_ (_08960_, _08959_, _08923_);
  nor _60397_ (_08961_, _08960_, _03474_);
  or _60398_ (_08962_, _08961_, _03437_);
  or _60399_ (_08963_, _08962_, _08958_);
  and _60400_ (_08964_, _06087_, _05208_);
  nor _60401_ (_08966_, _08964_, _08923_);
  nand _60402_ (_08967_, _08966_, _03437_);
  and _60403_ (_08968_, _08967_, _08963_);
  nor _60404_ (_08969_, _08968_, _03636_);
  and _60405_ (_08970_, _06305_, _05208_);
  or _60406_ (_08971_, _08923_, _04499_);
  nor _60407_ (_08972_, _08971_, _08970_);
  or _60408_ (_08973_, _08972_, _03769_);
  nor _60409_ (_08974_, _08973_, _08969_);
  nor _60410_ (_08975_, _08974_, _08926_);
  nor _60411_ (_08977_, _08975_, _04504_);
  not _60412_ (_08978_, _08923_);
  and _60413_ (_08979_, _08978_, _05281_);
  or _60414_ (_08980_, _08966_, _04505_);
  nor _60415_ (_08981_, _08980_, _08979_);
  nor _60416_ (_08982_, _08981_, _08977_);
  nor _60417_ (_08983_, _08982_, _03752_);
  or _60418_ (_08984_, _08979_, _03753_);
  nor _60419_ (_08985_, _08984_, _08928_);
  or _60420_ (_08986_, _08985_, _08983_);
  and _60421_ (_08988_, _08986_, _03759_);
  nor _60422_ (_08989_, _06304_, _08940_);
  nor _60423_ (_08990_, _08989_, _08923_);
  nor _60424_ (_08991_, _08990_, _03759_);
  or _60425_ (_08992_, _08991_, _08988_);
  and _60426_ (_08993_, _08992_, _04517_);
  nor _60427_ (_08994_, _06310_, _08940_);
  nor _60428_ (_08995_, _08994_, _08923_);
  nor _60429_ (_08996_, _08995_, _04517_);
  or _60430_ (_08997_, _08996_, _03790_);
  nor _60431_ (_08999_, _08997_, _08993_);
  and _60432_ (_09000_, _08936_, _03790_);
  or _60433_ (_09001_, _09000_, _03520_);
  nor _60434_ (_09002_, _09001_, _08999_);
  and _60435_ (_09003_, _05767_, _05208_);
  nor _60436_ (_09004_, _09003_, _08923_);
  nor _60437_ (_09005_, _09004_, _03521_);
  or _60438_ (_09006_, _09005_, _09002_);
  or _60439_ (_09007_, _09006_, _42967_);
  or _60440_ (_09008_, _42963_, \oc8051_golden_model_1.PCON [7]);
  and _60441_ (_09009_, _09008_, _41755_);
  and _60442_ (_40520_, _09009_, _09007_);
  not _60443_ (_09010_, \oc8051_golden_model_1.TCON [7]);
  nor _60444_ (_09011_, _05236_, _09010_);
  and _60445_ (_09012_, _06311_, _05236_);
  nor _60446_ (_09013_, _09012_, _09011_);
  nor _60447_ (_09014_, _09013_, _04501_);
  not _60448_ (_09015_, _05236_);
  nor _60449_ (_09016_, _09015_, _05176_);
  nor _60450_ (_09017_, _09016_, _09011_);
  and _60451_ (_09018_, _09017_, _07314_);
  nor _60452_ (_09019_, _05799_, _09010_);
  and _60453_ (_09020_, _05818_, _05799_);
  nor _60454_ (_09021_, _09020_, _09019_);
  nor _60455_ (_09022_, _09021_, _03513_);
  and _60456_ (_09023_, _05236_, \oc8051_golden_model_1.ACC [7]);
  nor _60457_ (_09024_, _09023_, _09011_);
  nor _60458_ (_09025_, _09024_, _04427_);
  nor _60459_ (_09026_, _04426_, _09010_);
  or _60460_ (_09027_, _09026_, _09025_);
  and _60461_ (_09028_, _09027_, _04444_);
  and _60462_ (_09029_, _05949_, _05236_);
  nor _60463_ (_09030_, _09029_, _09011_);
  nor _60464_ (_09031_, _09030_, _04444_);
  or _60465_ (_09032_, _09031_, _09028_);
  and _60466_ (_09033_, _09032_, _03517_);
  and _60467_ (_09034_, _05954_, _05799_);
  nor _60468_ (_09035_, _09034_, _09019_);
  nor _60469_ (_09036_, _09035_, _03517_);
  or _60470_ (_09037_, _09036_, _03568_);
  or _60471_ (_09038_, _09037_, _09033_);
  nand _60472_ (_09039_, _09017_, _03568_);
  and _60473_ (_09040_, _09039_, _09038_);
  and _60474_ (_09041_, _09040_, _03583_);
  nor _60475_ (_09042_, _09024_, _03583_);
  or _60476_ (_09043_, _09042_, _09041_);
  and _60477_ (_09044_, _09043_, _03513_);
  nor _60478_ (_09045_, _09044_, _09022_);
  nor _60479_ (_09046_, _09045_, _03505_);
  and _60480_ (_09047_, _05990_, _05799_);
  nor _60481_ (_09048_, _09047_, _09019_);
  nor _60482_ (_09049_, _09048_, _03506_);
  nor _60483_ (_09050_, _09049_, _09046_);
  nor _60484_ (_09051_, _09050_, _03499_);
  not _60485_ (_09052_, _05799_);
  nor _60486_ (_09053_, _06034_, _09052_);
  nor _60487_ (_09054_, _09053_, _09019_);
  nor _60488_ (_09055_, _09054_, _03500_);
  nor _60489_ (_09056_, _09055_, _07314_);
  not _60490_ (_09057_, _09056_);
  nor _60491_ (_09058_, _09057_, _09051_);
  nor _60492_ (_09059_, _09058_, _09018_);
  nor _60493_ (_09060_, _09059_, _03479_);
  and _60494_ (_09061_, _05935_, _05236_);
  nor _60495_ (_09062_, _09011_, _06044_);
  not _60496_ (_09063_, _09062_);
  nor _60497_ (_09064_, _09063_, _09061_);
  nor _60498_ (_09065_, _09064_, _03221_);
  not _60499_ (_09066_, _09065_);
  nor _60500_ (_09067_, _09066_, _09060_);
  nor _60501_ (_09068_, _06292_, _09015_);
  nor _60502_ (_09069_, _09068_, _09011_);
  nor _60503_ (_09070_, _09069_, _03474_);
  or _60504_ (_09071_, _09070_, _03437_);
  or _60505_ (_09072_, _09071_, _09067_);
  and _60506_ (_09073_, _06087_, _05236_);
  nor _60507_ (_09074_, _09073_, _09011_);
  nand _60508_ (_09075_, _09074_, _03437_);
  and _60509_ (_09076_, _09075_, _09072_);
  nor _60510_ (_09077_, _09076_, _03636_);
  and _60511_ (_09078_, _06305_, _05236_);
  or _60512_ (_09079_, _09011_, _04499_);
  nor _60513_ (_09080_, _09079_, _09078_);
  or _60514_ (_09081_, _09080_, _03769_);
  nor _60515_ (_09082_, _09081_, _09077_);
  nor _60516_ (_09083_, _09082_, _09014_);
  nor _60517_ (_09084_, _09083_, _04504_);
  not _60518_ (_09085_, _09011_);
  and _60519_ (_09086_, _09085_, _05281_);
  or _60520_ (_09087_, _09074_, _04505_);
  nor _60521_ (_09088_, _09087_, _09086_);
  nor _60522_ (_09089_, _09088_, _09084_);
  nor _60523_ (_09090_, _09089_, _03752_);
  or _60524_ (_09091_, _09086_, _03753_);
  nor _60525_ (_09092_, _09091_, _09024_);
  or _60526_ (_09093_, _09092_, _09090_);
  and _60527_ (_09094_, _09093_, _03759_);
  nor _60528_ (_09095_, _06304_, _09015_);
  nor _60529_ (_09096_, _09095_, _09011_);
  nor _60530_ (_09097_, _09096_, _03759_);
  or _60531_ (_09098_, _09097_, _09094_);
  and _60532_ (_09099_, _09098_, _04517_);
  nor _60533_ (_09100_, _06310_, _09015_);
  nor _60534_ (_09101_, _09100_, _09011_);
  nor _60535_ (_09102_, _09101_, _04517_);
  or _60536_ (_09103_, _09102_, _09099_);
  and _60537_ (_09104_, _09103_, _04192_);
  nor _60538_ (_09105_, _09030_, _04192_);
  or _60539_ (_09106_, _09105_, _09104_);
  and _60540_ (_09107_, _09106_, _03152_);
  nor _60541_ (_09108_, _09021_, _03152_);
  or _60542_ (_09109_, _09108_, _09107_);
  and _60543_ (_09110_, _09109_, _03521_);
  and _60544_ (_09111_, _05767_, _05236_);
  nor _60545_ (_09112_, _09111_, _09011_);
  nor _60546_ (_09113_, _09112_, _03521_);
  or _60547_ (_09114_, _09113_, _09110_);
  or _60548_ (_09115_, _09114_, _42967_);
  or _60549_ (_09116_, _42963_, \oc8051_golden_model_1.TCON [7]);
  and _60550_ (_09117_, _09116_, _41755_);
  and _60551_ (_40521_, _09117_, _09115_);
  not _60552_ (_09118_, \oc8051_golden_model_1.TL0 [7]);
  nor _60553_ (_09119_, _05258_, _09118_);
  and _60554_ (_09120_, _06311_, _05258_);
  nor _60555_ (_09121_, _09120_, _09119_);
  nor _60556_ (_09122_, _09121_, _04501_);
  and _60557_ (_09123_, _05258_, \oc8051_golden_model_1.ACC [7]);
  nor _60558_ (_09124_, _09123_, _09119_);
  nor _60559_ (_09125_, _09124_, _03583_);
  nor _60560_ (_09126_, _09124_, _04427_);
  nor _60561_ (_09127_, _04426_, _09118_);
  or _60562_ (_09128_, _09127_, _09126_);
  and _60563_ (_09129_, _09128_, _04444_);
  and _60564_ (_09130_, _05949_, _05258_);
  nor _60565_ (_09131_, _09130_, _09119_);
  nor _60566_ (_09132_, _09131_, _04444_);
  or _60567_ (_09133_, _09132_, _09129_);
  and _60568_ (_09134_, _09133_, _03983_);
  not _60569_ (_09135_, _05258_);
  nor _60570_ (_09136_, _09135_, _05176_);
  nor _60571_ (_09137_, _09136_, _09119_);
  nor _60572_ (_09138_, _09137_, _03983_);
  nor _60573_ (_09139_, _09138_, _09134_);
  nor _60574_ (_09140_, _09139_, _03575_);
  or _60575_ (_09141_, _09140_, _07314_);
  nor _60576_ (_09142_, _09141_, _09125_);
  and _60577_ (_09143_, _09137_, _07314_);
  nor _60578_ (_09144_, _09143_, _09142_);
  nor _60579_ (_09145_, _09144_, _03479_);
  and _60580_ (_09146_, _05935_, _05258_);
  nor _60581_ (_09147_, _09119_, _06044_);
  not _60582_ (_09148_, _09147_);
  nor _60583_ (_09149_, _09148_, _09146_);
  or _60584_ (_09150_, _09149_, _03221_);
  nor _60585_ (_09151_, _09150_, _09145_);
  nor _60586_ (_09152_, _06292_, _09135_);
  nor _60587_ (_09153_, _09152_, _09119_);
  nor _60588_ (_09154_, _09153_, _03474_);
  or _60589_ (_09155_, _09154_, _03437_);
  or _60590_ (_09156_, _09155_, _09151_);
  and _60591_ (_09157_, _06087_, _05258_);
  nor _60592_ (_09158_, _09157_, _09119_);
  nand _60593_ (_09159_, _09158_, _03437_);
  and _60594_ (_09160_, _09159_, _09156_);
  nor _60595_ (_09161_, _09160_, _03636_);
  and _60596_ (_09162_, _06305_, _05258_);
  or _60597_ (_09163_, _09119_, _04499_);
  nor _60598_ (_09164_, _09163_, _09162_);
  or _60599_ (_09165_, _09164_, _03769_);
  nor _60600_ (_09166_, _09165_, _09161_);
  nor _60601_ (_09167_, _09166_, _09122_);
  nor _60602_ (_09168_, _09167_, _04504_);
  not _60603_ (_09169_, _09119_);
  and _60604_ (_09170_, _09169_, _05281_);
  or _60605_ (_09171_, _09158_, _04505_);
  nor _60606_ (_09172_, _09171_, _09170_);
  nor _60607_ (_09173_, _09172_, _09168_);
  nor _60608_ (_09174_, _09173_, _03752_);
  or _60609_ (_09175_, _09170_, _03753_);
  or _60610_ (_09176_, _09175_, _09124_);
  and _60611_ (_09177_, _09176_, _03759_);
  not _60612_ (_09178_, _09177_);
  nor _60613_ (_09179_, _09178_, _09174_);
  nor _60614_ (_09180_, _06304_, _09135_);
  or _60615_ (_09181_, _09119_, _03759_);
  nor _60616_ (_09182_, _09181_, _09180_);
  or _60617_ (_09183_, _09182_, _03760_);
  nor _60618_ (_09184_, _09183_, _09179_);
  nor _60619_ (_09185_, _06310_, _09135_);
  nor _60620_ (_09186_, _09185_, _09119_);
  nor _60621_ (_09187_, _09186_, _04517_);
  or _60622_ (_09188_, _09187_, _03790_);
  nor _60623_ (_09189_, _09188_, _09184_);
  and _60624_ (_09190_, _09131_, _03790_);
  or _60625_ (_09191_, _09190_, _03520_);
  nor _60626_ (_09192_, _09191_, _09189_);
  and _60627_ (_09193_, _05767_, _05258_);
  nor _60628_ (_09194_, _09193_, _09119_);
  nor _60629_ (_09195_, _09194_, _03521_);
  or _60630_ (_09196_, _09195_, _09192_);
  or _60631_ (_09197_, _09196_, _42967_);
  or _60632_ (_09198_, _42963_, \oc8051_golden_model_1.TL0 [7]);
  and _60633_ (_09199_, _09198_, _41755_);
  and _60634_ (_40522_, _09199_, _09197_);
  not _60635_ (_09200_, \oc8051_golden_model_1.TL1 [7]);
  nor _60636_ (_09201_, _05242_, _09200_);
  and _60637_ (_09202_, _06311_, _05444_);
  nor _60638_ (_09203_, _09202_, _09201_);
  nor _60639_ (_09204_, _09203_, _04501_);
  not _60640_ (_09205_, _05444_);
  nor _60641_ (_09206_, _09205_, _05176_);
  nor _60642_ (_09207_, _09206_, _09201_);
  and _60643_ (_09208_, _09207_, _07314_);
  and _60644_ (_09209_, _05242_, \oc8051_golden_model_1.ACC [7]);
  nor _60645_ (_09210_, _09209_, _09201_);
  nor _60646_ (_09211_, _09210_, _03583_);
  nor _60647_ (_09212_, _09210_, _04427_);
  nor _60648_ (_09213_, _04426_, _09200_);
  or _60649_ (_09214_, _09213_, _09212_);
  and _60650_ (_09215_, _09214_, _04444_);
  and _60651_ (_09216_, _05949_, _05444_);
  nor _60652_ (_09217_, _09216_, _09201_);
  nor _60653_ (_09218_, _09217_, _04444_);
  or _60654_ (_09219_, _09218_, _09215_);
  and _60655_ (_09220_, _09219_, _03983_);
  nor _60656_ (_09221_, _09207_, _03983_);
  nor _60657_ (_09222_, _09221_, _09220_);
  nor _60658_ (_09223_, _09222_, _03575_);
  or _60659_ (_09224_, _09223_, _07314_);
  nor _60660_ (_09225_, _09224_, _09211_);
  nor _60661_ (_09226_, _09225_, _09208_);
  nor _60662_ (_09227_, _09226_, _03479_);
  nor _60663_ (_09228_, _09201_, _06044_);
  not _60664_ (_09229_, _05242_);
  or _60665_ (_09230_, _06004_, _09229_);
  and _60666_ (_09231_, _09230_, _09228_);
  or _60667_ (_09232_, _09231_, _03221_);
  nor _60668_ (_09233_, _09232_, _09227_);
  nor _60669_ (_09234_, _06292_, _09229_);
  nor _60670_ (_09235_, _09234_, _09201_);
  nor _60671_ (_09236_, _09235_, _03474_);
  or _60672_ (_09237_, _09236_, _03437_);
  or _60673_ (_09238_, _09237_, _09233_);
  and _60674_ (_09239_, _06087_, _05242_);
  nor _60675_ (_09240_, _09239_, _09201_);
  nand _60676_ (_09241_, _09240_, _03437_);
  and _60677_ (_09242_, _09241_, _09238_);
  nor _60678_ (_09243_, _09242_, _03636_);
  nand _60679_ (_09244_, _06305_, _05444_);
  nor _60680_ (_09245_, _09201_, _04499_);
  and _60681_ (_09246_, _09245_, _09244_);
  or _60682_ (_09247_, _09246_, _03769_);
  nor _60683_ (_09248_, _09247_, _09243_);
  nor _60684_ (_09249_, _09248_, _09204_);
  nor _60685_ (_09250_, _09249_, _04504_);
  not _60686_ (_09251_, _09201_);
  and _60687_ (_09252_, _09251_, _05281_);
  or _60688_ (_09253_, _09240_, _04505_);
  nor _60689_ (_09254_, _09253_, _09252_);
  nor _60690_ (_09255_, _09254_, _09250_);
  nor _60691_ (_09256_, _09255_, _03752_);
  or _60692_ (_09257_, _09252_, _03753_);
  or _60693_ (_09258_, _09257_, _09210_);
  and _60694_ (_09259_, _09258_, _03759_);
  not _60695_ (_09260_, _09259_);
  nor _60696_ (_09261_, _09260_, _09256_);
  or _60697_ (_09262_, _06304_, _09205_);
  nor _60698_ (_09263_, _09201_, _03759_);
  and _60699_ (_09264_, _09263_, _09262_);
  or _60700_ (_09265_, _09264_, _03760_);
  nor _60701_ (_09266_, _09265_, _09261_);
  nor _60702_ (_09267_, _06310_, _09205_);
  nor _60703_ (_09268_, _09267_, _09201_);
  nor _60704_ (_09269_, _09268_, _04517_);
  or _60705_ (_09270_, _09269_, _03790_);
  nor _60706_ (_09271_, _09270_, _09266_);
  and _60707_ (_09272_, _09217_, _03790_);
  or _60708_ (_09273_, _09272_, _03520_);
  nor _60709_ (_09274_, _09273_, _09271_);
  and _60710_ (_09275_, _05767_, _05242_);
  nor _60711_ (_09276_, _09275_, _09201_);
  nor _60712_ (_09277_, _09276_, _03521_);
  or _60713_ (_09278_, _09277_, _09274_);
  or _60714_ (_09279_, _09278_, _42967_);
  or _60715_ (_09280_, _42963_, \oc8051_golden_model_1.TL1 [7]);
  and _60716_ (_09281_, _09280_, _41755_);
  and _60717_ (_40523_, _09281_, _09279_);
  not _60718_ (_09282_, \oc8051_golden_model_1.TH0 [7]);
  nor _60719_ (_09283_, _05234_, _09282_);
  and _60720_ (_09284_, _06311_, _05234_);
  nor _60721_ (_09285_, _09284_, _09283_);
  nor _60722_ (_09286_, _09285_, _04501_);
  and _60723_ (_09287_, _05234_, \oc8051_golden_model_1.ACC [7]);
  nor _60724_ (_09288_, _09287_, _09283_);
  nor _60725_ (_09289_, _09288_, _03583_);
  nor _60726_ (_09290_, _09288_, _04427_);
  nor _60727_ (_09291_, _04426_, _09282_);
  or _60728_ (_09292_, _09291_, _09290_);
  and _60729_ (_09293_, _09292_, _04444_);
  and _60730_ (_09294_, _05949_, _05234_);
  nor _60731_ (_09295_, _09294_, _09283_);
  nor _60732_ (_09296_, _09295_, _04444_);
  or _60733_ (_09297_, _09296_, _09293_);
  and _60734_ (_09298_, _09297_, _03983_);
  not _60735_ (_09299_, _05234_);
  nor _60736_ (_09300_, _09299_, _05176_);
  nor _60737_ (_09301_, _09300_, _09283_);
  nor _60738_ (_09302_, _09301_, _03983_);
  nor _60739_ (_09303_, _09302_, _09298_);
  nor _60740_ (_09304_, _09303_, _03575_);
  or _60741_ (_09305_, _09304_, _07314_);
  nor _60742_ (_09306_, _09305_, _09289_);
  and _60743_ (_09307_, _09301_, _07314_);
  nor _60744_ (_09308_, _09307_, _09306_);
  nor _60745_ (_09309_, _09308_, _03479_);
  and _60746_ (_09310_, _05935_, _05234_);
  nor _60747_ (_09311_, _09283_, _06044_);
  not _60748_ (_09312_, _09311_);
  nor _60749_ (_09313_, _09312_, _09310_);
  or _60750_ (_09314_, _09313_, _03221_);
  nor _60751_ (_09315_, _09314_, _09309_);
  nor _60752_ (_09316_, _06292_, _09299_);
  nor _60753_ (_09317_, _09316_, _09283_);
  nor _60754_ (_09318_, _09317_, _03474_);
  or _60755_ (_09319_, _09318_, _03437_);
  or _60756_ (_09320_, _09319_, _09315_);
  and _60757_ (_09321_, _06087_, _05234_);
  nor _60758_ (_09322_, _09321_, _09283_);
  nand _60759_ (_09323_, _09322_, _03437_);
  and _60760_ (_09324_, _09323_, _09320_);
  nor _60761_ (_09325_, _09324_, _03636_);
  and _60762_ (_09326_, _06305_, _05234_);
  or _60763_ (_09327_, _09283_, _04499_);
  nor _60764_ (_09328_, _09327_, _09326_);
  or _60765_ (_09329_, _09328_, _03769_);
  nor _60766_ (_09330_, _09329_, _09325_);
  nor _60767_ (_09331_, _09330_, _09286_);
  nor _60768_ (_09332_, _09331_, _04504_);
  not _60769_ (_09333_, _09283_);
  and _60770_ (_09334_, _09333_, _05281_);
  or _60771_ (_09335_, _09322_, _04505_);
  nor _60772_ (_09336_, _09335_, _09334_);
  nor _60773_ (_09337_, _09336_, _09332_);
  nor _60774_ (_09338_, _09337_, _03752_);
  or _60775_ (_09339_, _09334_, _03753_);
  or _60776_ (_09340_, _09339_, _09288_);
  and _60777_ (_09341_, _09340_, _03759_);
  not _60778_ (_09342_, _09341_);
  nor _60779_ (_09343_, _09342_, _09338_);
  nor _60780_ (_09344_, _06304_, _09299_);
  or _60781_ (_09345_, _09283_, _03759_);
  nor _60782_ (_09346_, _09345_, _09344_);
  or _60783_ (_09347_, _09346_, _03760_);
  nor _60784_ (_09348_, _09347_, _09343_);
  nor _60785_ (_09349_, _06310_, _09299_);
  nor _60786_ (_09350_, _09349_, _09283_);
  nor _60787_ (_09351_, _09350_, _04517_);
  or _60788_ (_09352_, _09351_, _03790_);
  nor _60789_ (_09353_, _09352_, _09348_);
  and _60790_ (_09354_, _09295_, _03790_);
  or _60791_ (_09355_, _09354_, _03520_);
  nor _60792_ (_09356_, _09355_, _09353_);
  and _60793_ (_09357_, _05767_, _05234_);
  nor _60794_ (_09358_, _09357_, _09283_);
  nor _60795_ (_09359_, _09358_, _03521_);
  or _60796_ (_09360_, _09359_, _09356_);
  or _60797_ (_09361_, _09360_, _42967_);
  or _60798_ (_09362_, _42963_, \oc8051_golden_model_1.TH0 [7]);
  and _60799_ (_09363_, _09362_, _41755_);
  and _60800_ (_40524_, _09363_, _09361_);
  not _60801_ (_09364_, \oc8051_golden_model_1.TH1 [7]);
  nor _60802_ (_09365_, _05251_, _09364_);
  and _60803_ (_09366_, _06311_, _05251_);
  nor _60804_ (_09367_, _09366_, _09365_);
  nor _60805_ (_09368_, _09367_, _04501_);
  and _60806_ (_09369_, _05251_, \oc8051_golden_model_1.ACC [7]);
  nor _60807_ (_09370_, _09369_, _09365_);
  nor _60808_ (_09371_, _09370_, _03583_);
  nor _60809_ (_09372_, _09370_, _04427_);
  nor _60810_ (_09373_, _04426_, _09364_);
  or _60811_ (_09374_, _09373_, _09372_);
  and _60812_ (_09375_, _09374_, _04444_);
  and _60813_ (_09376_, _05949_, _05251_);
  nor _60814_ (_09377_, _09376_, _09365_);
  nor _60815_ (_09378_, _09377_, _04444_);
  or _60816_ (_09379_, _09378_, _09375_);
  and _60817_ (_09380_, _09379_, _03983_);
  not _60818_ (_09381_, _05251_);
  nor _60819_ (_09382_, _09381_, _05176_);
  nor _60820_ (_09383_, _09382_, _09365_);
  nor _60821_ (_09384_, _09383_, _03983_);
  nor _60822_ (_09385_, _09384_, _09380_);
  nor _60823_ (_09386_, _09385_, _03575_);
  or _60824_ (_09387_, _09386_, _07314_);
  nor _60825_ (_09388_, _09387_, _09371_);
  and _60826_ (_09389_, _09383_, _07314_);
  nor _60827_ (_09390_, _09389_, _09388_);
  nor _60828_ (_09391_, _09390_, _03479_);
  and _60829_ (_09392_, _05935_, _05251_);
  nor _60830_ (_09393_, _09365_, _06044_);
  not _60831_ (_09394_, _09393_);
  nor _60832_ (_09395_, _09394_, _09392_);
  or _60833_ (_09396_, _09395_, _03221_);
  nor _60834_ (_09397_, _09396_, _09391_);
  nor _60835_ (_09398_, _06292_, _09381_);
  nor _60836_ (_09399_, _09398_, _09365_);
  nor _60837_ (_09400_, _09399_, _03474_);
  or _60838_ (_09401_, _09400_, _03437_);
  or _60839_ (_09402_, _09401_, _09397_);
  and _60840_ (_09403_, _06087_, _05251_);
  nor _60841_ (_09404_, _09403_, _09365_);
  nand _60842_ (_09405_, _09404_, _03437_);
  and _60843_ (_09406_, _09405_, _09402_);
  nor _60844_ (_09407_, _09406_, _03636_);
  and _60845_ (_09408_, _06305_, _05251_);
  or _60846_ (_09409_, _09365_, _04499_);
  nor _60847_ (_09410_, _09409_, _09408_);
  or _60848_ (_09411_, _09410_, _03769_);
  nor _60849_ (_09412_, _09411_, _09407_);
  nor _60850_ (_09413_, _09412_, _09368_);
  nor _60851_ (_09414_, _09413_, _04504_);
  not _60852_ (_09415_, _09365_);
  and _60853_ (_09416_, _09415_, _05281_);
  or _60854_ (_09417_, _09404_, _04505_);
  nor _60855_ (_09418_, _09417_, _09416_);
  nor _60856_ (_09419_, _09418_, _09414_);
  nor _60857_ (_09420_, _09419_, _03752_);
  or _60858_ (_09421_, _09416_, _03753_);
  nor _60859_ (_09422_, _09421_, _09370_);
  or _60860_ (_09423_, _09422_, _09420_);
  and _60861_ (_09424_, _09423_, _03759_);
  nor _60862_ (_09425_, _06304_, _09381_);
  nor _60863_ (_09426_, _09425_, _09365_);
  nor _60864_ (_09427_, _09426_, _03759_);
  or _60865_ (_09428_, _09427_, _09424_);
  and _60866_ (_09429_, _09428_, _04517_);
  nor _60867_ (_09430_, _06310_, _09381_);
  nor _60868_ (_09431_, _09430_, _09365_);
  nor _60869_ (_09432_, _09431_, _04517_);
  or _60870_ (_09433_, _09432_, _03790_);
  nor _60871_ (_09434_, _09433_, _09429_);
  and _60872_ (_09435_, _09377_, _03790_);
  or _60873_ (_09436_, _09435_, _03520_);
  nor _60874_ (_09437_, _09436_, _09434_);
  and _60875_ (_09438_, _05767_, _05251_);
  nor _60876_ (_09439_, _09438_, _09365_);
  nor _60877_ (_09440_, _09439_, _03521_);
  or _60878_ (_09441_, _09440_, _09437_);
  or _60879_ (_09442_, _09441_, _42967_);
  or _60880_ (_09443_, _42963_, \oc8051_golden_model_1.TH1 [7]);
  and _60881_ (_09444_, _09443_, _41755_);
  and _60882_ (_40526_, _09444_, _09442_);
  not _60883_ (_09445_, \oc8051_golden_model_1.TMOD [7]);
  nor _60884_ (_09446_, _05254_, _09445_);
  and _60885_ (_09447_, _06311_, _05254_);
  nor _60886_ (_09448_, _09447_, _09446_);
  nor _60887_ (_09449_, _09448_, _04501_);
  and _60888_ (_09450_, _05254_, \oc8051_golden_model_1.ACC [7]);
  nor _60889_ (_09451_, _09450_, _09446_);
  nor _60890_ (_09452_, _09451_, _03583_);
  nor _60891_ (_09453_, _09451_, _04427_);
  nor _60892_ (_09454_, _04426_, _09445_);
  or _60893_ (_09455_, _09454_, _09453_);
  and _60894_ (_09456_, _09455_, _04444_);
  and _60895_ (_09457_, _05949_, _05254_);
  nor _60896_ (_09458_, _09457_, _09446_);
  nor _60897_ (_09459_, _09458_, _04444_);
  or _60898_ (_09460_, _09459_, _09456_);
  and _60899_ (_09461_, _09460_, _03983_);
  not _60900_ (_09462_, _05254_);
  nor _60901_ (_09463_, _09462_, _05176_);
  nor _60902_ (_09464_, _09463_, _09446_);
  nor _60903_ (_09465_, _09464_, _03983_);
  nor _60904_ (_09466_, _09465_, _09461_);
  nor _60905_ (_09467_, _09466_, _03575_);
  or _60906_ (_09468_, _09467_, _07314_);
  nor _60907_ (_09469_, _09468_, _09452_);
  and _60908_ (_09470_, _09464_, _07314_);
  nor _60909_ (_09471_, _09470_, _09469_);
  nor _60910_ (_09472_, _09471_, _03479_);
  and _60911_ (_09473_, _05935_, _05254_);
  nor _60912_ (_09474_, _09446_, _06044_);
  not _60913_ (_09475_, _09474_);
  nor _60914_ (_09476_, _09475_, _09473_);
  or _60915_ (_09477_, _09476_, _03221_);
  nor _60916_ (_09478_, _09477_, _09472_);
  nor _60917_ (_09479_, _06292_, _09462_);
  nor _60918_ (_09480_, _09479_, _09446_);
  nor _60919_ (_09481_, _09480_, _03474_);
  or _60920_ (_09482_, _09481_, _03437_);
  or _60921_ (_09483_, _09482_, _09478_);
  and _60922_ (_09484_, _06087_, _05254_);
  nor _60923_ (_09485_, _09484_, _09446_);
  nand _60924_ (_09486_, _09485_, _03437_);
  and _60925_ (_09487_, _09486_, _09483_);
  nor _60926_ (_09488_, _09487_, _03636_);
  and _60927_ (_09489_, _06305_, _05254_);
  or _60928_ (_09490_, _09446_, _04499_);
  nor _60929_ (_09491_, _09490_, _09489_);
  or _60930_ (_09492_, _09491_, _03769_);
  nor _60931_ (_09493_, _09492_, _09488_);
  nor _60932_ (_09494_, _09493_, _09449_);
  nor _60933_ (_09495_, _09494_, _04504_);
  not _60934_ (_09496_, _09446_);
  and _60935_ (_09497_, _09496_, _05281_);
  or _60936_ (_09498_, _09485_, _04505_);
  nor _60937_ (_09499_, _09498_, _09497_);
  nor _60938_ (_09500_, _09499_, _09495_);
  nor _60939_ (_09501_, _09500_, _03752_);
  or _60940_ (_09502_, _09497_, _03753_);
  nor _60941_ (_09503_, _09502_, _09451_);
  or _60942_ (_09504_, _09503_, _09501_);
  and _60943_ (_09505_, _09504_, _03759_);
  nor _60944_ (_09506_, _06304_, _09462_);
  nor _60945_ (_09507_, _09506_, _09446_);
  nor _60946_ (_09508_, _09507_, _03759_);
  or _60947_ (_09509_, _09508_, _09505_);
  and _60948_ (_09510_, _09509_, _04517_);
  nor _60949_ (_09511_, _06310_, _09462_);
  nor _60950_ (_09512_, _09511_, _09446_);
  nor _60951_ (_09513_, _09512_, _04517_);
  or _60952_ (_09514_, _09513_, _03790_);
  nor _60953_ (_09515_, _09514_, _09510_);
  and _60954_ (_09516_, _09458_, _03790_);
  or _60955_ (_09517_, _09516_, _03520_);
  nor _60956_ (_09518_, _09517_, _09515_);
  and _60957_ (_09519_, _05767_, _05254_);
  nor _60958_ (_09520_, _09519_, _09446_);
  nor _60959_ (_09521_, _09520_, _03521_);
  or _60960_ (_09522_, _09521_, _09518_);
  or _60961_ (_09523_, _09522_, _42967_);
  or _60962_ (_09524_, _42963_, \oc8051_golden_model_1.TMOD [7]);
  and _60963_ (_09525_, _09524_, _41755_);
  and _60964_ (_40527_, _09525_, _09523_);
  not _60965_ (_09526_, \oc8051_golden_model_1.IE [7]);
  nor _60966_ (_09527_, _05193_, _09526_);
  and _60967_ (_09528_, _06311_, _05193_);
  nor _60968_ (_09529_, _09528_, _09527_);
  nor _60969_ (_09530_, _09529_, _04501_);
  not _60970_ (_09531_, _05193_);
  nor _60971_ (_09532_, _09531_, _05176_);
  nor _60972_ (_09533_, _09532_, _09527_);
  and _60973_ (_09534_, _09533_, _07314_);
  nor _60974_ (_09535_, _05807_, _09526_);
  and _60975_ (_09536_, _05818_, _05807_);
  nor _60976_ (_09537_, _09536_, _09535_);
  nor _60977_ (_09538_, _09537_, _03513_);
  and _60978_ (_09539_, _05193_, \oc8051_golden_model_1.ACC [7]);
  nor _60979_ (_09540_, _09539_, _09527_);
  nor _60980_ (_09541_, _09540_, _04427_);
  nor _60981_ (_09543_, _04426_, _09526_);
  or _60982_ (_09544_, _09543_, _09541_);
  and _60983_ (_09545_, _09544_, _04444_);
  and _60984_ (_09546_, _05949_, _05193_);
  nor _60985_ (_09547_, _09546_, _09527_);
  nor _60986_ (_09548_, _09547_, _04444_);
  or _60987_ (_09549_, _09548_, _09545_);
  and _60988_ (_09550_, _09549_, _03517_);
  and _60989_ (_09551_, _05954_, _05807_);
  nor _60990_ (_09552_, _09551_, _09535_);
  nor _60991_ (_09553_, _09552_, _03517_);
  or _60992_ (_09554_, _09553_, _03568_);
  or _60993_ (_09555_, _09554_, _09550_);
  nand _60994_ (_09556_, _09533_, _03568_);
  and _60995_ (_09557_, _09556_, _09555_);
  and _60996_ (_09558_, _09557_, _03583_);
  nor _60997_ (_09559_, _09540_, _03583_);
  or _60998_ (_09560_, _09559_, _09558_);
  and _60999_ (_09561_, _09560_, _03513_);
  nor _61000_ (_09562_, _09561_, _09538_);
  nor _61001_ (_09564_, _09562_, _03505_);
  nor _61002_ (_09565_, _09535_, _05989_);
  or _61003_ (_09566_, _09552_, _03506_);
  nor _61004_ (_09567_, _09566_, _09565_);
  nor _61005_ (_09568_, _09567_, _09564_);
  nor _61006_ (_09569_, _09568_, _03499_);
  not _61007_ (_09570_, _05807_);
  nor _61008_ (_09571_, _06034_, _09570_);
  nor _61009_ (_09572_, _09571_, _09535_);
  nor _61010_ (_09573_, _09572_, _03500_);
  nor _61011_ (_09574_, _09573_, _07314_);
  not _61012_ (_09575_, _09574_);
  nor _61013_ (_09576_, _09575_, _09569_);
  nor _61014_ (_09577_, _09576_, _09534_);
  nor _61015_ (_09578_, _09577_, _03479_);
  and _61016_ (_09579_, _05935_, _05193_);
  nor _61017_ (_09580_, _09527_, _06044_);
  not _61018_ (_09581_, _09580_);
  nor _61019_ (_09582_, _09581_, _09579_);
  nor _61020_ (_09583_, _09582_, _03221_);
  not _61021_ (_09584_, _09583_);
  nor _61022_ (_09585_, _09584_, _09578_);
  nor _61023_ (_09586_, _06292_, _09531_);
  nor _61024_ (_09587_, _09586_, _09527_);
  nor _61025_ (_09588_, _09587_, _03474_);
  or _61026_ (_09589_, _09588_, _03437_);
  or _61027_ (_09590_, _09589_, _09585_);
  and _61028_ (_09591_, _06087_, _05193_);
  nor _61029_ (_09592_, _09591_, _09527_);
  nand _61030_ (_09593_, _09592_, _03437_);
  and _61031_ (_09594_, _09593_, _09590_);
  nor _61032_ (_09595_, _09594_, _03636_);
  and _61033_ (_09596_, _06305_, _05193_);
  or _61034_ (_09597_, _09527_, _04499_);
  nor _61035_ (_09598_, _09597_, _09596_);
  or _61036_ (_09599_, _09598_, _03769_);
  nor _61037_ (_09600_, _09599_, _09595_);
  nor _61038_ (_09601_, _09600_, _09530_);
  nor _61039_ (_09602_, _09601_, _04504_);
  not _61040_ (_09603_, _09527_);
  and _61041_ (_09604_, _09603_, _05281_);
  or _61042_ (_09605_, _09592_, _04505_);
  nor _61043_ (_09606_, _09605_, _09604_);
  nor _61044_ (_09607_, _09606_, _09602_);
  nor _61045_ (_09608_, _09607_, _03752_);
  or _61046_ (_09609_, _09604_, _03753_);
  nor _61047_ (_09610_, _09609_, _09540_);
  or _61048_ (_09611_, _09610_, _09608_);
  and _61049_ (_09612_, _09611_, _03759_);
  nor _61050_ (_09613_, _06304_, _09531_);
  nor _61051_ (_09614_, _09613_, _09527_);
  nor _61052_ (_09615_, _09614_, _03759_);
  or _61053_ (_09616_, _09615_, _09612_);
  and _61054_ (_09617_, _09616_, _04517_);
  nor _61055_ (_09618_, _06310_, _09531_);
  nor _61056_ (_09619_, _09618_, _09527_);
  nor _61057_ (_09620_, _09619_, _04517_);
  or _61058_ (_09621_, _09620_, _09617_);
  and _61059_ (_09622_, _09621_, _04192_);
  nor _61060_ (_09623_, _09547_, _04192_);
  or _61061_ (_09624_, _09623_, _09622_);
  and _61062_ (_09625_, _09624_, _03152_);
  nor _61063_ (_09626_, _09537_, _03152_);
  or _61064_ (_09627_, _09626_, _09625_);
  and _61065_ (_09628_, _09627_, _03521_);
  and _61066_ (_09629_, _05767_, _05193_);
  nor _61067_ (_09630_, _09629_, _09527_);
  nor _61068_ (_09631_, _09630_, _03521_);
  or _61069_ (_09632_, _09631_, _09628_);
  or _61070_ (_09633_, _09632_, _42967_);
  or _61071_ (_09634_, _42963_, \oc8051_golden_model_1.IE [7]);
  and _61072_ (_09635_, _09634_, _41755_);
  and _61073_ (_40528_, _09635_, _09633_);
  not _61074_ (_09636_, \oc8051_golden_model_1.IP [7]);
  nor _61075_ (_09637_, _05224_, _09636_);
  and _61076_ (_09638_, _06311_, _05224_);
  nor _61077_ (_09639_, _09638_, _09637_);
  nor _61078_ (_09640_, _09639_, _04501_);
  not _61079_ (_09641_, _05224_);
  nor _61080_ (_09642_, _09641_, _05176_);
  nor _61081_ (_09643_, _09642_, _09637_);
  and _61082_ (_09644_, _09643_, _07314_);
  nor _61083_ (_09645_, _05790_, _09636_);
  and _61084_ (_09646_, _05818_, _05790_);
  nor _61085_ (_09647_, _09646_, _09645_);
  nor _61086_ (_09648_, _09647_, _03513_);
  and _61087_ (_09649_, _05224_, \oc8051_golden_model_1.ACC [7]);
  nor _61088_ (_09650_, _09649_, _09637_);
  nor _61089_ (_09651_, _09650_, _04427_);
  nor _61090_ (_09652_, _04426_, _09636_);
  or _61091_ (_09653_, _09652_, _09651_);
  and _61092_ (_09654_, _09653_, _04444_);
  and _61093_ (_09655_, _05949_, _05224_);
  nor _61094_ (_09656_, _09655_, _09637_);
  nor _61095_ (_09657_, _09656_, _04444_);
  or _61096_ (_09658_, _09657_, _09654_);
  and _61097_ (_09659_, _09658_, _03517_);
  and _61098_ (_09660_, _05954_, _05790_);
  nor _61099_ (_09661_, _09660_, _09645_);
  nor _61100_ (_09662_, _09661_, _03517_);
  or _61101_ (_09663_, _09662_, _03568_);
  or _61102_ (_09664_, _09663_, _09659_);
  nand _61103_ (_09665_, _09643_, _03568_);
  and _61104_ (_09666_, _09665_, _09664_);
  and _61105_ (_09667_, _09666_, _03583_);
  nor _61106_ (_09668_, _09650_, _03583_);
  or _61107_ (_09669_, _09668_, _09667_);
  and _61108_ (_09670_, _09669_, _03513_);
  nor _61109_ (_09671_, _09670_, _09648_);
  nor _61110_ (_09672_, _09671_, _03505_);
  nor _61111_ (_09673_, _09645_, _05989_);
  or _61112_ (_09674_, _09661_, _03506_);
  nor _61113_ (_09675_, _09674_, _09673_);
  nor _61114_ (_09676_, _09675_, _09672_);
  nor _61115_ (_09677_, _09676_, _03499_);
  not _61116_ (_09678_, _05790_);
  nor _61117_ (_09679_, _06034_, _09678_);
  nor _61118_ (_09680_, _09679_, _09645_);
  nor _61119_ (_09681_, _09680_, _03500_);
  nor _61120_ (_09682_, _09681_, _07314_);
  not _61121_ (_09683_, _09682_);
  nor _61122_ (_09684_, _09683_, _09677_);
  nor _61123_ (_09685_, _09684_, _09644_);
  nor _61124_ (_09686_, _09685_, _03479_);
  and _61125_ (_09687_, _05935_, _05224_);
  nor _61126_ (_09688_, _09637_, _06044_);
  not _61127_ (_09689_, _09688_);
  nor _61128_ (_09690_, _09689_, _09687_);
  nor _61129_ (_09691_, _09690_, _03221_);
  not _61130_ (_09692_, _09691_);
  nor _61131_ (_09693_, _09692_, _09686_);
  nor _61132_ (_09694_, _06292_, _09641_);
  nor _61133_ (_09695_, _09694_, _09637_);
  nor _61134_ (_09696_, _09695_, _03474_);
  or _61135_ (_09697_, _09696_, _03437_);
  or _61136_ (_09698_, _09697_, _09693_);
  and _61137_ (_09699_, _06087_, _05224_);
  nor _61138_ (_09700_, _09699_, _09637_);
  nand _61139_ (_09701_, _09700_, _03437_);
  and _61140_ (_09702_, _09701_, _09698_);
  nor _61141_ (_09703_, _09702_, _03636_);
  and _61142_ (_09704_, _06305_, _05224_);
  or _61143_ (_09705_, _09637_, _04499_);
  nor _61144_ (_09706_, _09705_, _09704_);
  or _61145_ (_09707_, _09706_, _03769_);
  nor _61146_ (_09708_, _09707_, _09703_);
  nor _61147_ (_09709_, _09708_, _09640_);
  nor _61148_ (_09710_, _09709_, _04504_);
  not _61149_ (_09711_, _09637_);
  and _61150_ (_09712_, _09711_, _05281_);
  or _61151_ (_09713_, _09700_, _04505_);
  nor _61152_ (_09714_, _09713_, _09712_);
  nor _61153_ (_09715_, _09714_, _09710_);
  nor _61154_ (_09716_, _09715_, _03752_);
  or _61155_ (_09717_, _09712_, _03753_);
  nor _61156_ (_09718_, _09717_, _09650_);
  or _61157_ (_09719_, _09718_, _09716_);
  and _61158_ (_09720_, _09719_, _03759_);
  nor _61159_ (_09721_, _06304_, _09641_);
  nor _61160_ (_09722_, _09721_, _09637_);
  nor _61161_ (_09723_, _09722_, _03759_);
  or _61162_ (_09724_, _09723_, _09720_);
  and _61163_ (_09725_, _09724_, _04517_);
  nor _61164_ (_09726_, _06310_, _09641_);
  nor _61165_ (_09727_, _09726_, _09637_);
  nor _61166_ (_09728_, _09727_, _04517_);
  or _61167_ (_09729_, _09728_, _09725_);
  and _61168_ (_09730_, _09729_, _04192_);
  nor _61169_ (_09731_, _09656_, _04192_);
  or _61170_ (_09732_, _09731_, _09730_);
  and _61171_ (_09733_, _09732_, _03152_);
  nor _61172_ (_09734_, _09647_, _03152_);
  or _61173_ (_09735_, _09734_, _09733_);
  and _61174_ (_09736_, _09735_, _03521_);
  and _61175_ (_09737_, _05767_, _05224_);
  nor _61176_ (_09738_, _09737_, _09637_);
  nor _61177_ (_09739_, _09738_, _03521_);
  or _61178_ (_09740_, _09739_, _09736_);
  or _61179_ (_09741_, _09740_, _42967_);
  or _61180_ (_09742_, _42963_, \oc8051_golden_model_1.IP [7]);
  and _61181_ (_09743_, _09742_, _41755_);
  and _61182_ (_40529_, _09743_, _09741_);
  or _61183_ (_09744_, _42963_, \oc8051_golden_model_1.DPL [7]);
  and _61184_ (_09745_, _09744_, _41755_);
  not _61185_ (_09746_, \oc8051_golden_model_1.DPL [7]);
  nor _61186_ (_09747_, _05272_, _09746_);
  and _61187_ (_09748_, _06311_, _05272_);
  or _61188_ (_09749_, _09748_, _09747_);
  and _61189_ (_09750_, _09749_, _03769_);
  not _61190_ (_09751_, _05272_);
  nor _61191_ (_09752_, _09751_, _05176_);
  or _61192_ (_09753_, _09752_, _09747_);
  or _61193_ (_09754_, _09753_, _06039_);
  not _61194_ (_09755_, _03632_);
  and _61195_ (_09756_, _05949_, _05272_);
  or _61196_ (_09757_, _09756_, _09747_);
  or _61197_ (_09758_, _09757_, _04444_);
  and _61198_ (_09759_, _05272_, \oc8051_golden_model_1.ACC [7]);
  or _61199_ (_09760_, _09759_, _09747_);
  and _61200_ (_09761_, _09760_, _04426_);
  nor _61201_ (_09762_, _04426_, _09746_);
  or _61202_ (_09763_, _09762_, _03570_);
  or _61203_ (_09764_, _09763_, _09761_);
  and _61204_ (_09765_, _09764_, _03983_);
  and _61205_ (_09766_, _09765_, _09758_);
  and _61206_ (_09767_, _09753_, _03568_);
  or _61207_ (_09768_, _09767_, _03575_);
  or _61208_ (_09769_, _09768_, _09766_);
  nor _61209_ (_09770_, _03229_, _03212_);
  not _61210_ (_09771_, _09770_);
  or _61211_ (_09772_, _09760_, _03583_);
  and _61212_ (_09773_, _09772_, _09771_);
  and _61213_ (_09774_, _09773_, _09769_);
  and _61214_ (_09775_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and _61215_ (_09776_, _09775_, \oc8051_golden_model_1.DPL [2]);
  and _61216_ (_09777_, _09776_, \oc8051_golden_model_1.DPL [3]);
  and _61217_ (_09778_, _09777_, \oc8051_golden_model_1.DPL [4]);
  and _61218_ (_09779_, _09778_, \oc8051_golden_model_1.DPL [5]);
  and _61219_ (_09780_, _09779_, \oc8051_golden_model_1.DPL [6]);
  nor _61220_ (_09781_, _09780_, \oc8051_golden_model_1.DPL [7]);
  and _61221_ (_09782_, _09780_, \oc8051_golden_model_1.DPL [7]);
  nor _61222_ (_09783_, _09782_, _09781_);
  and _61223_ (_09784_, _09783_, _09770_);
  or _61224_ (_09785_, _09784_, _09774_);
  and _61225_ (_09786_, _09785_, _09755_);
  nor _61226_ (_09787_, _06086_, _09755_);
  or _61227_ (_09788_, _09787_, _07314_);
  or _61228_ (_09789_, _09788_, _09786_);
  and _61229_ (_09790_, _09789_, _09754_);
  or _61230_ (_09791_, _09790_, _03479_);
  and _61231_ (_09792_, _05935_, _05272_);
  or _61232_ (_09793_, _09747_, _06044_);
  or _61233_ (_09794_, _09793_, _09792_);
  and _61234_ (_09795_, _09794_, _03474_);
  and _61235_ (_09796_, _09795_, _09791_);
  nor _61236_ (_09797_, _06292_, _09751_);
  or _61237_ (_09798_, _09797_, _09747_);
  and _61238_ (_09799_, _09798_, _03221_);
  or _61239_ (_09800_, _09799_, _03437_);
  or _61240_ (_09801_, _09800_, _09796_);
  and _61241_ (_09802_, _06087_, _05272_);
  or _61242_ (_09803_, _09802_, _09747_);
  or _61243_ (_09804_, _09803_, _03438_);
  and _61244_ (_09805_, _09804_, _09801_);
  or _61245_ (_09806_, _09805_, _03636_);
  and _61246_ (_09807_, _06305_, _05272_);
  or _61247_ (_09808_, _09807_, _09747_);
  or _61248_ (_09809_, _09808_, _04499_);
  and _61249_ (_09810_, _09809_, _04501_);
  and _61250_ (_09811_, _09810_, _09806_);
  or _61251_ (_09812_, _09811_, _09750_);
  and _61252_ (_09813_, _09812_, _05769_);
  or _61253_ (_09814_, _09747_, _05282_);
  and _61254_ (_09815_, _09814_, _03754_);
  and _61255_ (_09816_, _09815_, _09803_);
  or _61256_ (_09817_, _09816_, _09813_);
  and _61257_ (_09818_, _09817_, _03753_);
  and _61258_ (_09819_, _09760_, _03752_);
  and _61259_ (_09820_, _09819_, _09814_);
  or _61260_ (_09821_, _09820_, _03758_);
  or _61261_ (_09822_, _09821_, _09818_);
  nor _61262_ (_09823_, _06304_, _09751_);
  or _61263_ (_09824_, _09747_, _03759_);
  or _61264_ (_09825_, _09824_, _09823_);
  and _61265_ (_09826_, _09825_, _04517_);
  and _61266_ (_09827_, _09826_, _09822_);
  nor _61267_ (_09828_, _06310_, _09751_);
  or _61268_ (_09829_, _09828_, _09747_);
  and _61269_ (_09830_, _09829_, _03760_);
  or _61270_ (_09831_, _09830_, _03790_);
  or _61271_ (_09832_, _09831_, _09827_);
  or _61272_ (_09833_, _09757_, _04192_);
  and _61273_ (_09834_, _09833_, _03521_);
  and _61274_ (_09835_, _09834_, _09832_);
  and _61275_ (_09836_, _05767_, _05272_);
  or _61276_ (_09837_, _09836_, _09747_);
  and _61277_ (_09838_, _09837_, _03520_);
  or _61278_ (_09839_, _09838_, _42967_);
  or _61279_ (_09840_, _09839_, _09835_);
  and _61280_ (_40530_, _09840_, _09745_);
  or _61281_ (_09841_, _42963_, \oc8051_golden_model_1.DPH [7]);
  and _61282_ (_09842_, _09841_, _41755_);
  not _61283_ (_09843_, \oc8051_golden_model_1.DPH [7]);
  nor _61284_ (_09844_, _05266_, _09843_);
  and _61285_ (_09845_, _06311_, _05266_);
  or _61286_ (_09846_, _09845_, _09844_);
  and _61287_ (_09847_, _09846_, _03769_);
  not _61288_ (_09848_, _05266_);
  nor _61289_ (_09849_, _09848_, _05176_);
  or _61290_ (_09850_, _09849_, _09844_);
  or _61291_ (_09851_, _09850_, _06039_);
  and _61292_ (_09852_, _05949_, _05266_);
  or _61293_ (_09853_, _09852_, _09844_);
  or _61294_ (_09854_, _09853_, _04444_);
  and _61295_ (_09855_, _05266_, \oc8051_golden_model_1.ACC [7]);
  or _61296_ (_09856_, _09855_, _09844_);
  and _61297_ (_09857_, _09856_, _04426_);
  nor _61298_ (_09858_, _04426_, _09843_);
  or _61299_ (_09859_, _09858_, _03570_);
  or _61300_ (_09860_, _09859_, _09857_);
  and _61301_ (_09861_, _09860_, _03983_);
  and _61302_ (_09862_, _09861_, _09854_);
  and _61303_ (_09863_, _09850_, _03568_);
  or _61304_ (_09864_, _09863_, _03575_);
  or _61305_ (_09865_, _09864_, _09862_);
  or _61306_ (_09866_, _09856_, _03583_);
  and _61307_ (_09867_, _09866_, _09771_);
  and _61308_ (_09868_, _09867_, _09865_);
  and _61309_ (_09869_, _09782_, \oc8051_golden_model_1.DPH [0]);
  and _61310_ (_09870_, _09869_, \oc8051_golden_model_1.DPH [1]);
  and _61311_ (_09871_, _09870_, \oc8051_golden_model_1.DPH [2]);
  and _61312_ (_09872_, _09871_, \oc8051_golden_model_1.DPH [3]);
  and _61313_ (_09873_, _09872_, \oc8051_golden_model_1.DPH [4]);
  and _61314_ (_09874_, _09873_, \oc8051_golden_model_1.DPH [5]);
  nand _61315_ (_09875_, _09874_, \oc8051_golden_model_1.DPH [6]);
  or _61316_ (_09876_, _09875_, _09843_);
  nand _61317_ (_09877_, _09875_, _09843_);
  and _61318_ (_09878_, _09877_, _09770_);
  and _61319_ (_09879_, _09878_, _09876_);
  or _61320_ (_09880_, _09879_, _09868_);
  and _61321_ (_09881_, _09880_, _09755_);
  and _61322_ (_09882_, _03632_, _03401_);
  or _61323_ (_09883_, _09882_, _07314_);
  or _61324_ (_09884_, _09883_, _09881_);
  and _61325_ (_09885_, _09884_, _09851_);
  or _61326_ (_09886_, _09885_, _03479_);
  and _61327_ (_09887_, _05935_, _05266_);
  or _61328_ (_09888_, _09844_, _06044_);
  or _61329_ (_09889_, _09888_, _09887_);
  and _61330_ (_09890_, _09889_, _03474_);
  and _61331_ (_09891_, _09890_, _09886_);
  nor _61332_ (_09892_, _06292_, _09848_);
  or _61333_ (_09893_, _09892_, _09844_);
  and _61334_ (_09894_, _09893_, _03221_);
  or _61335_ (_09895_, _09894_, _03437_);
  or _61336_ (_09896_, _09895_, _09891_);
  and _61337_ (_09897_, _06087_, _05266_);
  or _61338_ (_09898_, _09897_, _09844_);
  or _61339_ (_09899_, _09898_, _03438_);
  and _61340_ (_09900_, _09899_, _09896_);
  or _61341_ (_09901_, _09900_, _03636_);
  and _61342_ (_09902_, _06305_, _05266_);
  or _61343_ (_09903_, _09902_, _09844_);
  or _61344_ (_09904_, _09903_, _04499_);
  and _61345_ (_09905_, _09904_, _04501_);
  and _61346_ (_09906_, _09905_, _09901_);
  or _61347_ (_09907_, _09906_, _09847_);
  and _61348_ (_09908_, _09907_, _05769_);
  or _61349_ (_09909_, _09844_, _05282_);
  and _61350_ (_09910_, _09909_, _03754_);
  and _61351_ (_09911_, _09910_, _09898_);
  or _61352_ (_09912_, _09911_, _09908_);
  and _61353_ (_09913_, _09912_, _03753_);
  and _61354_ (_09914_, _09856_, _03752_);
  and _61355_ (_09915_, _09914_, _09909_);
  or _61356_ (_09916_, _09915_, _03758_);
  or _61357_ (_09917_, _09916_, _09913_);
  nor _61358_ (_09918_, _06304_, _09848_);
  or _61359_ (_09919_, _09844_, _03759_);
  or _61360_ (_09920_, _09919_, _09918_);
  and _61361_ (_09921_, _09920_, _04517_);
  and _61362_ (_09922_, _09921_, _09917_);
  nor _61363_ (_09923_, _06310_, _09848_);
  or _61364_ (_09924_, _09923_, _09844_);
  and _61365_ (_09925_, _09924_, _03760_);
  or _61366_ (_09926_, _09925_, _03790_);
  or _61367_ (_09927_, _09926_, _09922_);
  or _61368_ (_09928_, _09853_, _04192_);
  and _61369_ (_09929_, _09928_, _03521_);
  and _61370_ (_09930_, _09929_, _09927_);
  and _61371_ (_09931_, _05767_, _05266_);
  or _61372_ (_09932_, _09931_, _09844_);
  and _61373_ (_09933_, _09932_, _03520_);
  or _61374_ (_09934_, _09933_, _42967_);
  or _61375_ (_09935_, _09934_, _09930_);
  and _61376_ (_40532_, _09935_, _09842_);
  nor _61377_ (_09936_, _08597_, _03524_);
  not _61378_ (_09937_, _09936_);
  not _61379_ (_09938_, _02874_);
  and _61380_ (_09939_, _05837_, _09938_);
  and _61381_ (_09940_, _09939_, \oc8051_golden_model_1.PC [7]);
  and _61382_ (_09941_, _09940_, _06740_);
  and _61383_ (_09942_, _09941_, _06737_);
  and _61384_ (_09943_, _09942_, \oc8051_golden_model_1.PC [14]);
  and _61385_ (_09944_, _09943_, _06736_);
  nor _61386_ (_09945_, _09943_, _06736_);
  or _61387_ (_09946_, _09945_, _09944_);
  and _61388_ (_09947_, _04712_, _04002_);
  and _61389_ (_09948_, _09947_, _07777_);
  or _61390_ (_09949_, _09948_, _04178_);
  or _61391_ (_09950_, _09949_, _09946_);
  and _61392_ (_09951_, _08495_, _07830_);
  or _61393_ (_09952_, _09951_, _09946_);
  nor _61394_ (_09953_, _08456_, _04319_);
  and _61395_ (_09954_, _03476_, _03182_);
  nor _61396_ (_09955_, _08469_, _09954_);
  and _61397_ (_09956_, _09955_, _09953_);
  or _61398_ (_09957_, _09956_, _09946_);
  and _61399_ (_09958_, _03191_, _03150_);
  not _61400_ (_09959_, _09958_);
  nor _61401_ (_09960_, _03752_, _03192_);
  or _61402_ (_09961_, _09960_, _06746_);
  and _61403_ (_09962_, _09961_, _09959_);
  and _61404_ (_09963_, _05839_, \oc8051_golden_model_1.PC [8]);
  and _61405_ (_09964_, _09963_, \oc8051_golden_model_1.PC [9]);
  and _61406_ (_09965_, _09964_, \oc8051_golden_model_1.PC [10]);
  and _61407_ (_09966_, _09965_, \oc8051_golden_model_1.PC [11]);
  and _61408_ (_09967_, _09966_, \oc8051_golden_model_1.PC [12]);
  and _61409_ (_09968_, _09967_, \oc8051_golden_model_1.PC [13]);
  and _61410_ (_09969_, _09968_, \oc8051_golden_model_1.PC [14]);
  nor _61411_ (_09970_, _09968_, \oc8051_golden_model_1.PC [14]);
  nor _61412_ (_09971_, _09970_, _09969_);
  and _61413_ (_09972_, _09971_, _03401_);
  nor _61414_ (_09973_, _09971_, _03401_);
  nor _61415_ (_09974_, _09973_, _09972_);
  not _61416_ (_09975_, _09974_);
  nor _61417_ (_09976_, _09967_, \oc8051_golden_model_1.PC [13]);
  nor _61418_ (_09977_, _09976_, _09968_);
  and _61419_ (_09978_, _09977_, _03401_);
  nor _61420_ (_09979_, _09977_, _03401_);
  nor _61421_ (_09980_, _09966_, \oc8051_golden_model_1.PC [12]);
  nor _61422_ (_09981_, _09980_, _09967_);
  and _61423_ (_09982_, _09981_, _03401_);
  nor _61424_ (_09983_, _09965_, \oc8051_golden_model_1.PC [11]);
  nor _61425_ (_09984_, _09983_, _09966_);
  and _61426_ (_09985_, _09984_, _03401_);
  nor _61427_ (_09986_, _09984_, _03401_);
  nor _61428_ (_09987_, _09986_, _09985_);
  nor _61429_ (_09988_, _09964_, \oc8051_golden_model_1.PC [10]);
  nor _61430_ (_09989_, _09988_, _09965_);
  and _61431_ (_09990_, _09989_, _03401_);
  nor _61432_ (_09991_, _09989_, _03401_);
  nor _61433_ (_09992_, _09991_, _09990_);
  and _61434_ (_09993_, _09992_, _09987_);
  nor _61435_ (_09994_, _09963_, \oc8051_golden_model_1.PC [9]);
  nor _61436_ (_09995_, _09994_, _09964_);
  and _61437_ (_09996_, _09995_, _03401_);
  nor _61438_ (_09997_, _09995_, _03401_);
  nor _61439_ (_09998_, _09997_, _09996_);
  and _61440_ (_09999_, _05841_, _03401_);
  nor _61441_ (_10000_, _05841_, _03401_);
  and _61442_ (_10001_, _05836_, _03278_);
  nor _61443_ (_10002_, _10001_, \oc8051_golden_model_1.PC [6]);
  nor _61444_ (_10003_, _10002_, _05838_);
  not _61445_ (_10004_, _10003_);
  nor _61446_ (_10005_, _10004_, _03561_);
  and _61447_ (_10006_, _10004_, _03561_);
  nor _61448_ (_10007_, _10006_, _10005_);
  and _61449_ (_10008_, _03278_, \oc8051_golden_model_1.PC [4]);
  nor _61450_ (_10009_, _10008_, \oc8051_golden_model_1.PC [5]);
  nor _61451_ (_10010_, _10009_, _10001_);
  not _61452_ (_10011_, _10010_);
  nor _61453_ (_10012_, _10011_, _03834_);
  and _61454_ (_10013_, _10011_, _03834_);
  nor _61455_ (_10014_, _03278_, \oc8051_golden_model_1.PC [4]);
  nor _61456_ (_10015_, _10014_, _10008_);
  not _61457_ (_10016_, _10015_);
  nor _61458_ (_10017_, _10016_, _04249_);
  nor _61459_ (_10018_, _03432_, _03675_);
  and _61460_ (_10019_, _03432_, _03675_);
  nor _61461_ (_10020_, _03877_, _03626_);
  nor _61462_ (_10021_, _04284_, \oc8051_golden_model_1.PC [1]);
  nor _61463_ (_10022_, _03471_, _02887_);
  and _61464_ (_10023_, _04284_, \oc8051_golden_model_1.PC [1]);
  nor _61465_ (_10024_, _10023_, _10021_);
  and _61466_ (_10025_, _10024_, _10022_);
  nor _61467_ (_10026_, _10025_, _10021_);
  and _61468_ (_10027_, _03877_, _03626_);
  nor _61469_ (_10028_, _10027_, _10020_);
  not _61470_ (_10029_, _10028_);
  nor _61471_ (_10030_, _10029_, _10026_);
  nor _61472_ (_10031_, _10030_, _10020_);
  nor _61473_ (_10032_, _10031_, _10019_);
  nor _61474_ (_10033_, _10032_, _10018_);
  not _61475_ (_10034_, _10033_);
  and _61476_ (_10035_, _10016_, _04249_);
  nor _61477_ (_10036_, _10035_, _10017_);
  and _61478_ (_10037_, _10036_, _10034_);
  nor _61479_ (_10038_, _10037_, _10017_);
  nor _61480_ (_10039_, _10038_, _10013_);
  nor _61481_ (_10040_, _10039_, _10012_);
  not _61482_ (_10041_, _10040_);
  and _61483_ (_10042_, _10041_, _10007_);
  nor _61484_ (_10043_, _10042_, _10005_);
  nor _61485_ (_10044_, _10043_, _10000_);
  or _61486_ (_10045_, _10044_, _09999_);
  nor _61487_ (_10046_, _05839_, \oc8051_golden_model_1.PC [8]);
  nor _61488_ (_10047_, _10046_, _09963_);
  and _61489_ (_10048_, _10047_, _03401_);
  nor _61490_ (_10049_, _10047_, _03401_);
  nor _61491_ (_10050_, _10049_, _10048_);
  and _61492_ (_10051_, _10050_, _10045_);
  and _61493_ (_10052_, _10051_, _09998_);
  and _61494_ (_10053_, _10052_, _09993_);
  nor _61495_ (_10054_, _10048_, _09996_);
  not _61496_ (_10055_, _10054_);
  and _61497_ (_10056_, _10055_, _09993_);
  or _61498_ (_10057_, _10056_, _09990_);
  or _61499_ (_10058_, _10057_, _10053_);
  nor _61500_ (_10059_, _10058_, _09985_);
  nor _61501_ (_10060_, _09981_, _03401_);
  nor _61502_ (_10061_, _10060_, _09982_);
  not _61503_ (_10062_, _10061_);
  nor _61504_ (_10063_, _10062_, _10059_);
  nor _61505_ (_10064_, _10063_, _09982_);
  nor _61506_ (_10065_, _10064_, _09979_);
  nor _61507_ (_10066_, _10065_, _09978_);
  nor _61508_ (_10067_, _10066_, _09975_);
  nor _61509_ (_10068_, _10067_, _09972_);
  nor _61510_ (_10069_, _06746_, _03401_);
  and _61511_ (_10070_, _06746_, _03401_);
  nor _61512_ (_10071_, _10070_, _10069_);
  and _61513_ (_10072_, _10071_, _10068_);
  nor _61514_ (_10073_, _10071_, _10068_);
  or _61515_ (_10074_, _10073_, _10072_);
  or _61516_ (_10075_, _10074_, _08698_);
  and _61517_ (_10076_, _03188_, _03150_);
  not _61518_ (_10077_, _08698_);
  or _61519_ (_10078_, _10077_, _06746_);
  and _61520_ (_10079_, _10078_, _10076_);
  and _61521_ (_10080_, _10079_, _10075_);
  nor _61522_ (_10081_, _07328_, _03231_);
  and _61523_ (_10082_, _06754_, _03221_);
  nor _61524_ (_10083_, _03229_, _03199_);
  not _61525_ (_10084_, _10083_);
  not _61526_ (_10085_, _03638_);
  and _61527_ (_10086_, _06478_, _03472_);
  not _61528_ (_10087_, _10086_);
  or _61529_ (_10088_, _05935_, _05215_);
  or _61530_ (_10089_, _06713_, _03561_);
  and _61531_ (_10090_, _10089_, _10088_);
  or _61532_ (_10091_, _06388_, _04956_);
  or _61533_ (_10092_, _06616_, _05190_);
  and _61534_ (_10093_, _10092_, _10091_);
  and _61535_ (_10094_, _10093_, _10090_);
  or _61536_ (_10095_, _06721_, _03834_);
  or _61537_ (_10096_, _06722_, _04249_);
  and _61538_ (_10097_, _10096_, _10095_);
  or _61539_ (_10098_, _06661_, _05182_);
  and _61540_ (_10099_, _10098_, _06005_);
  and _61541_ (_10100_, _10099_, _10097_);
  and _61542_ (_10101_, _10100_, _10094_);
  or _61543_ (_10102_, _06717_, _03432_);
  or _61544_ (_10103_, _06524_, _03563_);
  and _61545_ (_10104_, _10103_, _10102_);
  or _61546_ (_10105_, _06569_, _04965_);
  or _61547_ (_10106_, _06718_, _03877_);
  and _61548_ (_10107_, _10106_, _10105_);
  and _61549_ (_10108_, _10107_, _10104_);
  or _61550_ (_10109_, _06478_, _03472_);
  or _61551_ (_10110_, _06714_, _04284_);
  or _61552_ (_10111_, _06433_, _04548_);
  and _61553_ (_10112_, _10111_, _10110_);
  and _61554_ (_10113_, _10112_, _10109_);
  and _61555_ (_10114_, _10113_, _10108_);
  and _61556_ (_10115_, _10114_, _10101_);
  and _61557_ (_10116_, _10115_, _10087_);
  and _61558_ (_10117_, _10116_, _06754_);
  and _61559_ (_10118_, _06677_, \oc8051_golden_model_1.PC [8]);
  and _61560_ (_10119_, _10118_, \oc8051_golden_model_1.PC [9]);
  and _61561_ (_10120_, _10119_, \oc8051_golden_model_1.PC [10]);
  and _61562_ (_10121_, _10120_, \oc8051_golden_model_1.PC [11]);
  and _61563_ (_10122_, _10121_, \oc8051_golden_model_1.PC [12]);
  and _61564_ (_10123_, _10122_, \oc8051_golden_model_1.PC [13]);
  and _61565_ (_10124_, _10123_, \oc8051_golden_model_1.PC [14]);
  nor _61566_ (_10125_, _10123_, \oc8051_golden_model_1.PC [14]);
  nor _61567_ (_10126_, _10125_, _10124_);
  not _61568_ (_10127_, _10126_);
  nor _61569_ (_10128_, _10127_, _06086_);
  and _61570_ (_10129_, _10127_, _06086_);
  nor _61571_ (_10130_, _10129_, _10128_);
  not _61572_ (_10131_, _10130_);
  nor _61573_ (_10132_, _10122_, \oc8051_golden_model_1.PC [13]);
  nor _61574_ (_10133_, _10132_, _10123_);
  not _61575_ (_10134_, _10133_);
  nor _61576_ (_10135_, _10134_, _06086_);
  and _61577_ (_10136_, _10134_, _06086_);
  nor _61578_ (_10137_, _10121_, \oc8051_golden_model_1.PC [12]);
  nor _61579_ (_10138_, _10137_, _10122_);
  not _61580_ (_10139_, _10138_);
  nor _61581_ (_10140_, _10139_, _06086_);
  nor _61582_ (_10141_, _10119_, \oc8051_golden_model_1.PC [10]);
  nor _61583_ (_10142_, _10141_, _10120_);
  not _61584_ (_10143_, _10142_);
  nor _61585_ (_10144_, _10143_, _06086_);
  not _61586_ (_10145_, _10144_);
  nor _61587_ (_10146_, _10120_, \oc8051_golden_model_1.PC [11]);
  nor _61588_ (_10147_, _10146_, _10121_);
  not _61589_ (_10148_, _10147_);
  nor _61590_ (_10149_, _10148_, _06086_);
  and _61591_ (_10150_, _10148_, _06086_);
  nor _61592_ (_10151_, _10150_, _10149_);
  and _61593_ (_10152_, _10143_, _06086_);
  nor _61594_ (_10153_, _10152_, _10144_);
  and _61595_ (_10154_, _10153_, _10151_);
  nor _61596_ (_10155_, _10118_, \oc8051_golden_model_1.PC [9]);
  nor _61597_ (_10156_, _10155_, _10119_);
  not _61598_ (_10157_, _10156_);
  nor _61599_ (_10158_, _10157_, _06086_);
  and _61600_ (_10159_, _10157_, _06086_);
  nor _61601_ (_10160_, _10159_, _10158_);
  nor _61602_ (_10161_, _06680_, _06086_);
  and _61603_ (_10162_, _06680_, _06086_);
  and _61604_ (_10163_, _06675_, _05836_);
  nor _61605_ (_10164_, _10163_, \oc8051_golden_model_1.PC [6]);
  nor _61606_ (_10165_, _10164_, _06676_);
  not _61607_ (_10166_, _10165_);
  nor _61608_ (_10167_, _10166_, _06132_);
  and _61609_ (_10168_, _10166_, _06132_);
  nor _61610_ (_10169_, _10168_, _10167_);
  not _61611_ (_10170_, _10169_);
  and _61612_ (_10171_, _06675_, \oc8051_golden_model_1.PC [4]);
  nor _61613_ (_10172_, _10171_, \oc8051_golden_model_1.PC [5]);
  nor _61614_ (_10173_, _10172_, _10163_);
  not _61615_ (_10174_, _10173_);
  nor _61616_ (_10175_, _10174_, _06164_);
  and _61617_ (_10176_, _10174_, _06164_);
  nor _61618_ (_10177_, _06675_, \oc8051_golden_model_1.PC [4]);
  nor _61619_ (_10178_, _10177_, _10171_);
  not _61620_ (_10179_, _10178_);
  nor _61621_ (_10180_, _10179_, _06195_);
  nor _61622_ (_10181_, _06674_, \oc8051_golden_model_1.PC [3]);
  nor _61623_ (_10182_, _10181_, _06675_);
  not _61624_ (_10183_, _10182_);
  nor _61625_ (_10184_, _10183_, _03742_);
  and _61626_ (_10185_, _10183_, _03742_);
  nor _61627_ (_10186_, _02891_, \oc8051_golden_model_1.PC [2]);
  nor _61628_ (_10187_, _10186_, _06674_);
  not _61629_ (_10188_, _10187_);
  nor _61630_ (_10189_, _10188_, _03920_);
  not _61631_ (_10190_, _03234_);
  nor _61632_ (_10191_, _04317_, _10190_);
  nor _61633_ (_10192_, _04109_, \oc8051_golden_model_1.PC [0]);
  and _61634_ (_10193_, _04317_, _10190_);
  nor _61635_ (_10194_, _10193_, _10191_);
  and _61636_ (_10195_, _10194_, _10192_);
  nor _61637_ (_10196_, _10195_, _10191_);
  and _61638_ (_10197_, _10188_, _03920_);
  nor _61639_ (_10198_, _10197_, _10189_);
  not _61640_ (_10199_, _10198_);
  nor _61641_ (_10200_, _10199_, _10196_);
  nor _61642_ (_10201_, _10200_, _10189_);
  nor _61643_ (_10202_, _10201_, _10185_);
  nor _61644_ (_10203_, _10202_, _10184_);
  and _61645_ (_10204_, _10179_, _06195_);
  nor _61646_ (_10205_, _10204_, _10180_);
  not _61647_ (_10206_, _10205_);
  nor _61648_ (_10207_, _10206_, _10203_);
  nor _61649_ (_10208_, _10207_, _10180_);
  nor _61650_ (_10209_, _10208_, _10176_);
  nor _61651_ (_10210_, _10209_, _10175_);
  nor _61652_ (_10211_, _10210_, _10170_);
  nor _61653_ (_10212_, _10211_, _10167_);
  nor _61654_ (_10213_, _10212_, _10162_);
  or _61655_ (_10214_, _10213_, _10161_);
  nor _61656_ (_10215_, _06677_, \oc8051_golden_model_1.PC [8]);
  nor _61657_ (_10216_, _10215_, _10118_);
  not _61658_ (_10217_, _10216_);
  nor _61659_ (_10218_, _10217_, _06086_);
  and _61660_ (_10219_, _10217_, _06086_);
  nor _61661_ (_10220_, _10219_, _10218_);
  and _61662_ (_10221_, _10220_, _10214_);
  and _61663_ (_10222_, _10221_, _10160_);
  and _61664_ (_10223_, _10222_, _10154_);
  nor _61665_ (_10224_, _10218_, _10158_);
  not _61666_ (_10225_, _10224_);
  and _61667_ (_10226_, _10225_, _10154_);
  or _61668_ (_10227_, _10226_, _10149_);
  nor _61669_ (_10228_, _10227_, _10223_);
  and _61670_ (_10229_, _10228_, _10145_);
  and _61671_ (_10230_, _10139_, _06086_);
  nor _61672_ (_10231_, _10230_, _10140_);
  not _61673_ (_10232_, _10231_);
  nor _61674_ (_10233_, _10232_, _10229_);
  nor _61675_ (_10234_, _10233_, _10140_);
  nor _61676_ (_10235_, _10234_, _10136_);
  nor _61677_ (_10236_, _10235_, _10135_);
  nor _61678_ (_10237_, _10236_, _10131_);
  nor _61679_ (_10238_, _10237_, _10128_);
  not _61680_ (_10239_, _06754_);
  and _61681_ (_10240_, _10239_, _06086_);
  nor _61682_ (_10241_, _10239_, _06086_);
  nor _61683_ (_10242_, _10241_, _10240_);
  and _61684_ (_10243_, _10242_, _10238_);
  nor _61685_ (_10244_, _10242_, _10238_);
  nor _61686_ (_10245_, _10244_, _10243_);
  nor _61687_ (_10246_, _10245_, _10116_);
  or _61688_ (_10247_, _10246_, _10117_);
  and _61689_ (_10248_, _10247_, _03657_);
  not _61690_ (_10249_, _03206_);
  nor _61691_ (_10250_, _03511_, _10249_);
  and _61692_ (_10251_, _10250_, _03513_);
  or _61693_ (_10252_, _10251_, _06746_);
  and _61694_ (_10253_, _06746_, _03575_);
  nor _61695_ (_10254_, _03229_, _03202_);
  nor _61696_ (_10255_, _10254_, _07948_);
  not _61697_ (_10256_, _10255_);
  and _61698_ (_10257_, _05617_, _05940_);
  and _61699_ (_10258_, _05943_, _10257_);
  and _61700_ (_10259_, _05376_, _05281_);
  and _61701_ (_10260_, _10259_, _05939_);
  and _61702_ (_10261_, _10260_, _10258_);
  nor _61703_ (_10262_, _10261_, _10245_);
  and _61704_ (_10263_, _10261_, _06754_);
  or _61705_ (_10264_, _10263_, _04444_);
  or _61706_ (_10265_, _10264_, _10262_);
  and _61707_ (_10266_, _05824_, _05822_);
  and _61708_ (_10267_, _04603_, _04419_);
  and _61709_ (_10268_, _06699_, _10267_);
  and _61710_ (_10269_, _10268_, _10266_);
  or _61711_ (_10270_, _10269_, _10074_);
  nand _61712_ (_10271_, _10268_, _10266_);
  or _61713_ (_10272_, _10271_, _06746_);
  and _61714_ (_10273_, _10272_, _05833_);
  and _61715_ (_10274_, _10273_, _10270_);
  not _61716_ (_10275_, _04012_);
  nand _61717_ (_10276_, _06747_, _04426_);
  and _61718_ (_10277_, _10276_, _10275_);
  nor _61719_ (_10278_, _04720_, _04713_);
  nand _61720_ (_10279_, _10278_, _06736_);
  or _61721_ (_10280_, _10278_, _09946_);
  and _61722_ (_10281_, _10280_, _10279_);
  or _61723_ (_10282_, _10281_, _04426_);
  and _61724_ (_10283_, _10282_, _10277_);
  and _61725_ (_10284_, _09946_, _04012_);
  or _61726_ (_10285_, _10284_, _10283_);
  and _61727_ (_10286_, _10285_, _04762_);
  nand _61728_ (_10287_, _06746_, _03923_);
  not _61729_ (_10288_, _07933_);
  nor _61730_ (_10289_, _07935_, _07945_);
  and _61731_ (_10290_, _10289_, _10288_);
  nand _61732_ (_10291_, _10290_, _10287_);
  or _61733_ (_10292_, _10291_, _10286_);
  or _61734_ (_10293_, _10290_, _09946_);
  and _61735_ (_10294_, _10293_, _05831_);
  and _61736_ (_10295_, _10294_, _10292_);
  nor _61737_ (_10296_, _04438_, _03570_);
  not _61738_ (_10297_, _10296_);
  or _61739_ (_10298_, _10297_, _10295_);
  or _61740_ (_10299_, _10298_, _10274_);
  and _61741_ (_10300_, _10299_, _10265_);
  or _61742_ (_10301_, _10300_, _10256_);
  and _61743_ (_10302_, _03576_, _03203_);
  and _61744_ (_10303_, _10255_, _05847_);
  or _61745_ (_10304_, _10303_, _09946_);
  and _61746_ (_10305_, _10304_, _10302_);
  and _61747_ (_10306_, _10305_, _10301_);
  and _61748_ (_10307_, _07927_, _07987_);
  or _61749_ (_10308_, _10302_, _06747_);
  nand _61750_ (_10309_, _10308_, _10307_);
  or _61751_ (_10310_, _10309_, _10306_);
  or _61752_ (_10311_, _10307_, _09946_);
  and _61753_ (_10312_, _10311_, _03583_);
  and _61754_ (_10313_, _10312_, _10310_);
  or _61755_ (_10314_, _10313_, _10253_);
  nor _61756_ (_10315_, _03229_, _03205_);
  nor _61757_ (_10316_, _10315_, _07991_);
  and _61758_ (_10317_, _10316_, _10314_);
  not _61759_ (_10318_, _09946_);
  or _61760_ (_10319_, _10316_, _10318_);
  nand _61761_ (_10320_, _10319_, _10251_);
  or _61762_ (_10321_, _10320_, _10317_);
  and _61763_ (_10322_, _10321_, _10252_);
  and _61764_ (_10323_, _03476_, _03504_);
  nor _61765_ (_10324_, _07778_, _03199_);
  nor _61766_ (_10325_, _10324_, _10323_);
  not _61767_ (_10326_, _10325_);
  or _61768_ (_10327_, _10326_, _10322_);
  not _61769_ (_10328_, _03657_);
  and _61770_ (_10329_, _05176_, _03401_);
  not _61771_ (_10330_, _10329_);
  and _61772_ (_10331_, _10330_, _05177_);
  nor _61773_ (_10332_, _05327_, _04956_);
  and _61774_ (_10333_, _05327_, _04956_);
  nor _61775_ (_10334_, _10333_, _10332_);
  and _61776_ (_10335_, _10334_, _10331_);
  and _61777_ (_10336_, _05422_, _05190_);
  not _61778_ (_10337_, _10336_);
  or _61779_ (_10338_, _05422_, _05190_);
  and _61780_ (_10339_, _10338_, _10337_);
  and _61781_ (_10340_, _05712_, _05182_);
  nor _61782_ (_10341_, _05712_, _05182_);
  nor _61783_ (_10342_, _10341_, _10340_);
  and _61784_ (_10343_, _10342_, _10339_);
  and _61785_ (_10344_, _10343_, _10335_);
  and _61786_ (_10345_, _04843_, _03563_);
  and _61787_ (_10346_, _05026_, _04965_);
  nor _61788_ (_10347_, _10346_, _10345_);
  or _61789_ (_10348_, _04843_, _03563_);
  or _61790_ (_10349_, _05026_, _04965_);
  and _61791_ (_10350_, _10349_, _10348_);
  and _61792_ (_10351_, _10350_, _10347_);
  or _61793_ (_10352_, _04439_, _03472_);
  nor _61794_ (_10353_, _04603_, _04548_);
  and _61795_ (_10354_, _04603_, _04548_);
  nor _61796_ (_10355_, _10354_, _10353_);
  and _61797_ (_10356_, _10355_, _10352_);
  or _61798_ (_10357_, _04419_, _03471_);
  and _61799_ (_10358_, _10357_, _10356_);
  and _61800_ (_10359_, _10358_, _10351_);
  and _61801_ (_10360_, _10359_, _10344_);
  and _61802_ (_10361_, _10360_, _06754_);
  nor _61803_ (_10362_, _10360_, _10245_);
  or _61804_ (_10363_, _10362_, _10361_);
  or _61805_ (_10364_, _10363_, _10325_);
  and _61806_ (_10365_, _10364_, _10328_);
  and _61807_ (_10366_, _10365_, _10327_);
  or _61808_ (_10367_, _10366_, _10248_);
  and _61809_ (_10368_, _10367_, _03998_);
  nor _61810_ (_10369_, _08143_, \oc8051_golden_model_1.ACC [3]);
  and _61811_ (_10370_, _08143_, \oc8051_golden_model_1.ACC [3]);
  nor _61812_ (_10371_, _10370_, _10369_);
  and _61813_ (_10372_, _10371_, _08621_);
  nor _61814_ (_10373_, _08191_, \oc8051_golden_model_1.ACC [0]);
  and _61815_ (_10374_, _08191_, \oc8051_golden_model_1.ACC [0]);
  nor _61816_ (_10375_, _10374_, _10373_);
  and _61817_ (_10376_, _10375_, _08625_);
  and _61818_ (_10377_, _10376_, _10372_);
  and _61819_ (_10378_, _08610_, _08614_);
  not _61820_ (_10379_, _08601_);
  and _61821_ (_10380_, _08605_, _10379_);
  and _61822_ (_10381_, _10380_, _10378_);
  and _61823_ (_10382_, _10381_, _10377_);
  nor _61824_ (_10383_, _10382_, _10245_);
  and _61825_ (_10384_, _10382_, _06754_);
  or _61826_ (_10385_, _10384_, _10383_);
  and _61827_ (_10386_, _10385_, _03527_);
  or _61828_ (_10387_, _10386_, _10368_);
  and _61829_ (_10388_, _10387_, _10085_);
  nor _61830_ (_10389_, _08652_, _08656_);
  nor _61831_ (_10390_, _08649_, _08422_);
  and _61832_ (_10391_, _10390_, _10389_);
  nor _61833_ (_10392_, _08657_, _08658_);
  nor _61834_ (_10393_, _10392_, _08661_);
  and _61835_ (_10394_, _03471_, _03321_);
  nor _61836_ (_10395_, _10394_, _08666_);
  nor _61837_ (_10396_, _10395_, _08665_);
  and _61838_ (_10397_, _10396_, _10393_);
  and _61839_ (_10398_, _10397_, _10391_);
  not _61840_ (_10399_, _10398_);
  nand _61841_ (_10400_, _10399_, _10245_);
  nand _61842_ (_10401_, _10398_, _10239_);
  and _61843_ (_10402_, _10401_, _03638_);
  and _61844_ (_10403_, _10402_, _10400_);
  or _61845_ (_10404_, _10403_, _10388_);
  and _61846_ (_10405_, _10404_, _10084_);
  nand _61847_ (_10406_, _10083_, _09946_);
  and _61848_ (_10407_, _04897_, _03593_);
  and _61849_ (_10408_, _10407_, _03602_);
  nand _61850_ (_10409_, _10408_, _10406_);
  or _61851_ (_10410_, _10409_, _10405_);
  or _61852_ (_10411_, _10408_, _06746_);
  and _61853_ (_10412_, _03220_, _03596_);
  not _61854_ (_10413_, _10412_);
  nor _61855_ (_10414_, _09770_, _06794_);
  and _61856_ (_10415_, _10414_, _10413_);
  and _61857_ (_10416_, _10415_, _10411_);
  and _61858_ (_10417_, _10416_, _10410_);
  nor _61859_ (_10418_, _10415_, _10318_);
  not _61860_ (_10419_, _03607_);
  not _61861_ (_10420_, _03213_);
  nor _61862_ (_10421_, _03606_, _10420_);
  and _61863_ (_10422_, _10421_, _10419_);
  not _61864_ (_10423_, _10422_);
  or _61865_ (_10424_, _10423_, _10418_);
  or _61866_ (_10425_, _10424_, _10417_);
  nor _61867_ (_10426_, _08035_, _07923_);
  or _61868_ (_10427_, _10422_, _06746_);
  and _61869_ (_10428_, _10427_, _10426_);
  and _61870_ (_10429_, _10428_, _10425_);
  nor _61871_ (_10430_, _08108_, _03614_);
  not _61872_ (_10431_, _10430_);
  nor _61873_ (_10432_, _10426_, _10318_);
  or _61874_ (_10433_, _10432_, _10431_);
  or _61875_ (_10434_, _10433_, _10429_);
  or _61876_ (_10435_, _10430_, _06746_);
  and _61877_ (_10436_, _10435_, _03254_);
  and _61878_ (_10437_, _10436_, _10434_);
  or _61879_ (_10438_, _10318_, _03254_);
  nor _61880_ (_10439_, _03499_, _03223_);
  nand _61881_ (_10440_, _10439_, _10438_);
  or _61882_ (_10441_, _10440_, _10437_);
  or _61883_ (_10442_, _10439_, _06746_);
  and _61884_ (_10443_, _10442_, _09755_);
  and _61885_ (_10444_, _10443_, _10441_);
  nand _61886_ (_10445_, _06754_, _03632_);
  nand _61887_ (_10446_, _10445_, _03493_);
  or _61888_ (_10447_, _10446_, _10444_);
  or _61889_ (_10448_, _06746_, _03493_);
  and _61890_ (_10449_, _10448_, _03474_);
  and _61891_ (_10450_, _10449_, _10447_);
  or _61892_ (_10451_, _10450_, _10082_);
  and _61893_ (_10452_, _10451_, _10081_);
  nor _61894_ (_10453_, _03745_, _03187_);
  not _61895_ (_10454_, _10453_);
  nor _61896_ (_10455_, _10081_, _10318_);
  or _61897_ (_10456_, _10455_, _10454_);
  or _61898_ (_10457_, _10456_, _10452_);
  and _61899_ (_10458_, _03186_, _03150_);
  not _61900_ (_10459_, _10458_);
  or _61901_ (_10460_, _10453_, _06746_);
  and _61902_ (_10461_, _10460_, _10459_);
  and _61903_ (_10462_, _10461_, _10457_);
  and _61904_ (_10463_, _10458_, _10074_);
  or _61905_ (_10464_, _10463_, _06055_);
  or _61906_ (_10465_, _10464_, _10462_);
  or _61907_ (_10466_, _06746_, _05775_);
  and _61908_ (_10467_, _10466_, _03438_);
  and _61909_ (_10468_, _10467_, _10465_);
  and _61910_ (_10469_, _06754_, _03437_);
  or _61911_ (_10470_, _10469_, _08385_);
  or _61912_ (_10471_, _10470_, _10468_);
  and _61913_ (_10472_, _03230_, _03188_);
  and _61914_ (_10473_, _08385_, _06747_);
  nor _61915_ (_10474_, _10473_, _10472_);
  and _61916_ (_10475_, _10474_, _10471_);
  not _61917_ (_10476_, \oc8051_golden_model_1.DPH [0]);
  and _61918_ (_10477_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor _61919_ (_10478_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and _61920_ (_10479_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _61921_ (_10480_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _61922_ (_10481_, _10480_, _10479_);
  and _61923_ (_10482_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _61924_ (_10483_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _61925_ (_10484_, _10483_, _10482_);
  not _61926_ (_10485_, _10484_);
  and _61927_ (_10486_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _61928_ (_10487_, _03287_, _03283_);
  not _61929_ (_10488_, _10487_);
  nor _61930_ (_10489_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _61931_ (_10490_, _10489_, _10486_);
  and _61932_ (_10491_, _10490_, _10488_);
  nor _61933_ (_10492_, _10491_, _10486_);
  nor _61934_ (_10493_, _10492_, _10485_);
  nor _61935_ (_10494_, _10493_, _10482_);
  not _61936_ (_10495_, _10494_);
  and _61937_ (_10496_, _10495_, _10481_);
  nor _61938_ (_10497_, _10496_, _10479_);
  nor _61939_ (_10498_, _10497_, _10478_);
  nor _61940_ (_10499_, _10498_, _10477_);
  nor _61941_ (_10500_, _10499_, _10476_);
  and _61942_ (_10501_, _10500_, \oc8051_golden_model_1.DPH [1]);
  and _61943_ (_10502_, _10501_, \oc8051_golden_model_1.DPH [2]);
  and _61944_ (_10503_, _10502_, \oc8051_golden_model_1.DPH [3]);
  and _61945_ (_10504_, _10503_, \oc8051_golden_model_1.DPH [4]);
  and _61946_ (_10505_, _10504_, \oc8051_golden_model_1.DPH [5]);
  and _61947_ (_10506_, _10505_, \oc8051_golden_model_1.DPH [6]);
  nand _61948_ (_10507_, _10506_, \oc8051_golden_model_1.DPH [7]);
  or _61949_ (_10508_, _10506_, \oc8051_golden_model_1.DPH [7]);
  and _61950_ (_10509_, _10508_, _10472_);
  and _61951_ (_10510_, _10509_, _10507_);
  nor _61952_ (_10511_, _03744_, _03189_);
  not _61953_ (_10512_, _10511_);
  or _61954_ (_10513_, _10512_, _10510_);
  or _61955_ (_10514_, _10513_, _10475_);
  not _61956_ (_10515_, _10076_);
  or _61957_ (_10516_, _10511_, _06746_);
  and _61958_ (_10517_, _10516_, _10515_);
  and _61959_ (_10518_, _10517_, _10514_);
  or _61960_ (_10519_, _10518_, _10080_);
  and _61961_ (_10520_, _08409_, _08397_);
  and _61962_ (_10521_, _10520_, _10519_);
  nor _61963_ (_10522_, _10520_, _10318_);
  nor _61964_ (_10523_, _08415_, _03767_);
  not _61965_ (_10524_, _10523_);
  or _61966_ (_10525_, _10524_, _10522_);
  or _61967_ (_10526_, _10525_, _10521_);
  or _61968_ (_10527_, _10523_, _06746_);
  and _61969_ (_10528_, _10527_, _04499_);
  and _61970_ (_10529_, _10528_, _10526_);
  nand _61971_ (_10530_, _06754_, _03636_);
  nor _61972_ (_10531_, _03769_, _03194_);
  nand _61973_ (_10532_, _10531_, _10530_);
  or _61974_ (_10533_, _10532_, _10529_);
  and _61975_ (_10534_, _03193_, _03150_);
  not _61976_ (_10535_, _10534_);
  or _61977_ (_10536_, _10531_, _06746_);
  and _61978_ (_10537_, _10536_, _10535_);
  and _61979_ (_10538_, _10537_, _10533_);
  or _61980_ (_10539_, _10074_, _10077_);
  or _61981_ (_10540_, _08698_, _06746_);
  and _61982_ (_10541_, _10540_, _10534_);
  and _61983_ (_10542_, _10541_, _10539_);
  or _61984_ (_10543_, _10542_, _10538_);
  not _61985_ (_10544_, _03191_);
  nor _61986_ (_10545_, _09948_, _10544_);
  not _61987_ (_10546_, _10545_);
  and _61988_ (_10547_, _10546_, _10543_);
  nor _61989_ (_10548_, _07909_, _03755_);
  not _61990_ (_10549_, _10548_);
  and _61991_ (_10550_, _10545_, _09946_);
  or _61992_ (_10551_, _10550_, _10549_);
  or _61993_ (_10552_, _10551_, _10547_);
  or _61994_ (_10553_, _10548_, _06746_);
  and _61995_ (_10554_, _10553_, _05769_);
  and _61996_ (_10555_, _10554_, _10552_);
  nand _61997_ (_10556_, _06754_, _03754_);
  nand _61998_ (_10557_, _10556_, _09960_);
  or _61999_ (_10558_, _10557_, _10555_);
  and _62000_ (_10559_, _10558_, _09962_);
  not _62001_ (_10560_, _09956_);
  or _62002_ (_10561_, _10074_, \oc8051_golden_model_1.PSW [7]);
  or _62003_ (_10562_, _06746_, _07888_);
  and _62004_ (_10563_, _10562_, _09958_);
  and _62005_ (_10564_, _10563_, _10561_);
  or _62006_ (_10565_, _10564_, _10560_);
  or _62007_ (_10566_, _10565_, _10559_);
  and _62008_ (_10567_, _10566_, _09957_);
  or _62009_ (_10568_, _10567_, _08479_);
  or _62010_ (_10569_, _08478_, _06746_);
  and _62011_ (_10570_, _10569_, _03759_);
  and _62012_ (_10571_, _10570_, _10568_);
  nand _62013_ (_10572_, _06754_, _03758_);
  nor _62014_ (_10573_, _03760_, _03183_);
  nand _62015_ (_10574_, _10573_, _10572_);
  or _62016_ (_10575_, _10574_, _10571_);
  and _62017_ (_10576_, _03182_, _03150_);
  not _62018_ (_10577_, _10576_);
  or _62019_ (_10578_, _10573_, _06746_);
  and _62020_ (_10579_, _10578_, _10577_);
  and _62021_ (_10580_, _10579_, _10575_);
  not _62022_ (_10581_, _09951_);
  or _62023_ (_10582_, _10074_, _07888_);
  or _62024_ (_10583_, _06746_, \oc8051_golden_model_1.PSW [7]);
  and _62025_ (_10584_, _10583_, _10576_);
  and _62026_ (_10585_, _10584_, _10582_);
  or _62027_ (_10586_, _10585_, _10581_);
  or _62028_ (_10587_, _10586_, _10580_);
  and _62029_ (_10588_, _10587_, _09952_);
  or _62030_ (_10589_, _10588_, _08525_);
  or _62031_ (_10590_, _08524_, _06746_);
  and _62032_ (_10591_, _10590_, _08556_);
  and _62033_ (_10592_, _10591_, _10589_);
  and _62034_ (_10593_, _09946_, _08555_);
  or _62035_ (_10594_, _10593_, _03775_);
  or _62036_ (_10595_, _10594_, _10592_);
  nand _62037_ (_10596_, _05176_, _03775_);
  and _62038_ (_10597_, _10596_, _10595_);
  or _62039_ (_10598_, _10597_, _03179_);
  not _62040_ (_10599_, _03627_);
  nand _62041_ (_10600_, _06747_, _03179_);
  and _62042_ (_10601_, _10600_, _10599_);
  and _62043_ (_10602_, _10601_, _10598_);
  not _62044_ (_10603_, _09949_);
  not _62045_ (_10604_, _05271_);
  and _62046_ (_10605_, _05799_, \oc8051_golden_model_1.TCON [2]);
  and _62047_ (_10606_, _05785_, \oc8051_golden_model_1.B [2]);
  nor _62048_ (_10607_, _10606_, _10605_);
  and _62049_ (_10608_, _05790_, \oc8051_golden_model_1.IP [2]);
  not _62050_ (_10609_, _10608_);
  and _62051_ (_10610_, _05783_, \oc8051_golden_model_1.PSW [2]);
  and _62052_ (_10611_, _05792_, \oc8051_golden_model_1.ACC [2]);
  nor _62053_ (_10612_, _10611_, _10610_);
  and _62054_ (_10613_, _10612_, _10609_);
  and _62055_ (_10614_, _10613_, _10607_);
  and _62056_ (_10615_, _05805_, \oc8051_golden_model_1.SCON [2]);
  and _62057_ (_10616_, _05807_, \oc8051_golden_model_1.IE [2]);
  nor _62058_ (_10617_, _10616_, _10615_);
  and _62059_ (_10618_, _05811_, \oc8051_golden_model_1.P1INREG [2]);
  and _62060_ (_10619_, _05796_, \oc8051_golden_model_1.P3INREG [2]);
  nor _62061_ (_10620_, _10619_, _10618_);
  and _62062_ (_10621_, _05205_, \oc8051_golden_model_1.P0INREG [2]);
  and _62063_ (_10622_, _05801_, \oc8051_golden_model_1.P2INREG [2]);
  nor _62064_ (_10623_, _10622_, _10621_);
  and _62065_ (_10624_, _10623_, _10620_);
  and _62066_ (_10625_, _10624_, _10617_);
  and _62067_ (_10626_, _10625_, _10614_);
  and _62068_ (_10627_, _10626_, _05619_);
  nor _62069_ (_10628_, _10627_, _10604_);
  not _62070_ (_10629_, _05179_);
  and _62071_ (_10630_, _05805_, \oc8051_golden_model_1.SCON [1]);
  and _62072_ (_10631_, _05807_, \oc8051_golden_model_1.IE [1]);
  nor _62073_ (_10632_, _10631_, _10630_);
  and _62074_ (_10633_, _05799_, \oc8051_golden_model_1.TCON [1]);
  and _62075_ (_10634_, _05796_, \oc8051_golden_model_1.P3INREG [1]);
  nor _62076_ (_10635_, _10634_, _10633_);
  and _62077_ (_10636_, _10635_, _10632_);
  and _62078_ (_10637_, _05790_, \oc8051_golden_model_1.IP [1]);
  and _62079_ (_10638_, _05785_, \oc8051_golden_model_1.B [1]);
  nor _62080_ (_10639_, _10638_, _10637_);
  and _62081_ (_10640_, _05783_, \oc8051_golden_model_1.PSW [1]);
  and _62082_ (_10641_, _05792_, \oc8051_golden_model_1.ACC [1]);
  nor _62083_ (_10642_, _10641_, _10640_);
  and _62084_ (_10643_, _10642_, _10639_);
  and _62085_ (_10644_, _05811_, \oc8051_golden_model_1.P1INREG [1]);
  and _62086_ (_10645_, _05801_, \oc8051_golden_model_1.P2INREG [1]);
  and _62087_ (_10646_, _05205_, \oc8051_golden_model_1.P0INREG [1]);
  or _62088_ (_10647_, _10646_, _10645_);
  nor _62089_ (_10648_, _10647_, _10644_);
  and _62090_ (_10649_, _10648_, _10643_);
  and _62091_ (_10650_, _10649_, _10636_);
  and _62092_ (_10651_, _10650_, _05522_);
  nor _62093_ (_10652_, _10651_, _10629_);
  nor _62094_ (_10653_, _10652_, _10628_);
  and _62095_ (_10654_, _05187_, _04965_);
  not _62096_ (_10655_, _10654_);
  and _62097_ (_10656_, _05805_, \oc8051_golden_model_1.SCON [4]);
  and _62098_ (_10657_, _05807_, \oc8051_golden_model_1.IE [4]);
  nor _62099_ (_10658_, _10657_, _10656_);
  and _62100_ (_10659_, _05799_, \oc8051_golden_model_1.TCON [4]);
  and _62101_ (_10660_, _05796_, \oc8051_golden_model_1.P3INREG [4]);
  nor _62102_ (_10661_, _10660_, _10659_);
  and _62103_ (_10662_, _10661_, _10658_);
  and _62104_ (_10663_, _05783_, \oc8051_golden_model_1.PSW [4]);
  and _62105_ (_10664_, _05792_, \oc8051_golden_model_1.ACC [4]);
  nor _62106_ (_10665_, _10664_, _10663_);
  and _62107_ (_10666_, _05790_, \oc8051_golden_model_1.IP [4]);
  and _62108_ (_10667_, _05785_, \oc8051_golden_model_1.B [4]);
  nor _62109_ (_10668_, _10667_, _10666_);
  and _62110_ (_10669_, _10668_, _10665_);
  and _62111_ (_10670_, _05811_, \oc8051_golden_model_1.P1INREG [4]);
  and _62112_ (_10671_, _05801_, \oc8051_golden_model_1.P2INREG [4]);
  and _62113_ (_10672_, _05205_, \oc8051_golden_model_1.P0INREG [4]);
  or _62114_ (_10673_, _10672_, _10671_);
  nor _62115_ (_10674_, _10673_, _10670_);
  and _62116_ (_10675_, _10674_, _10669_);
  and _62117_ (_10676_, _10675_, _10662_);
  and _62118_ (_10677_, _10676_, _05713_);
  nor _62119_ (_10678_, _10677_, _10655_);
  nor _62120_ (_10679_, _06029_, _05953_);
  nor _62121_ (_10680_, _10679_, _10678_);
  and _62122_ (_10681_, _10680_, _10653_);
  not _62123_ (_10682_, _05188_);
  and _62124_ (_10683_, _05799_, \oc8051_golden_model_1.TCON [0]);
  and _62125_ (_10684_, _05785_, \oc8051_golden_model_1.B [0]);
  nor _62126_ (_10685_, _10684_, _10683_);
  and _62127_ (_10686_, _05783_, \oc8051_golden_model_1.PSW [0]);
  not _62128_ (_10687_, _10686_);
  and _62129_ (_10688_, _05790_, \oc8051_golden_model_1.IP [0]);
  and _62130_ (_10689_, _05792_, \oc8051_golden_model_1.ACC [0]);
  nor _62131_ (_10691_, _10689_, _10688_);
  and _62132_ (_10692_, _10691_, _10687_);
  and _62133_ (_10693_, _10692_, _10685_);
  and _62134_ (_10694_, _05805_, \oc8051_golden_model_1.SCON [0]);
  and _62135_ (_10695_, _05807_, \oc8051_golden_model_1.IE [0]);
  nor _62136_ (_10696_, _10695_, _10694_);
  and _62137_ (_10697_, _05205_, \oc8051_golden_model_1.P0INREG [0]);
  and _62138_ (_10698_, _05801_, \oc8051_golden_model_1.P2INREG [0]);
  nor _62139_ (_10699_, _10698_, _10697_);
  and _62140_ (_10700_, _05811_, \oc8051_golden_model_1.P1INREG [0]);
  and _62141_ (_10702_, _05796_, \oc8051_golden_model_1.P3INREG [0]);
  nor _62142_ (_10703_, _10702_, _10700_);
  and _62143_ (_10704_, _10703_, _10699_);
  and _62144_ (_10705_, _10704_, _10696_);
  and _62145_ (_10706_, _10705_, _10693_);
  and _62146_ (_10707_, _10706_, _05570_);
  nor _62147_ (_10708_, _10707_, _10682_);
  and _62148_ (_10709_, _05256_, _04965_);
  not _62149_ (_10710_, _10709_);
  and _62150_ (_10711_, _05799_, \oc8051_golden_model_1.TCON [6]);
  and _62151_ (_10713_, _05785_, \oc8051_golden_model_1.B [6]);
  nor _62152_ (_10714_, _10713_, _10711_);
  and _62153_ (_10715_, _05790_, \oc8051_golden_model_1.IP [6]);
  not _62154_ (_10716_, _10715_);
  and _62155_ (_10717_, _05783_, \oc8051_golden_model_1.PSW [6]);
  and _62156_ (_10718_, _05792_, \oc8051_golden_model_1.ACC [6]);
  nor _62157_ (_10719_, _10718_, _10717_);
  and _62158_ (_10720_, _10719_, _10716_);
  and _62159_ (_10721_, _10720_, _10714_);
  and _62160_ (_10722_, _05805_, \oc8051_golden_model_1.SCON [6]);
  and _62161_ (_10724_, _05807_, \oc8051_golden_model_1.IE [6]);
  nor _62162_ (_10725_, _10724_, _10722_);
  and _62163_ (_10726_, _05205_, \oc8051_golden_model_1.P0INREG [6]);
  and _62164_ (_10727_, _05801_, \oc8051_golden_model_1.P2INREG [6]);
  nor _62165_ (_10728_, _10727_, _10726_);
  and _62166_ (_10729_, _05811_, \oc8051_golden_model_1.P1INREG [6]);
  and _62167_ (_10730_, _05796_, \oc8051_golden_model_1.P3INREG [6]);
  nor _62168_ (_10731_, _10730_, _10729_);
  and _62169_ (_10732_, _10731_, _10728_);
  and _62170_ (_10733_, _10732_, _10725_);
  and _62171_ (_10735_, _10733_, _10721_);
  and _62172_ (_10736_, _10735_, _05328_);
  nor _62173_ (_10737_, _10736_, _10710_);
  nor _62174_ (_10738_, _10737_, _10708_);
  not _62175_ (_10739_, _05265_);
  and _62176_ (_10740_, _05783_, \oc8051_golden_model_1.PSW [3]);
  and _62177_ (_10741_, _05792_, \oc8051_golden_model_1.ACC [3]);
  nor _62178_ (_10742_, _10741_, _10740_);
  and _62179_ (_10743_, _05790_, \oc8051_golden_model_1.IP [3]);
  and _62180_ (_10744_, _05785_, \oc8051_golden_model_1.B [3]);
  nor _62181_ (_10746_, _10744_, _10743_);
  and _62182_ (_10747_, _10746_, _10742_);
  and _62183_ (_10748_, _05801_, \oc8051_golden_model_1.P2INREG [3]);
  not _62184_ (_10749_, _10748_);
  and _62185_ (_10750_, _05205_, \oc8051_golden_model_1.P0INREG [3]);
  and _62186_ (_10751_, _05796_, \oc8051_golden_model_1.P3INREG [3]);
  nor _62187_ (_10752_, _10751_, _10750_);
  and _62188_ (_10753_, _10752_, _10749_);
  and _62189_ (_10754_, _05805_, \oc8051_golden_model_1.SCON [3]);
  and _62190_ (_10755_, _05807_, \oc8051_golden_model_1.IE [3]);
  nor _62191_ (_10757_, _10755_, _10754_);
  and _62192_ (_10758_, _05799_, \oc8051_golden_model_1.TCON [3]);
  and _62193_ (_10759_, _05811_, \oc8051_golden_model_1.P1INREG [3]);
  nor _62194_ (_10760_, _10759_, _10758_);
  and _62195_ (_10761_, _10760_, _10757_);
  and _62196_ (_10762_, _10761_, _10753_);
  and _62197_ (_10763_, _10762_, _10747_);
  and _62198_ (_10764_, _10763_, _05473_);
  nor _62199_ (_10765_, _10764_, _10739_);
  and _62200_ (_10766_, _05178_, _04965_);
  not _62201_ (_10767_, _10766_);
  and _62202_ (_10768_, _05799_, \oc8051_golden_model_1.TCON [5]);
  and _62203_ (_10769_, _05785_, \oc8051_golden_model_1.B [5]);
  nor _62204_ (_10770_, _10769_, _10768_);
  and _62205_ (_10771_, _05783_, \oc8051_golden_model_1.PSW [5]);
  not _62206_ (_10772_, _10771_);
  and _62207_ (_10773_, _05790_, \oc8051_golden_model_1.IP [5]);
  and _62208_ (_10774_, _05792_, \oc8051_golden_model_1.ACC [5]);
  nor _62209_ (_10775_, _10774_, _10773_);
  and _62210_ (_10776_, _10775_, _10772_);
  and _62211_ (_10777_, _10776_, _10770_);
  and _62212_ (_10778_, _05805_, \oc8051_golden_model_1.SCON [5]);
  and _62213_ (_10779_, _05807_, \oc8051_golden_model_1.IE [5]);
  nor _62214_ (_10780_, _10779_, _10778_);
  and _62215_ (_10781_, _05205_, \oc8051_golden_model_1.P0INREG [5]);
  and _62216_ (_10782_, _05801_, \oc8051_golden_model_1.P2INREG [5]);
  nor _62217_ (_10783_, _10782_, _10781_);
  and _62218_ (_10784_, _05811_, \oc8051_golden_model_1.P1INREG [5]);
  and _62219_ (_10785_, _05796_, \oc8051_golden_model_1.P3INREG [5]);
  nor _62220_ (_10786_, _10785_, _10784_);
  and _62221_ (_10787_, _10786_, _10783_);
  and _62222_ (_10788_, _10787_, _10780_);
  and _62223_ (_10789_, _10788_, _10777_);
  and _62224_ (_10790_, _10789_, _05423_);
  nor _62225_ (_10791_, _10790_, _10767_);
  nor _62226_ (_10792_, _10791_, _10765_);
  and _62227_ (_10793_, _10792_, _10738_);
  and _62228_ (_10794_, _10793_, _10681_);
  nand _62229_ (_10795_, _10794_, _10245_);
  or _62230_ (_10796_, _10794_, _06754_);
  and _62231_ (_10797_, _10796_, _03627_);
  and _62232_ (_10798_, _10797_, _10795_);
  or _62233_ (_10799_, _10798_, _10603_);
  or _62234_ (_10800_, _10799_, _10602_);
  and _62235_ (_10801_, _10800_, _09950_);
  or _62236_ (_10802_, _10801_, _09937_);
  not _62237_ (_10803_, _07729_);
  or _62238_ (_10804_, _09936_, _06746_);
  and _62239_ (_10805_, _10804_, _10803_);
  and _62240_ (_10806_, _10805_, _10802_);
  and _62241_ (_10807_, _09946_, _07729_);
  or _62242_ (_10808_, _10807_, _03522_);
  or _62243_ (_10809_, _10808_, _10806_);
  nand _62244_ (_10810_, _05176_, _03522_);
  and _62245_ (_10811_, _10810_, _10809_);
  or _62246_ (_10812_, _10811_, _03172_);
  nand _62247_ (_10813_, _06747_, _03172_);
  and _62248_ (_10814_, _10813_, _03791_);
  and _62249_ (_10815_, _10814_, _10812_);
  and _62250_ (_10816_, _10794_, _06754_);
  nor _62251_ (_10817_, _10794_, _10245_);
  or _62252_ (_10818_, _10817_, _10816_);
  and _62253_ (_10819_, _10818_, _03628_);
  and _62254_ (_10820_, _03147_, _03010_);
  nor _62255_ (_10821_, _10820_, _04527_);
  not _62256_ (_10822_, _10821_);
  or _62257_ (_10823_, _10822_, _10819_);
  or _62258_ (_10824_, _10823_, _10815_);
  or _62259_ (_10825_, _10821_, _09946_);
  and _62260_ (_10826_, _10825_, _04192_);
  and _62261_ (_10827_, _10826_, _10824_);
  nor _62262_ (_10828_, _08692_, _08687_);
  nand _62263_ (_10829_, _06746_, _03790_);
  nand _62264_ (_10830_, _10829_, _10828_);
  or _62265_ (_10831_, _10830_, _10827_);
  not _62266_ (_10832_, _03641_);
  or _62267_ (_10833_, _09946_, _10828_);
  and _62268_ (_10834_, _10833_, _10832_);
  and _62269_ (_10835_, _10834_, _10831_);
  and _62270_ (_10836_, _03641_, _03401_);
  or _62271_ (_10837_, _10836_, _03160_);
  or _62272_ (_10838_, _10837_, _10835_);
  nand _62273_ (_10839_, _06747_, _03160_);
  and _62274_ (_10840_, _10839_, _03152_);
  and _62275_ (_10841_, _10840_, _10838_);
  and _62276_ (_10842_, _10818_, _03151_);
  nor _62277_ (_10843_, _04967_, _04766_);
  and _62278_ (_10844_, _10843_, _06712_);
  not _62279_ (_10845_, _10844_);
  or _62280_ (_10846_, _10845_, _10842_);
  or _62281_ (_10847_, _10846_, _10841_);
  or _62282_ (_10848_, _10844_, _09946_);
  and _62283_ (_10849_, _10848_, _03521_);
  and _62284_ (_10850_, _10849_, _10847_);
  nor _62285_ (_10851_, _08716_, _08709_);
  nand _62286_ (_10852_, _06746_, _03520_);
  nand _62287_ (_10853_, _10852_, _10851_);
  or _62288_ (_10854_, _10853_, _10850_);
  not _62289_ (_10855_, _03645_);
  or _62290_ (_10856_, _09946_, _10851_);
  and _62291_ (_10857_, _10856_, _10855_);
  and _62292_ (_10858_, _10857_, _10854_);
  and _62293_ (_10859_, _03645_, _03401_);
  or _62294_ (_10860_, _10859_, _03166_);
  or _62295_ (_10861_, _10860_, _10858_);
  and _62296_ (_10862_, _03165_, _03150_);
  not _62297_ (_10863_, _10862_);
  nand _62298_ (_10864_, _06747_, _03166_);
  and _62299_ (_10865_, _10864_, _10863_);
  and _62300_ (_10866_, _10865_, _10861_);
  and _62301_ (_10867_, _10862_, _09946_);
  or _62302_ (_10868_, _10867_, _10866_);
  or _62303_ (_10869_, _10868_, _42967_);
  or _62304_ (_10870_, _42963_, \oc8051_golden_model_1.PC [15]);
  and _62305_ (_10871_, _10870_, _41755_);
  and _62306_ (_40533_, _10871_, _10869_);
  not _62307_ (_10872_, _05210_);
  and _62308_ (_10873_, _10872_, \oc8051_golden_model_1.P2 [7]);
  and _62309_ (_10874_, _06311_, _05210_);
  or _62310_ (_10875_, _10874_, _10873_);
  and _62311_ (_10876_, _10875_, _03769_);
  nor _62312_ (_10877_, _10872_, _05176_);
  or _62313_ (_10878_, _10877_, _10873_);
  or _62314_ (_10879_, _10878_, _06039_);
  not _62315_ (_10880_, _05801_);
  and _62316_ (_10881_, _10880_, \oc8051_golden_model_1.P2 [7]);
  and _62317_ (_10882_, _05818_, _05801_);
  or _62318_ (_10883_, _10882_, _10881_);
  and _62319_ (_10884_, _10883_, _03512_);
  and _62320_ (_10885_, _05949_, _05210_);
  or _62321_ (_10886_, _10885_, _10873_);
  or _62322_ (_10887_, _10886_, _04444_);
  and _62323_ (_10888_, _05210_, \oc8051_golden_model_1.ACC [7]);
  or _62324_ (_10889_, _10888_, _10873_);
  and _62325_ (_10890_, _10889_, _04426_);
  and _62326_ (_10891_, _04427_, \oc8051_golden_model_1.P2 [7]);
  or _62327_ (_10892_, _10891_, _03570_);
  or _62328_ (_10893_, _10892_, _10890_);
  and _62329_ (_10894_, _10893_, _03517_);
  and _62330_ (_10895_, _10894_, _10887_);
  and _62331_ (_10896_, _05954_, _05801_);
  or _62332_ (_10897_, _10896_, _10881_);
  and _62333_ (_10898_, _10897_, _03516_);
  or _62334_ (_10899_, _10898_, _03568_);
  or _62335_ (_10900_, _10899_, _10895_);
  or _62336_ (_10901_, _10878_, _03983_);
  and _62337_ (_10902_, _10901_, _10900_);
  or _62338_ (_10903_, _10902_, _03575_);
  or _62339_ (_10904_, _10889_, _03583_);
  and _62340_ (_10905_, _10904_, _03513_);
  and _62341_ (_10906_, _10905_, _10903_);
  or _62342_ (_10907_, _10906_, _10884_);
  and _62343_ (_10908_, _10907_, _03506_);
  and _62344_ (_10909_, _05990_, _05801_);
  or _62345_ (_10910_, _10909_, _10881_);
  and _62346_ (_10911_, _10910_, _03505_);
  or _62347_ (_10912_, _10911_, _10908_);
  and _62348_ (_10913_, _10912_, _03500_);
  or _62349_ (_10914_, _06032_, _05818_);
  and _62350_ (_10915_, _10914_, _05801_);
  or _62351_ (_10916_, _10915_, _10881_);
  and _62352_ (_10917_, _10916_, _03499_);
  or _62353_ (_10918_, _10917_, _07314_);
  or _62354_ (_10919_, _10918_, _10913_);
  and _62355_ (_10920_, _10919_, _10879_);
  or _62356_ (_10921_, _10920_, _03479_);
  and _62357_ (_10922_, _05935_, _05210_);
  or _62358_ (_10923_, _10873_, _06044_);
  or _62359_ (_10924_, _10923_, _10922_);
  and _62360_ (_10925_, _10924_, _03474_);
  and _62361_ (_10926_, _10925_, _10921_);
  and _62362_ (_10927_, _06214_, \oc8051_golden_model_1.P2 [7]);
  and _62363_ (_10928_, _06242_, \oc8051_golden_model_1.P0 [7]);
  or _62364_ (_10929_, _10928_, _06221_);
  or _62365_ (_10930_, _10929_, _10927_);
  and _62366_ (_10931_, _06245_, \oc8051_golden_model_1.P1 [7]);
  and _62367_ (_10932_, _06249_, \oc8051_golden_model_1.P3 [7]);
  or _62368_ (_10933_, _10932_, _10931_);
  nor _62369_ (_10934_, _10933_, _06226_);
  nand _62370_ (_10935_, _10934_, _06241_);
  nor _62371_ (_10936_, _10935_, _10930_);
  and _62372_ (_10937_, _10936_, _06208_);
  nand _62373_ (_10938_, _10937_, _06289_);
  or _62374_ (_10939_, _10938_, _06088_);
  and _62375_ (_10940_, _10939_, _05210_);
  or _62376_ (_10941_, _10940_, _10873_);
  and _62377_ (_10942_, _10941_, _03221_);
  or _62378_ (_10943_, _10942_, _03437_);
  or _62379_ (_10944_, _10943_, _10926_);
  and _62380_ (_10945_, _06087_, _05210_);
  or _62381_ (_10946_, _10945_, _10873_);
  or _62382_ (_10947_, _10946_, _03438_);
  and _62383_ (_10948_, _10947_, _10944_);
  or _62384_ (_10949_, _10948_, _03636_);
  and _62385_ (_10950_, _06305_, _05210_);
  or _62386_ (_10951_, _10950_, _10873_);
  or _62387_ (_10952_, _10951_, _04499_);
  and _62388_ (_10953_, _10952_, _04501_);
  and _62389_ (_10954_, _10953_, _10949_);
  or _62390_ (_10955_, _10954_, _10876_);
  and _62391_ (_10956_, _10955_, _05769_);
  or _62392_ (_10957_, _10873_, _05282_);
  and _62393_ (_10958_, _10957_, _03754_);
  and _62394_ (_10959_, _10958_, _10946_);
  or _62395_ (_10960_, _10959_, _10956_);
  and _62396_ (_10961_, _10960_, _03753_);
  and _62397_ (_10962_, _10889_, _03752_);
  and _62398_ (_10963_, _10962_, _10957_);
  or _62399_ (_10964_, _10963_, _03758_);
  or _62400_ (_10965_, _10964_, _10961_);
  nor _62401_ (_10966_, _06304_, _10872_);
  or _62402_ (_10967_, _10873_, _03759_);
  or _62403_ (_10968_, _10967_, _10966_);
  and _62404_ (_10969_, _10968_, _04517_);
  and _62405_ (_10970_, _10969_, _10965_);
  nor _62406_ (_10971_, _06310_, _10872_);
  or _62407_ (_10972_, _10971_, _10873_);
  and _62408_ (_10973_, _10972_, _03760_);
  or _62409_ (_10974_, _10973_, _03790_);
  or _62410_ (_10975_, _10974_, _10970_);
  or _62411_ (_10976_, _10886_, _04192_);
  and _62412_ (_10977_, _10976_, _03152_);
  and _62413_ (_10978_, _10977_, _10975_);
  and _62414_ (_10979_, _10883_, _03151_);
  or _62415_ (_10980_, _10979_, _03520_);
  or _62416_ (_10981_, _10980_, _10978_);
  and _62417_ (_10982_, _05767_, _05210_);
  or _62418_ (_10983_, _10873_, _03521_);
  or _62419_ (_10984_, _10983_, _10982_);
  and _62420_ (_10985_, _10984_, _42963_);
  and _62421_ (_10986_, _10985_, _10981_);
  nor _62422_ (_10987_, \oc8051_golden_model_1.P2 [7], rst);
  nor _62423_ (_10988_, _10987_, _00000_);
  or _62424_ (_40534_, _10988_, _10986_);
  not _62425_ (_10989_, _05200_);
  and _62426_ (_10990_, _10989_, \oc8051_golden_model_1.P3 [7]);
  and _62427_ (_10991_, _06311_, _05200_);
  or _62428_ (_10992_, _10991_, _10990_);
  and _62429_ (_10993_, _10992_, _03769_);
  nor _62430_ (_10994_, _10989_, _05176_);
  or _62431_ (_10995_, _10994_, _10990_);
  or _62432_ (_10996_, _10995_, _06039_);
  not _62433_ (_10997_, _05796_);
  and _62434_ (_10998_, _10997_, \oc8051_golden_model_1.P3 [7]);
  and _62435_ (_10999_, _05818_, _05796_);
  or _62436_ (_11000_, _10999_, _10998_);
  and _62437_ (_11001_, _11000_, _03512_);
  and _62438_ (_11002_, _05949_, _05200_);
  or _62439_ (_11003_, _11002_, _10990_);
  or _62440_ (_11004_, _11003_, _04444_);
  and _62441_ (_11005_, _05200_, \oc8051_golden_model_1.ACC [7]);
  or _62442_ (_11006_, _11005_, _10990_);
  and _62443_ (_11007_, _11006_, _04426_);
  and _62444_ (_11008_, _04427_, \oc8051_golden_model_1.P3 [7]);
  or _62445_ (_11009_, _11008_, _03570_);
  or _62446_ (_11010_, _11009_, _11007_);
  and _62447_ (_11011_, _11010_, _03517_);
  and _62448_ (_11012_, _11011_, _11004_);
  and _62449_ (_11013_, _05954_, _05796_);
  or _62450_ (_11014_, _11013_, _10998_);
  and _62451_ (_11015_, _11014_, _03516_);
  or _62452_ (_11016_, _11015_, _03568_);
  or _62453_ (_11017_, _11016_, _11012_);
  or _62454_ (_11018_, _10995_, _03983_);
  and _62455_ (_11019_, _11018_, _11017_);
  or _62456_ (_11020_, _11019_, _03575_);
  or _62457_ (_11021_, _11006_, _03583_);
  and _62458_ (_11022_, _11021_, _03513_);
  and _62459_ (_11023_, _11022_, _11020_);
  or _62460_ (_11024_, _11023_, _11001_);
  and _62461_ (_11025_, _11024_, _03506_);
  and _62462_ (_11026_, _05990_, _05796_);
  or _62463_ (_11027_, _11026_, _10998_);
  and _62464_ (_11028_, _11027_, _03505_);
  or _62465_ (_11029_, _11028_, _11025_);
  and _62466_ (_11030_, _11029_, _03500_);
  and _62467_ (_11031_, _10914_, _05796_);
  or _62468_ (_11032_, _11031_, _10998_);
  and _62469_ (_11033_, _11032_, _03499_);
  or _62470_ (_11034_, _11033_, _07314_);
  or _62471_ (_11035_, _11034_, _11030_);
  and _62472_ (_11036_, _11035_, _10996_);
  or _62473_ (_11037_, _11036_, _03479_);
  and _62474_ (_11038_, _05935_, _05200_);
  or _62475_ (_11039_, _10990_, _06044_);
  or _62476_ (_11040_, _11039_, _11038_);
  and _62477_ (_11041_, _11040_, _03474_);
  and _62478_ (_11042_, _11041_, _11037_);
  and _62479_ (_11043_, _10939_, _05200_);
  or _62480_ (_11044_, _11043_, _10990_);
  and _62481_ (_11045_, _11044_, _03221_);
  or _62482_ (_11046_, _11045_, _03437_);
  or _62483_ (_11047_, _11046_, _11042_);
  and _62484_ (_11048_, _06087_, _05200_);
  or _62485_ (_11049_, _11048_, _10990_);
  or _62486_ (_11050_, _11049_, _03438_);
  and _62487_ (_11051_, _11050_, _11047_);
  or _62488_ (_11052_, _11051_, _03636_);
  and _62489_ (_11053_, _06305_, _05200_);
  or _62490_ (_11054_, _11053_, _10990_);
  or _62491_ (_11055_, _11054_, _04499_);
  and _62492_ (_11056_, _11055_, _04501_);
  and _62493_ (_11057_, _11056_, _11052_);
  or _62494_ (_11058_, _11057_, _10993_);
  and _62495_ (_11059_, _11058_, _05769_);
  or _62496_ (_11060_, _10990_, _05282_);
  and _62497_ (_11061_, _11060_, _03754_);
  and _62498_ (_11062_, _11061_, _11049_);
  or _62499_ (_11063_, _11062_, _11059_);
  and _62500_ (_11064_, _11063_, _03753_);
  and _62501_ (_11065_, _11006_, _03752_);
  and _62502_ (_11066_, _11065_, _11060_);
  or _62503_ (_11067_, _11066_, _03758_);
  or _62504_ (_11068_, _11067_, _11064_);
  nor _62505_ (_11069_, _06304_, _10989_);
  or _62506_ (_11070_, _10990_, _03759_);
  or _62507_ (_11071_, _11070_, _11069_);
  and _62508_ (_11072_, _11071_, _04517_);
  and _62509_ (_11073_, _11072_, _11068_);
  nor _62510_ (_11074_, _06310_, _10989_);
  or _62511_ (_11075_, _11074_, _10990_);
  and _62512_ (_11076_, _11075_, _03760_);
  or _62513_ (_11077_, _11076_, _03790_);
  or _62514_ (_11078_, _11077_, _11073_);
  or _62515_ (_11079_, _11003_, _04192_);
  and _62516_ (_11080_, _11079_, _03152_);
  and _62517_ (_11081_, _11080_, _11078_);
  and _62518_ (_11082_, _11000_, _03151_);
  or _62519_ (_11083_, _11082_, _03520_);
  or _62520_ (_11084_, _11083_, _11081_);
  and _62521_ (_11085_, _05767_, _05200_);
  or _62522_ (_11086_, _10990_, _03521_);
  or _62523_ (_11087_, _11086_, _11085_);
  and _62524_ (_11088_, _11087_, _42963_);
  and _62525_ (_11089_, _11088_, _11084_);
  nor _62526_ (_11090_, \oc8051_golden_model_1.P3 [7], rst);
  nor _62527_ (_11091_, _11090_, _00000_);
  or _62528_ (_40535_, _11091_, _11089_);
  not _62529_ (_11092_, _05276_);
  and _62530_ (_11093_, _11092_, \oc8051_golden_model_1.P0 [7]);
  and _62531_ (_11094_, _06311_, _05276_);
  or _62532_ (_11095_, _11094_, _11093_);
  and _62533_ (_11096_, _11095_, _03769_);
  nor _62534_ (_11097_, _11092_, _05176_);
  or _62535_ (_11098_, _11097_, _11093_);
  or _62536_ (_11099_, _11098_, _06039_);
  not _62537_ (_11100_, _05205_);
  and _62538_ (_11101_, _11100_, \oc8051_golden_model_1.P0 [7]);
  and _62539_ (_11102_, _05818_, _05205_);
  or _62540_ (_11103_, _11102_, _11101_);
  and _62541_ (_11104_, _11103_, _03512_);
  and _62542_ (_11105_, _05949_, _05276_);
  or _62543_ (_11106_, _11105_, _11093_);
  or _62544_ (_11107_, _11106_, _04444_);
  and _62545_ (_11108_, _05276_, \oc8051_golden_model_1.ACC [7]);
  or _62546_ (_11109_, _11108_, _11093_);
  and _62547_ (_11110_, _11109_, _04426_);
  and _62548_ (_11111_, _04427_, \oc8051_golden_model_1.P0 [7]);
  or _62549_ (_11112_, _11111_, _03570_);
  or _62550_ (_11113_, _11112_, _11110_);
  and _62551_ (_11114_, _11113_, _03517_);
  and _62552_ (_11115_, _11114_, _11107_);
  and _62553_ (_11116_, _05954_, _05205_);
  or _62554_ (_11117_, _11116_, _11101_);
  and _62555_ (_11118_, _11117_, _03516_);
  or _62556_ (_11119_, _11118_, _03568_);
  or _62557_ (_11120_, _11119_, _11115_);
  or _62558_ (_11121_, _11098_, _03983_);
  and _62559_ (_11122_, _11121_, _11120_);
  or _62560_ (_11123_, _11122_, _03575_);
  or _62561_ (_11124_, _11109_, _03583_);
  and _62562_ (_11125_, _11124_, _03513_);
  and _62563_ (_11126_, _11125_, _11123_);
  or _62564_ (_11127_, _11126_, _11104_);
  and _62565_ (_11128_, _11127_, _03506_);
  or _62566_ (_11129_, _11101_, _05989_);
  and _62567_ (_11130_, _11129_, _03505_);
  and _62568_ (_11131_, _11130_, _11117_);
  or _62569_ (_11132_, _11131_, _11128_);
  and _62570_ (_11133_, _11132_, _03500_);
  and _62571_ (_11134_, _10914_, _05205_);
  or _62572_ (_11135_, _11134_, _11101_);
  and _62573_ (_11136_, _11135_, _03499_);
  or _62574_ (_11137_, _11136_, _07314_);
  or _62575_ (_11138_, _11137_, _11133_);
  and _62576_ (_11139_, _11138_, _11099_);
  or _62577_ (_11140_, _11139_, _03479_);
  and _62578_ (_11141_, _05935_, _05276_);
  or _62579_ (_11142_, _11093_, _06044_);
  or _62580_ (_11143_, _11142_, _11141_);
  and _62581_ (_11144_, _11143_, _03474_);
  and _62582_ (_11145_, _11144_, _11140_);
  and _62583_ (_11146_, _10939_, _05276_);
  or _62584_ (_11147_, _11146_, _11093_);
  and _62585_ (_11148_, _11147_, _03221_);
  or _62586_ (_11149_, _11148_, _03437_);
  or _62587_ (_11150_, _11149_, _11145_);
  and _62588_ (_11151_, _06087_, _05276_);
  or _62589_ (_11152_, _11151_, _11093_);
  or _62590_ (_11153_, _11152_, _03438_);
  and _62591_ (_11154_, _11153_, _11150_);
  or _62592_ (_11155_, _11154_, _03636_);
  and _62593_ (_11156_, _06305_, _05276_);
  or _62594_ (_11157_, _11156_, _11093_);
  or _62595_ (_11158_, _11157_, _04499_);
  and _62596_ (_11159_, _11158_, _04501_);
  and _62597_ (_11160_, _11159_, _11155_);
  or _62598_ (_11161_, _11160_, _11096_);
  and _62599_ (_11162_, _11161_, _05769_);
  or _62600_ (_11163_, _11093_, _05282_);
  and _62601_ (_11164_, _11163_, _03754_);
  and _62602_ (_11165_, _11164_, _11152_);
  or _62603_ (_11166_, _11165_, _11162_);
  and _62604_ (_11167_, _11166_, _03753_);
  and _62605_ (_11168_, _11109_, _03752_);
  and _62606_ (_11169_, _11168_, _11163_);
  or _62607_ (_11170_, _11169_, _03758_);
  or _62608_ (_11171_, _11170_, _11167_);
  nor _62609_ (_11172_, _06304_, _11092_);
  or _62610_ (_11173_, _11093_, _03759_);
  or _62611_ (_11174_, _11173_, _11172_);
  and _62612_ (_11175_, _11174_, _04517_);
  and _62613_ (_11176_, _11175_, _11171_);
  nor _62614_ (_11177_, _06310_, _11092_);
  or _62615_ (_11178_, _11177_, _11093_);
  and _62616_ (_11179_, _11178_, _03760_);
  or _62617_ (_11180_, _11179_, _03790_);
  or _62618_ (_11181_, _11180_, _11176_);
  or _62619_ (_11182_, _11106_, _04192_);
  and _62620_ (_11183_, _11182_, _03152_);
  and _62621_ (_11184_, _11183_, _11181_);
  and _62622_ (_11185_, _11103_, _03151_);
  or _62623_ (_11186_, _11185_, _03520_);
  or _62624_ (_11187_, _11186_, _11184_);
  and _62625_ (_11188_, _05767_, _05276_);
  or _62626_ (_11189_, _11093_, _03521_);
  or _62627_ (_11190_, _11189_, _11188_);
  and _62628_ (_11191_, _11190_, _42963_);
  and _62629_ (_11192_, _11191_, _11187_);
  nor _62630_ (_11193_, \oc8051_golden_model_1.P0 [7], rst);
  nor _62631_ (_11194_, _11193_, _00000_);
  or _62632_ (_40536_, _11194_, _11192_);
  nor _62633_ (_11195_, \oc8051_golden_model_1.P1 [7], rst);
  nor _62634_ (_11196_, _11195_, _00000_);
  not _62635_ (_11197_, _05244_);
  and _62636_ (_11198_, _11197_, \oc8051_golden_model_1.P1 [7]);
  and _62637_ (_11199_, _06311_, _05244_);
  or _62638_ (_11200_, _11199_, _11198_);
  and _62639_ (_11201_, _11200_, _03769_);
  nor _62640_ (_11202_, _11197_, _05176_);
  or _62641_ (_11203_, _11202_, _11198_);
  or _62642_ (_11204_, _11203_, _06039_);
  not _62643_ (_11205_, _05811_);
  and _62644_ (_11206_, _11205_, \oc8051_golden_model_1.P1 [7]);
  and _62645_ (_11207_, _05818_, _05811_);
  or _62646_ (_11208_, _11207_, _11206_);
  and _62647_ (_11209_, _11208_, _03512_);
  and _62648_ (_11210_, _05949_, _05244_);
  or _62649_ (_11211_, _11210_, _11198_);
  or _62650_ (_11212_, _11211_, _04444_);
  and _62651_ (_11213_, _05244_, \oc8051_golden_model_1.ACC [7]);
  or _62652_ (_11214_, _11213_, _11198_);
  and _62653_ (_11215_, _11214_, _04426_);
  and _62654_ (_11216_, _04427_, \oc8051_golden_model_1.P1 [7]);
  or _62655_ (_11217_, _11216_, _03570_);
  or _62656_ (_11218_, _11217_, _11215_);
  and _62657_ (_11219_, _11218_, _03517_);
  and _62658_ (_11220_, _11219_, _11212_);
  and _62659_ (_11221_, _05954_, _05811_);
  or _62660_ (_11222_, _11221_, _11206_);
  and _62661_ (_11223_, _11222_, _03516_);
  or _62662_ (_11224_, _11223_, _03568_);
  or _62663_ (_11225_, _11224_, _11220_);
  or _62664_ (_11226_, _11203_, _03983_);
  and _62665_ (_11227_, _11226_, _11225_);
  or _62666_ (_11228_, _11227_, _03575_);
  or _62667_ (_11229_, _11214_, _03583_);
  and _62668_ (_11230_, _11229_, _03513_);
  and _62669_ (_11231_, _11230_, _11228_);
  or _62670_ (_11232_, _11231_, _11209_);
  and _62671_ (_11233_, _11232_, _03506_);
  and _62672_ (_11234_, _05990_, _05811_);
  or _62673_ (_11235_, _11234_, _11206_);
  and _62674_ (_11236_, _11235_, _03505_);
  or _62675_ (_11237_, _11236_, _11233_);
  and _62676_ (_11238_, _11237_, _03500_);
  and _62677_ (_11239_, _10914_, _05811_);
  or _62678_ (_11240_, _11239_, _11206_);
  and _62679_ (_11241_, _11240_, _03499_);
  or _62680_ (_11242_, _11241_, _07314_);
  or _62681_ (_11243_, _11242_, _11238_);
  and _62682_ (_11244_, _11243_, _11204_);
  or _62683_ (_11245_, _11244_, _03479_);
  and _62684_ (_11246_, _05935_, _05244_);
  or _62685_ (_11247_, _11198_, _06044_);
  or _62686_ (_11248_, _11247_, _11246_);
  and _62687_ (_11249_, _11248_, _03474_);
  and _62688_ (_11250_, _11249_, _11245_);
  and _62689_ (_11251_, _10939_, _05244_);
  or _62690_ (_11252_, _11251_, _11198_);
  and _62691_ (_11253_, _11252_, _03221_);
  or _62692_ (_11254_, _11253_, _03437_);
  or _62693_ (_11255_, _11254_, _11250_);
  and _62694_ (_11256_, _06087_, _05244_);
  or _62695_ (_11257_, _11256_, _11198_);
  or _62696_ (_11258_, _11257_, _03438_);
  and _62697_ (_11259_, _11258_, _11255_);
  or _62698_ (_11260_, _11259_, _03636_);
  and _62699_ (_11261_, _06305_, _05244_);
  or _62700_ (_11262_, _11261_, _11198_);
  or _62701_ (_11263_, _11262_, _04499_);
  and _62702_ (_11264_, _11263_, _04501_);
  and _62703_ (_11265_, _11264_, _11260_);
  or _62704_ (_11266_, _11265_, _11201_);
  and _62705_ (_11267_, _11266_, _05769_);
  or _62706_ (_11268_, _11198_, _05282_);
  and _62707_ (_11269_, _11268_, _03754_);
  and _62708_ (_11270_, _11269_, _11257_);
  or _62709_ (_11271_, _11270_, _11267_);
  and _62710_ (_11272_, _11271_, _03753_);
  and _62711_ (_11273_, _11214_, _03752_);
  and _62712_ (_11274_, _11273_, _11268_);
  or _62713_ (_11275_, _11274_, _03758_);
  or _62714_ (_11276_, _11275_, _11272_);
  nor _62715_ (_11277_, _06304_, _11197_);
  or _62716_ (_11278_, _11198_, _03759_);
  or _62717_ (_11279_, _11278_, _11277_);
  and _62718_ (_11280_, _11279_, _04517_);
  and _62719_ (_11281_, _11280_, _11276_);
  nor _62720_ (_11282_, _06310_, _11197_);
  or _62721_ (_11283_, _11282_, _11198_);
  and _62722_ (_11284_, _11283_, _03760_);
  or _62723_ (_11285_, _11284_, _03790_);
  or _62724_ (_11286_, _11285_, _11281_);
  or _62725_ (_11287_, _11211_, _04192_);
  and _62726_ (_11288_, _11287_, _03152_);
  and _62727_ (_11289_, _11288_, _11286_);
  and _62728_ (_11290_, _11208_, _03151_);
  or _62729_ (_11291_, _11290_, _03520_);
  or _62730_ (_11292_, _11291_, _11289_);
  and _62731_ (_11293_, _05767_, _05244_);
  or _62732_ (_11294_, _11198_, _03521_);
  or _62733_ (_11295_, _11294_, _11293_);
  and _62734_ (_11296_, _11295_, _42963_);
  and _62735_ (_11297_, _11296_, _11292_);
  or _62736_ (_40538_, _11297_, _11196_);
  not _62737_ (_11298_, \oc8051_golden_model_1.SP [7]);
  nor _62738_ (_11299_, _42963_, _11298_);
  and _62739_ (_11300_, _04849_, \oc8051_golden_model_1.SP [4]);
  and _62740_ (_11301_, _11300_, \oc8051_golden_model_1.SP [5]);
  and _62741_ (_11302_, _11301_, \oc8051_golden_model_1.SP [6]);
  or _62742_ (_11303_, _11302_, \oc8051_golden_model_1.SP [7]);
  nand _62743_ (_11304_, _11302_, \oc8051_golden_model_1.SP [7]);
  and _62744_ (_11305_, _11304_, _11303_);
  or _62745_ (_11306_, _11305_, _04533_);
  nor _62746_ (_11307_, _05269_, _11298_);
  and _62747_ (_11308_, _06311_, _05269_);
  or _62748_ (_11309_, _11308_, _11307_);
  and _62749_ (_11310_, _11309_, _03769_);
  and _62750_ (_11311_, _05949_, _05269_);
  or _62751_ (_11312_, _11311_, _11307_);
  or _62752_ (_11313_, _11312_, _04444_);
  nor _62753_ (_11314_, _04426_, _11298_);
  and _62754_ (_11315_, _05269_, \oc8051_golden_model_1.ACC [7]);
  or _62755_ (_11316_, _11315_, _11307_);
  and _62756_ (_11317_, _11316_, _04426_);
  or _62757_ (_11318_, _11317_, _11314_);
  and _62758_ (_11319_, _11318_, _04762_);
  and _62759_ (_11320_, _11305_, _03923_);
  or _62760_ (_11321_, _11320_, _03570_);
  or _62761_ (_11322_, _11321_, _11319_);
  and _62762_ (_11323_, _11322_, _03203_);
  and _62763_ (_11324_, _11323_, _11313_);
  and _62764_ (_11325_, _11305_, _04746_);
  or _62765_ (_11326_, _11325_, _03568_);
  or _62766_ (_11327_, _11326_, _11324_);
  not _62767_ (_11328_, \oc8051_golden_model_1.SP [6]);
  not _62768_ (_11329_, \oc8051_golden_model_1.SP [5]);
  not _62769_ (_11330_, \oc8051_golden_model_1.SP [4]);
  and _62770_ (_11331_, _05852_, _11330_);
  and _62771_ (_11332_, _11331_, _11329_);
  and _62772_ (_11333_, _11332_, _11328_);
  and _62773_ (_11334_, _11333_, _03502_);
  nor _62774_ (_11335_, _11334_, _11298_);
  and _62775_ (_11336_, _11334_, _11298_);
  nor _62776_ (_11337_, _11336_, _11335_);
  nand _62777_ (_11338_, _11337_, _03568_);
  and _62778_ (_11339_, _11338_, _11327_);
  or _62779_ (_11340_, _11339_, _03575_);
  or _62780_ (_11341_, _11316_, _03583_);
  and _62781_ (_11342_, _11341_, _04887_);
  and _62782_ (_11343_, _11342_, _11340_);
  and _62783_ (_11344_, _11301_, \oc8051_golden_model_1.SP [0]);
  and _62784_ (_11345_, _11344_, \oc8051_golden_model_1.SP [6]);
  or _62785_ (_11346_, _11345_, \oc8051_golden_model_1.SP [7]);
  nand _62786_ (_11347_, _11345_, \oc8051_golden_model_1.SP [7]);
  and _62787_ (_11348_, _11347_, _11346_);
  and _62788_ (_11349_, _11348_, _03511_);
  or _62789_ (_11350_, _11349_, _04744_);
  or _62790_ (_11351_, _11350_, _11343_);
  or _62791_ (_11352_, _11305_, _04745_);
  and _62792_ (_11353_, _11352_, _06039_);
  and _62793_ (_11354_, _11353_, _11351_);
  not _62794_ (_11355_, _05269_);
  nor _62795_ (_11356_, _11355_, _05176_);
  or _62796_ (_11357_, _11356_, _11307_);
  and _62797_ (_11358_, _11357_, _07314_);
  or _62798_ (_11359_, _11358_, _03479_);
  or _62799_ (_11360_, _11359_, _11354_);
  and _62800_ (_11361_, _05935_, _05269_);
  or _62801_ (_11362_, _11307_, _06044_);
  or _62802_ (_11363_, _11362_, _11361_);
  and _62803_ (_11364_, _11363_, _03474_);
  and _62804_ (_11365_, _11364_, _11360_);
  nor _62805_ (_11366_, _06292_, _11355_);
  or _62806_ (_11367_, _11366_, _11307_);
  and _62807_ (_11368_, _11367_, _03221_);
  or _62808_ (_11369_, _11368_, _03437_);
  or _62809_ (_11370_, _11369_, _11365_);
  and _62810_ (_11371_, _06087_, _05269_);
  or _62811_ (_11372_, _11371_, _11307_);
  or _62812_ (_11373_, _11372_, _03438_);
  and _62813_ (_11374_, _11373_, _11370_);
  or _62814_ (_11375_, _11374_, _03189_);
  not _62815_ (_11376_, _03189_);
  or _62816_ (_11377_, _11305_, _11376_);
  and _62817_ (_11378_, _11377_, _11375_);
  or _62818_ (_11379_, _11378_, _03636_);
  and _62819_ (_11380_, _06305_, _05269_);
  or _62820_ (_11381_, _11380_, _11307_);
  or _62821_ (_11382_, _11381_, _04499_);
  and _62822_ (_11383_, _11382_, _04501_);
  and _62823_ (_11384_, _11383_, _11379_);
  or _62824_ (_11385_, _11384_, _11310_);
  and _62825_ (_11386_, _11385_, _05769_);
  or _62826_ (_11387_, _11307_, _05282_);
  and _62827_ (_11388_, _11387_, _03754_);
  and _62828_ (_11389_, _11388_, _11372_);
  or _62829_ (_11390_, _11389_, _11386_);
  and _62830_ (_11391_, _11390_, _09960_);
  and _62831_ (_11392_, _11316_, _03752_);
  and _62832_ (_11393_, _11392_, _11387_);
  and _62833_ (_11394_, _11305_, _03192_);
  or _62834_ (_11395_, _11394_, _03758_);
  or _62835_ (_11396_, _11395_, _11393_);
  or _62836_ (_11397_, _11396_, _11391_);
  nor _62837_ (_11398_, _06304_, _11355_);
  or _62838_ (_11399_, _11398_, _11307_);
  or _62839_ (_11400_, _11399_, _03759_);
  and _62840_ (_11401_, _11400_, _11397_);
  or _62841_ (_11402_, _11401_, _03760_);
  not _62842_ (_11403_, _03775_);
  nor _62843_ (_11404_, _06310_, _11355_);
  or _62844_ (_11405_, _11307_, _04517_);
  or _62845_ (_11406_, _11405_, _11404_);
  and _62846_ (_11407_, _11406_, _11403_);
  and _62847_ (_11408_, _11407_, _11402_);
  or _62848_ (_11409_, _11333_, \oc8051_golden_model_1.SP [7]);
  nand _62849_ (_11410_, _11333_, \oc8051_golden_model_1.SP [7]);
  and _62850_ (_11411_, _11410_, _11409_);
  and _62851_ (_11412_, _11411_, _03775_);
  or _62852_ (_11413_, _11412_, _03179_);
  or _62853_ (_11414_, _11413_, _11408_);
  or _62854_ (_11415_, _11305_, _06328_);
  and _62855_ (_11416_, _11415_, _11414_);
  or _62856_ (_11417_, _11416_, _03522_);
  or _62857_ (_11418_, _11411_, _03523_);
  and _62858_ (_11419_, _11418_, _04192_);
  and _62859_ (_11420_, _11419_, _11417_);
  and _62860_ (_11421_, _11312_, _03790_);
  or _62861_ (_11422_, _11421_, _04947_);
  or _62862_ (_11423_, _11422_, _11420_);
  and _62863_ (_11424_, _11423_, _11306_);
  or _62864_ (_11425_, _11424_, _03520_);
  and _62865_ (_11426_, _05767_, _05269_);
  or _62866_ (_11427_, _11307_, _03521_);
  or _62867_ (_11428_, _11427_, _11426_);
  and _62868_ (_11429_, _11428_, _42963_);
  and _62869_ (_11430_, _11429_, _11425_);
  or _62870_ (_11431_, _11430_, _11299_);
  and _62871_ (_40539_, _11431_, _41755_);
  nor _62872_ (_11432_, _42963_, _07888_);
  nor _62873_ (_11433_, _05783_, _07888_);
  and _62874_ (_11434_, _05818_, _05783_);
  or _62875_ (_11435_, _11434_, _11433_);
  or _62876_ (_11436_, _11435_, _03152_);
  not _62877_ (_11437_, _07782_);
  nor _62878_ (_11438_, _07818_, _07783_);
  nor _62879_ (_11439_, _11438_, _07780_);
  nand _62880_ (_11440_, _11439_, _11437_);
  and _62881_ (_11441_, _07851_, _07847_);
  and _62882_ (_11442_, _11441_, _06700_);
  nor _62883_ (_11443_, _07836_, _05834_);
  or _62884_ (_11444_, _11443_, _07905_);
  or _62885_ (_11445_, _11444_, _11442_);
  or _62886_ (_11446_, _11445_, _07830_);
  nor _62887_ (_11447_, _05218_, _07888_);
  and _62888_ (_11448_, _06311_, _05218_);
  or _62889_ (_11449_, _11448_, _11447_);
  and _62890_ (_11450_, _11449_, _03769_);
  not _62891_ (_11451_, _05218_);
  nor _62892_ (_11452_, _06292_, _11451_);
  or _62893_ (_11453_, _11452_, _11447_);
  and _62894_ (_11454_, _11453_, _03221_);
  nor _62895_ (_11455_, _11451_, _05176_);
  or _62896_ (_11456_, _11455_, _11447_);
  or _62897_ (_11457_, _11456_, _06039_);
  and _62898_ (_11458_, _08048_, _06713_);
  and _62899_ (_11459_, _11458_, _05935_);
  and _62900_ (_11460_, _08051_, _08044_);
  nor _62901_ (_11461_, _11460_, _08042_);
  nand _62902_ (_11462_, _08098_, _08044_);
  or _62903_ (_11463_, _11462_, _08096_);
  and _62904_ (_11464_, _11463_, _11461_);
  or _62905_ (_11465_, _11464_, _08037_);
  or _62906_ (_11466_, _11465_, _11459_);
  not _62907_ (_11467_, _03606_);
  nor _62908_ (_11468_, _10794_, _10419_);
  and _62909_ (_11469_, _10083_, _07888_);
  not _62910_ (_11470_, _08625_);
  nor _62911_ (_11471_, _10374_, _11470_);
  or _62912_ (_11472_, _11471_, _08623_);
  and _62913_ (_11473_, _11472_, _10372_);
  not _62914_ (_11474_, _10370_);
  and _62915_ (_11475_, _08620_, _11474_);
  or _62916_ (_11476_, _11475_, _10369_);
  or _62917_ (_11477_, _11476_, _11473_);
  and _62918_ (_11478_, _11477_, _10381_);
  not _62919_ (_11479_, _08609_);
  or _62920_ (_11480_, _08613_, _08608_);
  and _62921_ (_11481_, _11480_, _11479_);
  and _62922_ (_11482_, _11481_, _10380_);
  nor _62923_ (_11483_, _05984_, \oc8051_golden_model_1.ACC [7]);
  and _62924_ (_11484_, _08604_, _10379_);
  or _62925_ (_11485_, _11484_, _11483_);
  or _62926_ (_11486_, _11485_, _11482_);
  or _62927_ (_11487_, _11486_, _11478_);
  nor _62928_ (_11488_, _10382_, _03998_);
  and _62929_ (_11489_, _11488_, _11487_);
  nor _62930_ (_11490_, _04284_, \oc8051_golden_model_1.ACC [1]);
  and _62931_ (_11491_, _04284_, \oc8051_golden_model_1.ACC [1]);
  and _62932_ (_11492_, _03471_, \oc8051_golden_model_1.ACC [0]);
  nor _62933_ (_11493_, _11492_, _11491_);
  or _62934_ (_11494_, _11493_, _11490_);
  and _62935_ (_11495_, _11494_, _10393_);
  nand _62936_ (_11496_, _03432_, \oc8051_golden_model_1.ACC [3]);
  nor _62937_ (_11497_, _03432_, \oc8051_golden_model_1.ACC [3]);
  nor _62938_ (_11498_, _03877_, \oc8051_golden_model_1.ACC [2]);
  or _62939_ (_11499_, _11498_, _11497_);
  and _62940_ (_11500_, _11499_, _11496_);
  or _62941_ (_11501_, _11500_, _11495_);
  and _62942_ (_11502_, _11501_, _10391_);
  nand _62943_ (_11503_, _03834_, \oc8051_golden_model_1.ACC [5]);
  nor _62944_ (_11504_, _03834_, \oc8051_golden_model_1.ACC [5]);
  nor _62945_ (_11505_, _04249_, \oc8051_golden_model_1.ACC [4]);
  or _62946_ (_11506_, _11505_, _11504_);
  and _62947_ (_11507_, _11506_, _11503_);
  and _62948_ (_11508_, _11507_, _10390_);
  and _62949_ (_11509_, _03401_, _05834_);
  or _62950_ (_11510_, _03561_, \oc8051_golden_model_1.ACC [6]);
  nor _62951_ (_11511_, _11510_, _08422_);
  or _62952_ (_11512_, _11511_, _11509_);
  or _62953_ (_11513_, _11512_, _11508_);
  or _62954_ (_11514_, _11513_, _11502_);
  and _62955_ (_11515_, _11514_, _03638_);
  and _62956_ (_11516_, _11515_, _10399_);
  or _62957_ (_11517_, _11516_, _11489_);
  or _62958_ (_11518_, _11517_, _11469_);
  not _62959_ (_11519_, _10324_);
  or _62960_ (_11520_, _10333_, _10329_);
  and _62961_ (_11521_, _11520_, _05177_);
  or _62962_ (_11522_, _10340_, _10336_);
  and _62963_ (_11523_, _10338_, _11522_);
  and _62964_ (_11524_, _11523_, _10335_);
  or _62965_ (_11525_, _11524_, _11521_);
  or _62966_ (_11526_, _10356_, _10354_);
  and _62967_ (_11527_, _11526_, _10351_);
  and _62968_ (_11528_, _10348_, _10346_);
  or _62969_ (_11529_, _11528_, _10345_);
  or _62970_ (_11530_, _11529_, _11527_);
  and _62971_ (_11531_, _11530_, _10344_);
  nor _62972_ (_11532_, _11531_, _11525_);
  nor _62973_ (_11533_, _11532_, _10360_);
  or _62974_ (_11534_, _11533_, _11519_);
  and _62975_ (_11535_, _05949_, _05218_);
  or _62976_ (_11536_, _11535_, _11447_);
  or _62977_ (_11537_, _11536_, _04444_);
  not _62978_ (_11538_, _07948_);
  and _62979_ (_11539_, _05218_, \oc8051_golden_model_1.ACC [7]);
  or _62980_ (_11540_, _11539_, _11447_);
  and _62981_ (_11541_, _11540_, _04426_);
  nor _62982_ (_11542_, _04426_, _07888_);
  or _62983_ (_11543_, _11542_, _03570_);
  or _62984_ (_11544_, _11543_, _11541_);
  and _62985_ (_11545_, _11544_, _11538_);
  and _62986_ (_11546_, _11545_, _11537_);
  nor _62987_ (_11547_, _07958_, \oc8051_golden_model_1.PSW [7]);
  not _62988_ (_11548_, _11547_);
  nor _62989_ (_11549_, _11548_, _07968_);
  nor _62990_ (_11550_, _11549_, _11538_);
  not _62991_ (_11551_, _10254_);
  nand _62992_ (_11552_, _11551_, _03576_);
  or _62993_ (_11553_, _11552_, _11550_);
  or _62994_ (_11554_, _11553_, _11546_);
  and _62995_ (_11555_, _05954_, _05783_);
  or _62996_ (_11556_, _11555_, _11433_);
  or _62997_ (_11557_, _11556_, _03517_);
  or _62998_ (_11558_, _11456_, _03983_);
  and _62999_ (_11559_, _11558_, _11557_);
  and _63000_ (_11560_, _11559_, _11554_);
  or _63001_ (_11561_, _11560_, _03575_);
  or _63002_ (_11562_, _11540_, _03583_);
  nor _63003_ (_11563_, _10315_, _03512_);
  and _63004_ (_11564_, _11563_, _11562_);
  and _63005_ (_11565_, _11564_, _11561_);
  and _63006_ (_11566_, _11435_, _03512_);
  or _63007_ (_11567_, _11566_, _10324_);
  or _63008_ (_11568_, _11567_, _11565_);
  and _63009_ (_11569_, _11568_, _11534_);
  or _63010_ (_11570_, _11569_, _10323_);
  and _63011_ (_11571_, _04004_, _03504_);
  and _63012_ (_11572_, _03654_, _03219_);
  and _63013_ (_11573_, _11572_, _03504_);
  nor _63014_ (_11574_, _11573_, _11571_);
  not _63015_ (_11575_, _10323_);
  or _63016_ (_11576_, _11533_, _11575_);
  and _63017_ (_11577_, _11576_, _11574_);
  and _63018_ (_11578_, _11577_, _11570_);
  not _63019_ (_11579_, _10106_);
  nand _63020_ (_11580_, _11579_, _10103_);
  nand _63021_ (_11581_, _11580_, _10102_);
  not _63022_ (_11582_, _10110_);
  and _63023_ (_11583_, _11582_, _10108_);
  or _63024_ (_11584_, _11583_, _11581_);
  and _63025_ (_11585_, _11584_, _10101_);
  not _63026_ (_11586_, _10097_);
  nand _63027_ (_11587_, _11586_, _10094_);
  nand _63028_ (_11588_, _11587_, _10090_);
  and _63029_ (_11589_, _11588_, _06005_);
  or _63030_ (_11590_, _11589_, _10115_);
  or _63031_ (_11591_, _11590_, _11585_);
  nor _63032_ (_11592_, _10116_, _10328_);
  and _63033_ (_11593_, _11592_, _11591_);
  or _63034_ (_11594_, _11593_, _11578_);
  nor _63035_ (_11595_, _03638_, _03527_);
  and _63036_ (_11596_, _11595_, _10084_);
  and _63037_ (_11597_, _11596_, _11594_);
  or _63038_ (_11598_, _11597_, _11518_);
  and _63039_ (_11599_, _11598_, _03593_);
  and _63040_ (_11600_, _05801_, \oc8051_golden_model_1.P2 [2]);
  and _63041_ (_11601_, _05796_, \oc8051_golden_model_1.P3 [2]);
  nor _63042_ (_11602_, _11601_, _11600_);
  and _63043_ (_11603_, _05205_, \oc8051_golden_model_1.P0 [2]);
  and _63044_ (_11604_, _05811_, \oc8051_golden_model_1.P1 [2]);
  nor _63045_ (_11605_, _11604_, _11603_);
  and _63046_ (_11606_, _11605_, _11602_);
  and _63047_ (_11607_, _11606_, _10617_);
  and _63048_ (_11608_, _11607_, _10614_);
  and _63049_ (_11609_, _11608_, _05619_);
  nor _63050_ (_11610_, _11609_, _10604_);
  and _63051_ (_11611_, _05205_, \oc8051_golden_model_1.P0 [1]);
  and _63052_ (_11612_, _05811_, \oc8051_golden_model_1.P1 [1]);
  nor _63053_ (_11613_, _11612_, _11611_);
  and _63054_ (_11614_, _05796_, \oc8051_golden_model_1.P3 [1]);
  and _63055_ (_11615_, _05801_, \oc8051_golden_model_1.P2 [1]);
  or _63056_ (_11616_, _11615_, _11614_);
  nor _63057_ (_11617_, _11616_, _10633_);
  and _63058_ (_11618_, _11617_, _10643_);
  and _63059_ (_11619_, _11618_, _10632_);
  and _63060_ (_11620_, _11619_, _11613_);
  and _63061_ (_11621_, _11620_, _05522_);
  nor _63062_ (_11622_, _11621_, _10629_);
  nor _63063_ (_11623_, _11622_, _11610_);
  and _63064_ (_11624_, _05205_, \oc8051_golden_model_1.P0 [4]);
  and _63065_ (_11625_, _05811_, \oc8051_golden_model_1.P1 [4]);
  nor _63066_ (_11626_, _11625_, _11624_);
  and _63067_ (_11627_, _05796_, \oc8051_golden_model_1.P3 [4]);
  and _63068_ (_11628_, _05801_, \oc8051_golden_model_1.P2 [4]);
  or _63069_ (_11629_, _11628_, _11627_);
  nor _63070_ (_11630_, _11629_, _10659_);
  and _63071_ (_11631_, _11630_, _10669_);
  and _63072_ (_11632_, _11631_, _10658_);
  and _63073_ (_11633_, _11632_, _11626_);
  and _63074_ (_11634_, _11633_, _05713_);
  nor _63075_ (_11635_, _10655_, _11634_);
  nor _63076_ (_11636_, _11635_, _05988_);
  and _63077_ (_11637_, _11636_, _11623_);
  and _63078_ (_11638_, _05801_, \oc8051_golden_model_1.P2 [0]);
  and _63079_ (_11639_, _05796_, \oc8051_golden_model_1.P3 [0]);
  nor _63080_ (_11640_, _11639_, _11638_);
  and _63081_ (_11641_, _05205_, \oc8051_golden_model_1.P0 [0]);
  and _63082_ (_11642_, _05811_, \oc8051_golden_model_1.P1 [0]);
  nor _63083_ (_11643_, _11642_, _11641_);
  and _63084_ (_11644_, _11643_, _11640_);
  and _63085_ (_11645_, _11644_, _10696_);
  and _63086_ (_11646_, _11645_, _10693_);
  and _63087_ (_11647_, _11646_, _05570_);
  nor _63088_ (_11648_, _11647_, _10682_);
  and _63089_ (_11649_, _05801_, \oc8051_golden_model_1.P2 [6]);
  and _63090_ (_11650_, _05796_, \oc8051_golden_model_1.P3 [6]);
  nor _63091_ (_11651_, _11650_, _11649_);
  and _63092_ (_11652_, _05205_, \oc8051_golden_model_1.P0 [6]);
  and _63093_ (_11653_, _05811_, \oc8051_golden_model_1.P1 [6]);
  nor _63094_ (_11654_, _11653_, _11652_);
  and _63095_ (_11655_, _11654_, _11651_);
  and _63096_ (_11656_, _11655_, _10725_);
  and _63097_ (_11657_, _11656_, _10721_);
  and _63098_ (_11658_, _11657_, _05328_);
  nor _63099_ (_11659_, _10710_, _11658_);
  nor _63100_ (_11660_, _11659_, _11648_);
  and _63101_ (_11661_, _05205_, \oc8051_golden_model_1.P0 [3]);
  and _63102_ (_11662_, _05811_, \oc8051_golden_model_1.P1 [3]);
  nor _63103_ (_11663_, _11662_, _11661_);
  and _63104_ (_11664_, _05796_, \oc8051_golden_model_1.P3 [3]);
  and _63105_ (_11665_, _05801_, \oc8051_golden_model_1.P2 [3]);
  or _63106_ (_11666_, _11665_, _11664_);
  nor _63107_ (_11667_, _11666_, _10758_);
  and _63108_ (_11668_, _11667_, _10747_);
  and _63109_ (_11669_, _11668_, _10757_);
  and _63110_ (_11670_, _11669_, _11663_);
  and _63111_ (_11671_, _11670_, _05473_);
  nor _63112_ (_11672_, _11671_, _10739_);
  and _63113_ (_11673_, _05801_, \oc8051_golden_model_1.P2 [5]);
  and _63114_ (_11674_, _05796_, \oc8051_golden_model_1.P3 [5]);
  nor _63115_ (_11675_, _11674_, _11673_);
  and _63116_ (_11676_, _05205_, \oc8051_golden_model_1.P0 [5]);
  and _63117_ (_11677_, _05811_, \oc8051_golden_model_1.P1 [5]);
  nor _63118_ (_11678_, _11677_, _11676_);
  and _63119_ (_11679_, _11678_, _11675_);
  and _63120_ (_11680_, _11679_, _10780_);
  and _63121_ (_11681_, _11680_, _10777_);
  and _63122_ (_11682_, _11681_, _05423_);
  nor _63123_ (_11683_, _10767_, _11682_);
  nor _63124_ (_11684_, _11683_, _11672_);
  and _63125_ (_11685_, _11684_, _11660_);
  and _63126_ (_11686_, _11685_, _11637_);
  and _63127_ (_11687_, _11686_, \oc8051_golden_model_1.PSW [7]);
  and _63128_ (_11688_, _11687_, _03592_);
  or _63129_ (_11689_, _11433_, _05989_);
  and _63130_ (_11690_, _11689_, _03505_);
  and _63131_ (_11691_, _11690_, _11556_);
  or _63132_ (_11692_, _11691_, _11688_);
  or _63133_ (_11693_, _11692_, _11599_);
  nor _63134_ (_11694_, _06794_, _03607_);
  and _63135_ (_11695_, _11694_, _11693_);
  or _63136_ (_11696_, _11695_, _11468_);
  and _63137_ (_11697_, _11696_, _11467_);
  nand _63138_ (_11698_, _03484_, _03222_);
  or _63139_ (_11699_, _03666_, _03253_);
  nand _63140_ (_11700_, _11699_, _11698_);
  or _63141_ (_11701_, _11686_, \oc8051_golden_model_1.PSW [7]);
  and _63142_ (_11702_, _11701_, _03606_);
  or _63143_ (_11703_, _11702_, _11700_);
  or _63144_ (_11704_, _11703_, _11697_);
  and _63145_ (_11705_, _03650_, _03222_);
  not _63146_ (_11706_, _11705_);
  and _63147_ (_11707_, _07844_, _07839_);
  nor _63148_ (_11708_, _11707_, _07837_);
  nand _63149_ (_11709_, _07845_, _07839_);
  or _63150_ (_11710_, _11709_, _08027_);
  and _63151_ (_11711_, _11710_, _11708_);
  or _63152_ (_11712_, _11711_, _11442_);
  and _63153_ (_11713_, _11712_, _11706_);
  or _63154_ (_11714_, _11713_, _07922_);
  and _63155_ (_11715_, _11714_, _11704_);
  and _63156_ (_11716_, _11712_, _11705_);
  or _63157_ (_11717_, _11716_, _08035_);
  or _63158_ (_11718_, _11717_, _11715_);
  and _63159_ (_11719_, _11718_, _11466_);
  or _63160_ (_11720_, _11719_, _03614_);
  not _63161_ (_11721_, _05984_);
  and _63162_ (_11722_, _08237_, _08235_);
  and _63163_ (_11723_, _11722_, _08126_);
  and _63164_ (_11724_, _11723_, _11721_);
  and _63165_ (_11725_, _08234_, _08231_);
  nor _63166_ (_11726_, _11725_, _08229_);
  and _63167_ (_11727_, _08279_, _08231_);
  nand _63168_ (_11728_, _11727_, _08277_);
  and _63169_ (_11729_, _11728_, _11726_);
  or _63170_ (_11730_, _11729_, _11724_);
  or _63171_ (_11731_, _11730_, _03619_);
  and _63172_ (_11732_, _11731_, _08109_);
  and _63173_ (_11733_, _11732_, _11720_);
  and _63174_ (_11734_, _08289_, _05220_);
  and _63175_ (_11735_, _08301_, _08297_);
  nor _63176_ (_11736_, _11735_, _08295_);
  nand _63177_ (_11737_, _08345_, _08297_);
  or _63178_ (_11738_, _11737_, _08343_);
  and _63179_ (_11739_, _11738_, _11736_);
  or _63180_ (_11740_, _11739_, _11734_);
  and _63181_ (_11741_, _11740_, _08108_);
  or _63182_ (_11742_, _11741_, _07314_);
  or _63183_ (_11743_, _11742_, _11733_);
  and _63184_ (_11744_, _11743_, _11457_);
  or _63185_ (_11745_, _11744_, _03479_);
  and _63186_ (_11746_, _05935_, _05218_);
  or _63187_ (_11747_, _11447_, _06044_);
  or _63188_ (_11748_, _11747_, _11746_);
  and _63189_ (_11749_, _11748_, _03474_);
  and _63190_ (_11750_, _11749_, _11745_);
  or _63191_ (_11751_, _11750_, _11454_);
  nor _63192_ (_11752_, _07328_, _03745_);
  and _63193_ (_11753_, _11752_, _11751_);
  nor _63194_ (_11754_, _11686_, _07888_);
  and _63195_ (_11755_, _11754_, _03745_);
  or _63196_ (_11756_, _11755_, _03437_);
  or _63197_ (_11757_, _11756_, _11753_);
  and _63198_ (_11758_, _06087_, _05218_);
  or _63199_ (_11759_, _11758_, _11447_);
  or _63200_ (_11760_, _11759_, _03438_);
  and _63201_ (_11761_, _11760_, _11757_);
  or _63202_ (_11762_, _11761_, _03744_);
  nand _63203_ (_11763_, _11686_, _07888_);
  or _63204_ (_11764_, _11763_, _04118_);
  and _63205_ (_11765_, _11764_, _11762_);
  or _63206_ (_11766_, _11765_, _03636_);
  and _63207_ (_11767_, _06305_, _05218_);
  or _63208_ (_11768_, _11767_, _11447_);
  or _63209_ (_11769_, _11768_, _04499_);
  and _63210_ (_11770_, _11769_, _04501_);
  and _63211_ (_11771_, _11770_, _11766_);
  or _63212_ (_11772_, _11771_, _11450_);
  and _63213_ (_11773_, _11772_, _05769_);
  or _63214_ (_11774_, _11447_, _05282_);
  and _63215_ (_11775_, _11774_, _03754_);
  and _63216_ (_11776_, _11775_, _11759_);
  or _63217_ (_11777_, _11776_, _11773_);
  and _63218_ (_11778_, _11777_, _03753_);
  and _63219_ (_11779_, _11540_, _03752_);
  and _63220_ (_11780_, _11779_, _11774_);
  or _63221_ (_11781_, _11780_, _03758_);
  or _63222_ (_11782_, _11781_, _11778_);
  nor _63223_ (_11783_, _06304_, _11451_);
  or _63224_ (_11784_, _11447_, _03759_);
  or _63225_ (_11785_, _11784_, _11783_);
  and _63226_ (_11786_, _11785_, _04517_);
  and _63227_ (_11787_, _11786_, _11782_);
  nor _63228_ (_11788_, _06310_, _11451_);
  or _63229_ (_11789_, _11788_, _11447_);
  and _63230_ (_11790_, _11789_, _03760_);
  or _63231_ (_11791_, _11790_, _08490_);
  or _63232_ (_11792_, _11791_, _11787_);
  and _63233_ (_11793_, _11792_, _11446_);
  or _63234_ (_11794_, _11793_, _07825_);
  or _63235_ (_11795_, _08495_, _11459_);
  nor _63236_ (_11796_, _08041_, _05834_);
  or _63237_ (_11797_, _11796_, _08517_);
  or _63238_ (_11798_, _11797_, _11795_);
  and _63239_ (_11799_, _11798_, _03766_);
  and _63240_ (_11800_, _11799_, _11794_);
  nor _63241_ (_11801_, _08228_, _05834_);
  or _63242_ (_11802_, _11801_, _08549_);
  or _63243_ (_11803_, _11802_, _11724_);
  and _63244_ (_11804_, _11803_, _03765_);
  or _63245_ (_11805_, _11804_, _11800_);
  or _63246_ (_11806_, _11805_, _08523_);
  nor _63247_ (_11807_, _08294_, _05834_);
  or _63248_ (_11808_, _11807_, _08579_);
  or _63249_ (_11809_, _11808_, _11734_);
  or _63250_ (_11810_, _11809_, _08557_);
  and _63251_ (_11811_, _11810_, _08556_);
  and _63252_ (_11812_, _11811_, _11806_);
  nand _63253_ (_11813_, _08555_, \oc8051_golden_model_1.ACC [7]);
  nand _63254_ (_11814_, _11813_, _07780_);
  or _63255_ (_11815_, _11814_, _11812_);
  and _63256_ (_11816_, _11815_, _11440_);
  or _63257_ (_11817_, _11816_, _07731_);
  and _63258_ (_11818_, _07768_, _07735_);
  not _63259_ (_11819_, _07733_);
  and _63260_ (_11820_, _07736_, _11819_);
  or _63261_ (_11821_, _07734_, _07732_);
  or _63262_ (_11822_, _11821_, _11820_);
  or _63263_ (_11823_, _11822_, _11818_);
  and _63264_ (_11824_, _11823_, _03526_);
  and _63265_ (_11825_, _11824_, _11817_);
  not _63266_ (_11826_, _08599_);
  not _63267_ (_11827_, _08600_);
  nand _63268_ (_11828_, _08639_, _11827_);
  and _63269_ (_11829_, _11828_, _03524_);
  and _63270_ (_11830_, _11829_, _11826_);
  or _63271_ (_11831_, _11830_, _08597_);
  or _63272_ (_11832_, _11831_, _11825_);
  not _63273_ (_11833_, _08421_);
  or _63274_ (_11834_, _08678_, _08420_);
  and _63275_ (_11835_, _11834_, _08597_);
  nand _63276_ (_11836_, _11835_, _11833_);
  and _63277_ (_11837_, _11836_, _11832_);
  or _63278_ (_11838_, _11837_, _03790_);
  not _63279_ (_11839_, _08692_);
  or _63280_ (_11840_, _11536_, _04192_);
  and _63281_ (_11841_, _11840_, _11839_);
  and _63282_ (_11842_, _11841_, _11838_);
  and _63283_ (_11843_, _08692_, \oc8051_golden_model_1.ACC [0]);
  or _63284_ (_11844_, _11843_, _03151_);
  or _63285_ (_11845_, _11844_, _11842_);
  and _63286_ (_11846_, _11845_, _11436_);
  or _63287_ (_11847_, _11846_, _03520_);
  and _63288_ (_11848_, _05767_, _05218_);
  or _63289_ (_11849_, _11447_, _03521_);
  or _63290_ (_11850_, _11849_, _11848_);
  and _63291_ (_11851_, _11850_, _42963_);
  and _63292_ (_11852_, _11851_, _11847_);
  or _63293_ (_11853_, _11852_, _11432_);
  and _63294_ (_40540_, _11853_, _41755_);
  and _63295_ (_11854_, _42967_, \oc8051_golden_model_1.P0INREG [7]);
  or _63296_ (_11855_, _11854_, _00862_);
  and _63297_ (_40541_, _11855_, _41755_);
  and _63298_ (_11856_, _42967_, \oc8051_golden_model_1.P1INREG [7]);
  or _63299_ (_11857_, _11856_, _00969_);
  and _63300_ (_40542_, _11857_, _41755_);
  and _63301_ (_11858_, _42967_, \oc8051_golden_model_1.P2INREG [7]);
  or _63302_ (_11859_, _11858_, _00934_);
  and _63303_ (_40544_, _11859_, _41755_);
  and _63304_ (_11860_, _42967_, \oc8051_golden_model_1.P3INREG [7]);
  or _63305_ (_11861_, _11860_, _01115_);
  and _63306_ (_40545_, _11861_, _41755_);
  and _63307_ (_11862_, _04794_, _04547_);
  nor _63308_ (_11863_, _11862_, _04796_);
  nor _63309_ (_11864_, _04964_, _04795_);
  nor _63310_ (_11865_, _11864_, _05103_);
  and _63311_ (_11866_, _11865_, _11863_);
  and _63312_ (_11867_, _11866_, _04794_);
  not _63313_ (_11868_, _11867_);
  nand _63314_ (_11869_, _03160_, _02887_);
  and _63315_ (_11870_, _05941_, _03321_);
  nand _63316_ (_11871_, _11870_, _04518_);
  or _63317_ (_11872_, _06478_, _03401_);
  nand _63318_ (_11873_, _11872_, _08190_);
  and _63319_ (_11874_, _11873_, _04478_);
  nor _63320_ (_11875_, _11647_, _05188_);
  or _63321_ (_11876_, _11875_, _05778_);
  and _63322_ (_11877_, _05833_, _04439_);
  and _63323_ (_11878_, _03923_, \oc8051_golden_model_1.PC [0]);
  nor _63324_ (_11879_, _03923_, _03321_);
  or _63325_ (_11880_, _11879_, _11878_);
  and _63326_ (_11881_, _11880_, _05831_);
  or _63327_ (_11882_, _11881_, _11877_);
  and _63328_ (_11883_, _11882_, _04866_);
  and _63329_ (_11884_, _05941_, _04445_);
  or _63330_ (_11885_, _11884_, _11883_);
  and _63331_ (_11886_, _11885_, _05820_);
  nand _63332_ (_11887_, _11647_, _10682_);
  and _63333_ (_11888_, _11887_, _04443_);
  or _63334_ (_11889_, _11888_, _04746_);
  or _63335_ (_11890_, _11889_, _11886_);
  nor _63336_ (_11891_, _03203_, \oc8051_golden_model_1.PC [0]);
  nor _63337_ (_11892_, _11891_, _04454_);
  and _63338_ (_11893_, _11892_, _11890_);
  and _63339_ (_11894_, _04454_, _04419_);
  or _63340_ (_11895_, _11894_, _04462_);
  or _63341_ (_11896_, _11895_, _11893_);
  and _63342_ (_11897_, _11896_, _11876_);
  or _63343_ (_11898_, _11897_, _03511_);
  nand _63344_ (_11899_, _08191_, _03511_);
  and _63345_ (_11900_, _11899_, _03509_);
  and _63346_ (_11901_, _11900_, _11898_);
  nor _63347_ (_11902_, _11648_, _03509_);
  and _63348_ (_11903_, _11902_, _11887_);
  or _63349_ (_11904_, _11903_, _11901_);
  and _63350_ (_11905_, _11904_, _03200_);
  or _63351_ (_11906_, _03200_, _02887_);
  nand _63352_ (_11907_, _03602_, _11906_);
  or _63353_ (_11908_, _11907_, _11905_);
  nand _63354_ (_11909_, _08191_, _04053_);
  and _63355_ (_11910_, _11909_, _05857_);
  and _63356_ (_11911_, _11910_, _11908_);
  or _63357_ (_11912_, _11911_, _11874_);
  and _63358_ (_11913_, _11912_, _04901_);
  nor _63359_ (_11914_, _10707_, _05188_);
  and _63360_ (_11915_, _05188_, \oc8051_golden_model_1.PSW [7]);
  nor _63361_ (_11916_, _11915_, _11914_);
  nor _63362_ (_11917_, _11916_, _04901_);
  or _63363_ (_11918_, _11917_, _03223_);
  or _63364_ (_11919_, _11918_, _11913_);
  and _63365_ (_11920_, _03223_, _02887_);
  nor _63366_ (_11921_, _11920_, _06040_);
  and _63367_ (_11922_, _11921_, _11919_);
  and _63368_ (_11923_, _06040_, _04419_);
  or _63369_ (_11924_, _11923_, _06045_);
  or _63370_ (_11925_, _11924_, _11922_);
  or _63371_ (_11926_, _06715_, _06051_);
  and _63372_ (_11927_, _11926_, _06050_);
  and _63373_ (_11928_, _11927_, _11925_);
  and _63374_ (_11929_, _06086_, _04419_);
  and _63375_ (_11930_, _06269_, \oc8051_golden_model_1.IP [0]);
  and _63376_ (_11931_, _06273_, \oc8051_golden_model_1.B [0]);
  nor _63377_ (_11932_, _11931_, _11930_);
  and _63378_ (_11933_, _06276_, \oc8051_golden_model_1.PSW [0]);
  and _63379_ (_11934_, _06278_, \oc8051_golden_model_1.ACC [0]);
  nor _63380_ (_11935_, _11934_, _11933_);
  and _63381_ (_11936_, _11935_, _11932_);
  and _63382_ (_11937_, _06200_, \oc8051_golden_model_1.DPH [0]);
  and _63383_ (_11938_, _06206_, \oc8051_golden_model_1.TH1 [0]);
  nor _63384_ (_11939_, _11938_, _11937_);
  and _63385_ (_11940_, _06285_, \oc8051_golden_model_1.DPL [0]);
  and _63386_ (_11941_, _06225_, \oc8051_golden_model_1.TL0 [0]);
  nor _63387_ (_11942_, _11941_, _11940_);
  and _63388_ (_11943_, _11942_, _11939_);
  and _63389_ (_11944_, _11943_, _11936_);
  and _63390_ (_11945_, _06256_, \oc8051_golden_model_1.TH0 [0]);
  and _63391_ (_11946_, _06258_, \oc8051_golden_model_1.TL1 [0]);
  nor _63392_ (_11947_, _11946_, _11945_);
  and _63393_ (_11948_, _06263_, \oc8051_golden_model_1.PCON [0]);
  and _63394_ (_11949_, _06265_, \oc8051_golden_model_1.TCON [0]);
  nor _63395_ (_11950_, _11949_, _11948_);
  and _63396_ (_11951_, _11950_, _11947_);
  and _63397_ (_11952_, _06220_, \oc8051_golden_model_1.TMOD [0]);
  not _63398_ (_11953_, _11952_);
  and _63399_ (_11954_, _06245_, \oc8051_golden_model_1.P1INREG [0]);
  and _63400_ (_11955_, _06249_, \oc8051_golden_model_1.P3INREG [0]);
  nor _63401_ (_11956_, _11955_, _11954_);
  and _63402_ (_11957_, _11956_, _11953_);
  and _63403_ (_11958_, _06242_, \oc8051_golden_model_1.P0INREG [0]);
  and _63404_ (_11959_, _06214_, \oc8051_golden_model_1.P2INREG [0]);
  nor _63405_ (_11960_, _11959_, _11958_);
  and _63406_ (_11961_, _11960_, _11957_);
  and _63407_ (_11962_, _06283_, \oc8051_golden_model_1.SP [0]);
  not _63408_ (_11963_, _11962_);
  and _63409_ (_11964_, _06230_, \oc8051_golden_model_1.IE [0]);
  not _63410_ (_11965_, _11964_);
  and _63411_ (_11966_, _06236_, \oc8051_golden_model_1.SCON [0]);
  and _63412_ (_11967_, _06238_, \oc8051_golden_model_1.SBUF [0]);
  nor _63413_ (_11968_, _11967_, _11966_);
  and _63414_ (_11969_, _11968_, _11965_);
  and _63415_ (_11970_, _11969_, _11963_);
  and _63416_ (_11971_, _11970_, _11961_);
  and _63417_ (_11972_, _11971_, _11951_);
  and _63418_ (_11973_, _11972_, _11944_);
  not _63419_ (_11974_, _11973_);
  nor _63420_ (_11975_, _11974_, _11929_);
  nor _63421_ (_11976_, _11975_, _06050_);
  or _63422_ (_11977_, _11976_, _06055_);
  or _63423_ (_11978_, _11977_, _11928_);
  and _63424_ (_11979_, _06055_, _03471_);
  nor _63425_ (_11980_, _11979_, _03439_);
  and _63426_ (_11981_, _11980_, _11978_);
  and _63427_ (_11982_, _06202_, _03439_);
  or _63428_ (_11983_, _11982_, _03189_);
  or _63429_ (_11984_, _11983_, _11981_);
  and _63430_ (_11985_, _03189_, _02887_);
  nor _63431_ (_11986_, _11985_, _04500_);
  and _63432_ (_11987_, _11986_, _11984_);
  and _63433_ (_11988_, _05941_, _04109_);
  and _63434_ (_11989_, _05617_, _06202_);
  nor _63435_ (_11990_, _11989_, _11988_);
  nor _63436_ (_11991_, _11990_, _04502_);
  nor _63437_ (_11992_, _11991_, _04503_);
  or _63438_ (_11993_, _11992_, _11987_);
  and _63439_ (_11994_, _05617_, \oc8051_golden_model_1.ACC [0]);
  nor _63440_ (_11995_, _11994_, _11870_);
  or _63441_ (_11996_, _11995_, _05772_);
  and _63442_ (_11997_, _11996_, _04507_);
  and _63443_ (_11998_, _11997_, _11993_);
  and _63444_ (_11999_, _11989_, _05770_);
  or _63445_ (_12000_, _11999_, _11998_);
  and _63446_ (_12001_, _12000_, _04498_);
  and _63447_ (_12002_, _11994_, _04497_);
  or _63448_ (_12003_, _12002_, _03192_);
  or _63449_ (_12004_, _12003_, _12001_);
  and _63450_ (_12005_, _03192_, _02887_);
  nor _63451_ (_12006_, _12005_, _04516_);
  and _63452_ (_12007_, _12006_, _12004_);
  and _63453_ (_12008_, _11988_, _06324_);
  nor _63454_ (_12009_, _12008_, _04519_);
  or _63455_ (_12010_, _12009_, _12007_);
  and _63456_ (_12011_, _12010_, _11871_);
  or _63457_ (_12012_, _12011_, _03179_);
  not _63458_ (_12013_, _10820_);
  nand _63459_ (_12014_, _03179_, _02887_);
  and _63460_ (_12015_, _12014_, _12013_);
  and _63461_ (_12016_, _12015_, _12012_);
  nor _63462_ (_12017_, _12013_, _04419_);
  or _63463_ (_12018_, _12017_, _04527_);
  or _63464_ (_12019_, _12018_, _12016_);
  or _63465_ (_12020_, _06478_, _06343_);
  and _63466_ (_12021_, _12020_, _12019_);
  or _63467_ (_12022_, _12021_, _04526_);
  or _63468_ (_12023_, _05941_, _06342_);
  and _63469_ (_12024_, _12023_, _10832_);
  and _63470_ (_12025_, _12024_, _12022_);
  and _63471_ (_12026_, _03641_, _02887_);
  or _63472_ (_12027_, _12026_, _03160_);
  or _63473_ (_12028_, _12027_, _12025_);
  and _63474_ (_12029_, _12028_, _11869_);
  or _63475_ (_12030_, _12029_, _03435_);
  or _63476_ (_12031_, _11914_, _03436_);
  and _63477_ (_12032_, _12031_, _10843_);
  and _63478_ (_12033_, _12032_, _12030_);
  not _63479_ (_12034_, _10843_);
  and _63480_ (_12035_, _12034_, _04439_);
  or _63481_ (_12036_, _12035_, _12033_);
  and _63482_ (_12037_, _12036_, _06712_);
  and _63483_ (_12038_, _06478_, _04540_);
  or _63484_ (_12039_, _12038_, _04544_);
  or _63485_ (_12040_, _12039_, _12037_);
  or _63486_ (_12041_, _05941_, _06711_);
  and _63487_ (_12042_, _12041_, _04794_);
  and _63488_ (_12043_, _12042_, _12040_);
  or _63489_ (_12044_, _12043_, _11868_);
  or _63490_ (_12045_, _11867_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _63491_ (_12046_, _05110_, _05113_);
  and _63492_ (_12047_, _12046_, _05117_);
  and _63493_ (_12048_, _12047_, _04551_);
  not _63494_ (_12049_, _12048_);
  and _63495_ (_12050_, _12049_, _12045_);
  and _63496_ (_12051_, _12050_, _12044_);
  not _63497_ (_12052_, _10047_);
  nor _63498_ (_12053_, _12052_, _03641_);
  and _63499_ (_12054_, _10216_, _03641_);
  or _63500_ (_12055_, _12054_, _12053_);
  and _63501_ (_12056_, _12055_, _12048_);
  or _63502_ (_40560_, _12056_, _12051_);
  nor _63503_ (_12057_, _06716_, _06479_);
  or _63504_ (_12058_, _12057_, _06712_);
  or _63505_ (_12059_, _06716_, _06479_);
  and _63506_ (_12060_, _12059_, _04527_);
  not _63507_ (_12061_, _03010_);
  nor _63508_ (_12062_, _03665_, _12061_);
  or _63509_ (_12063_, _04707_, _04187_);
  not _63510_ (_12064_, _12063_);
  nor _63511_ (_12065_, _06692_, _05823_);
  nor _63512_ (_12066_, _12065_, _12064_);
  or _63513_ (_12067_, _12066_, _12062_);
  nand _63514_ (_12068_, _04603_, _06040_);
  nor _63515_ (_12069_, _11621_, _05179_);
  or _63516_ (_12070_, _12069_, _05778_);
  nand _63517_ (_12071_, _12065_, _05833_);
  nor _63518_ (_12072_, _03923_, _03233_);
  and _63519_ (_12073_, _03923_, _02860_);
  or _63520_ (_12074_, _12073_, _12072_);
  or _63521_ (_12075_, _12074_, _03979_);
  or _63522_ (_12076_, _12075_, _04979_);
  and _63523_ (_12077_, _12076_, _12071_);
  and _63524_ (_12078_, _12077_, _04866_);
  or _63525_ (_12079_, _05942_, _05618_);
  and _63526_ (_12080_, _12079_, _04445_);
  or _63527_ (_12081_, _12080_, _12078_);
  or _63528_ (_12082_, _12081_, _04443_);
  nand _63529_ (_12083_, _11621_, _10629_);
  or _63530_ (_12084_, _12083_, _05820_);
  and _63531_ (_12085_, _12084_, _12082_);
  or _63532_ (_12086_, _12085_, _04746_);
  nor _63533_ (_12087_, _03203_, _02860_);
  nor _63534_ (_12088_, _12087_, _04454_);
  and _63535_ (_12089_, _12088_, _12086_);
  and _63536_ (_12090_, _07880_, _04454_);
  or _63537_ (_12091_, _12090_, _04462_);
  or _63538_ (_12092_, _12091_, _12089_);
  and _63539_ (_12093_, _12092_, _12070_);
  or _63540_ (_12094_, _12093_, _03511_);
  nand _63541_ (_12095_, _08177_, _03511_);
  and _63542_ (_12096_, _12095_, _03509_);
  and _63543_ (_12097_, _12096_, _12094_);
  not _63544_ (_12098_, _11622_);
  and _63545_ (_12099_, _12083_, _12098_);
  and _63546_ (_12100_, _12099_, _03508_);
  or _63547_ (_12101_, _12100_, _12097_);
  and _63548_ (_12102_, _12101_, _03200_);
  or _63549_ (_12103_, _03200_, \oc8051_golden_model_1.PC [1]);
  nand _63550_ (_12104_, _03602_, _12103_);
  or _63551_ (_12105_, _12104_, _12102_);
  nand _63552_ (_12106_, _08177_, _04053_);
  and _63553_ (_12107_, _12106_, _05857_);
  and _63554_ (_12108_, _12107_, _12105_);
  or _63555_ (_12109_, _06433_, _03401_);
  nand _63556_ (_12110_, _12109_, _08176_);
  and _63557_ (_12111_, _12110_, _04478_);
  or _63558_ (_12112_, _12111_, _04476_);
  or _63559_ (_12113_, _12112_, _12108_);
  nor _63560_ (_12114_, _10651_, _05179_);
  and _63561_ (_12115_, _05179_, \oc8051_golden_model_1.PSW [7]);
  nor _63562_ (_12116_, _12115_, _12114_);
  nand _63563_ (_12117_, _12116_, _04476_);
  and _63564_ (_12118_, _12117_, _04853_);
  and _63565_ (_12119_, _12118_, _12113_);
  and _63566_ (_12120_, _03223_, _02860_);
  or _63567_ (_12121_, _06040_, _12120_);
  or _63568_ (_12122_, _12121_, _12119_);
  and _63569_ (_12123_, _12122_, _12068_);
  or _63570_ (_12124_, _12123_, _06045_);
  or _63571_ (_12125_, _06714_, _06051_);
  and _63572_ (_12126_, _12125_, _06050_);
  and _63573_ (_12127_, _12126_, _12124_);
  nor _63574_ (_12128_, _06087_, _04603_);
  and _63575_ (_12129_, _06283_, \oc8051_golden_model_1.SP [1]);
  not _63576_ (_12130_, _12129_);
  and _63577_ (_12131_, _06285_, \oc8051_golden_model_1.DPL [1]);
  not _63578_ (_12132_, _12131_);
  and _63579_ (_12133_, _06230_, \oc8051_golden_model_1.IE [1]);
  not _63580_ (_12134_, _12133_);
  and _63581_ (_12135_, _06236_, \oc8051_golden_model_1.SCON [1]);
  and _63582_ (_12136_, _06238_, \oc8051_golden_model_1.SBUF [1]);
  nor _63583_ (_12137_, _12136_, _12135_);
  and _63584_ (_12138_, _12137_, _12134_);
  and _63585_ (_12139_, _12138_, _12132_);
  and _63586_ (_12140_, _12139_, _12130_);
  and _63587_ (_12141_, _06269_, \oc8051_golden_model_1.IP [1]);
  and _63588_ (_12142_, _06278_, \oc8051_golden_model_1.ACC [1]);
  nor _63589_ (_12143_, _12142_, _12141_);
  and _63590_ (_12144_, _06276_, \oc8051_golden_model_1.PSW [1]);
  and _63591_ (_12145_, _06273_, \oc8051_golden_model_1.B [1]);
  nor _63592_ (_12146_, _12145_, _12144_);
  and _63593_ (_12147_, _12146_, _12143_);
  and _63594_ (_12148_, _06214_, \oc8051_golden_model_1.P2INREG [1]);
  not _63595_ (_12149_, _12148_);
  and _63596_ (_12150_, _06245_, \oc8051_golden_model_1.P1INREG [1]);
  and _63597_ (_12151_, _06249_, \oc8051_golden_model_1.P3INREG [1]);
  nor _63598_ (_12152_, _12151_, _12150_);
  and _63599_ (_12153_, _12152_, _12149_);
  and _63600_ (_12154_, _06242_, \oc8051_golden_model_1.P0INREG [1]);
  and _63601_ (_12155_, _06220_, \oc8051_golden_model_1.TMOD [1]);
  nor _63602_ (_12156_, _12155_, _12154_);
  and _63603_ (_12157_, _12156_, _12153_);
  and _63604_ (_12158_, _12157_, _12147_);
  and _63605_ (_12159_, _12158_, _12140_);
  and _63606_ (_12160_, _06256_, \oc8051_golden_model_1.TH0 [1]);
  and _63607_ (_12161_, _06258_, \oc8051_golden_model_1.TL1 [1]);
  nor _63608_ (_12162_, _12161_, _12160_);
  and _63609_ (_12163_, _06263_, \oc8051_golden_model_1.PCON [1]);
  and _63610_ (_12164_, _06265_, \oc8051_golden_model_1.TCON [1]);
  nor _63611_ (_12165_, _12164_, _12163_);
  and _63612_ (_12166_, _12165_, _12162_);
  and _63613_ (_12167_, _06200_, \oc8051_golden_model_1.DPH [1]);
  not _63614_ (_12168_, _12167_);
  and _63615_ (_12169_, _06225_, \oc8051_golden_model_1.TL0 [1]);
  and _63616_ (_12170_, _06206_, \oc8051_golden_model_1.TH1 [1]);
  nor _63617_ (_12171_, _12170_, _12169_);
  and _63618_ (_12172_, _12171_, _12168_);
  and _63619_ (_12173_, _12172_, _12166_);
  and _63620_ (_12174_, _12173_, _12159_);
  not _63621_ (_12175_, _12174_);
  nor _63622_ (_12176_, _12175_, _12128_);
  nor _63623_ (_12177_, _12176_, _06050_);
  or _63624_ (_12178_, _12177_, _06055_);
  or _63625_ (_12179_, _12178_, _12127_);
  and _63626_ (_12180_, _06055_, _04284_);
  nor _63627_ (_12181_, _12180_, _03439_);
  and _63628_ (_12182_, _12181_, _12179_);
  and _63629_ (_12183_, _06222_, _03439_);
  or _63630_ (_12184_, _12183_, _03189_);
  or _63631_ (_12185_, _12184_, _12182_);
  and _63632_ (_12186_, _03189_, \oc8051_golden_model_1.PC [1]);
  nor _63633_ (_12187_, _12186_, _04500_);
  and _63634_ (_12188_, _12187_, _12185_);
  and _63635_ (_12189_, _05940_, _04317_);
  and _63636_ (_12190_, _05569_, _06222_);
  nor _63637_ (_12191_, _12190_, _12189_);
  nor _63638_ (_12192_, _12191_, _04502_);
  nor _63639_ (_12193_, _12192_, _04503_);
  or _63640_ (_12194_, _12193_, _12188_);
  and _63641_ (_12195_, _05569_, \oc8051_golden_model_1.ACC [1]);
  and _63642_ (_12196_, _05940_, _03233_);
  nor _63643_ (_12197_, _12196_, _12195_);
  or _63644_ (_12198_, _12197_, _05772_);
  and _63645_ (_12199_, _12198_, _04507_);
  and _63646_ (_12200_, _12199_, _12194_);
  and _63647_ (_12201_, _12190_, _05770_);
  or _63648_ (_12202_, _12201_, _12200_);
  and _63649_ (_12203_, _12202_, _04498_);
  and _63650_ (_12204_, _12195_, _04497_);
  or _63651_ (_12205_, _12204_, _03192_);
  or _63652_ (_12206_, _12205_, _12203_);
  and _63653_ (_12207_, _03192_, \oc8051_golden_model_1.PC [1]);
  nor _63654_ (_12208_, _12207_, _04516_);
  and _63655_ (_12209_, _12208_, _12206_);
  and _63656_ (_12210_, _12189_, _06324_);
  nor _63657_ (_12211_, _12210_, _04519_);
  or _63658_ (_12212_, _12211_, _12209_);
  nand _63659_ (_12213_, _12196_, _04518_);
  and _63660_ (_12214_, _12213_, _06328_);
  and _63661_ (_12215_, _12214_, _12212_);
  and _63662_ (_12216_, _03179_, _02860_);
  or _63663_ (_12217_, _04705_, _12216_);
  or _63664_ (_12218_, _12217_, _12215_);
  nand _63665_ (_12219_, _12065_, _04705_);
  and _63666_ (_12220_, _12219_, _12064_);
  and _63667_ (_12221_, _12220_, _12218_);
  or _63668_ (_12222_, _12221_, _12067_);
  nor _63669_ (_12223_, _04681_, _04188_);
  nor _63670_ (_12224_, _12065_, _04194_);
  or _63671_ (_12225_, _12224_, _12223_);
  and _63672_ (_12226_, _12225_, _12222_);
  not _63673_ (_12227_, _04194_);
  nor _63674_ (_12228_, _12065_, _12227_);
  or _63675_ (_12229_, _12228_, _12226_);
  and _63676_ (_12230_, _12229_, _06343_);
  or _63677_ (_12231_, _12230_, _12060_);
  and _63678_ (_12232_, _12231_, _06342_);
  and _63679_ (_12233_, _12079_, _04526_);
  or _63680_ (_12234_, _12233_, _03641_);
  or _63681_ (_12235_, _12234_, _12232_);
  nand _63682_ (_12236_, _03641_, _10190_);
  and _63683_ (_12237_, _12236_, _03161_);
  and _63684_ (_12238_, _12237_, _12235_);
  and _63685_ (_12239_, _03160_, _02860_);
  or _63686_ (_12240_, _03435_, _12239_);
  or _63687_ (_12241_, _12240_, _12238_);
  or _63688_ (_12242_, _12114_, _03436_);
  and _63689_ (_12243_, _12242_, _10843_);
  and _63690_ (_12244_, _12243_, _12241_);
  and _63691_ (_12245_, _12065_, _12034_);
  or _63692_ (_12246_, _12245_, _04540_);
  or _63693_ (_12247_, _12246_, _12244_);
  and _63694_ (_12248_, _12247_, _12058_);
  or _63695_ (_12249_, _12248_, _04544_);
  or _63696_ (_12250_, _05941_, _05940_);
  or _63697_ (_12251_, _05617_, _05569_);
  and _63698_ (_12252_, _12251_, _12250_);
  or _63699_ (_12253_, _12252_, _06711_);
  and _63700_ (_12254_, _12253_, _04794_);
  and _63701_ (_12255_, _12254_, _12249_);
  or _63702_ (_12256_, _12255_, _11868_);
  or _63703_ (_12257_, _11867_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _63704_ (_12258_, _12257_, _12049_);
  and _63705_ (_12259_, _12258_, _12256_);
  not _63706_ (_12260_, _09995_);
  nor _63707_ (_12261_, _12260_, _03641_);
  and _63708_ (_12262_, _10156_, _03641_);
  or _63709_ (_12263_, _12262_, _12261_);
  and _63710_ (_12264_, _12263_, _12048_);
  or _63711_ (_40562_, _12264_, _12259_);
  not _63712_ (_12265_, _04212_);
  nor _63713_ (_12266_, _06716_, _06718_);
  nor _63714_ (_12267_, _12266_, _08068_);
  or _63715_ (_12268_, _12267_, _12265_);
  nor _63716_ (_12269_, _10627_, _05271_);
  or _63717_ (_12270_, _12269_, _03436_);
  nor _63718_ (_12271_, _05664_, _03920_);
  and _63719_ (_12272_, _05664_, _03920_);
  nor _63720_ (_12273_, _12272_, _12271_);
  and _63721_ (_12274_, _12273_, _04500_);
  nand _63722_ (_12275_, _05026_, _06040_);
  nor _63723_ (_12276_, _11609_, _05271_);
  or _63724_ (_12277_, _12276_, _05778_);
  nand _63725_ (_12278_, _11609_, _10604_);
  or _63726_ (_12279_, _12278_, _05820_);
  or _63727_ (_12280_, _12251_, _05665_);
  or _63728_ (_12281_, _05942_, _05664_);
  and _63729_ (_12282_, _12281_, _12280_);
  nor _63730_ (_12283_, _12282_, _04866_);
  and _63731_ (_12284_, _05823_, _05026_);
  nor _63732_ (_12285_, _05823_, _05026_);
  or _63733_ (_12286_, _12285_, _12284_);
  or _63734_ (_12287_, _12286_, _05831_);
  and _63735_ (_12288_, _03923_, _03155_);
  nor _63736_ (_12289_, _03923_, _07506_);
  or _63737_ (_12290_, _12289_, _12288_);
  nor _63738_ (_12291_, _12290_, _05833_);
  nor _63739_ (_12292_, _12291_, _04445_);
  and _63740_ (_12293_, _12292_, _12287_);
  or _63741_ (_12294_, _12293_, _04443_);
  or _63742_ (_12295_, _12294_, _12283_);
  and _63743_ (_12296_, _12295_, _12279_);
  or _63744_ (_12297_, _12296_, _04746_);
  nor _63745_ (_12298_, _03203_, _03155_);
  nor _63746_ (_12299_, _12298_, _04454_);
  and _63747_ (_12300_, _12299_, _12297_);
  and _63748_ (_12301_, _07865_, _04454_);
  or _63749_ (_12302_, _12301_, _04462_);
  or _63750_ (_12303_, _12302_, _12300_);
  and _63751_ (_12304_, _12303_, _12277_);
  or _63752_ (_12305_, _12304_, _03511_);
  nand _63753_ (_12306_, _08163_, _03511_);
  and _63754_ (_12307_, _12306_, _03509_);
  and _63755_ (_12308_, _12307_, _12305_);
  not _63756_ (_12309_, _11610_);
  and _63757_ (_12310_, _12278_, _12309_);
  and _63758_ (_12311_, _12310_, _03508_);
  or _63759_ (_12312_, _12311_, _12308_);
  and _63760_ (_12313_, _12312_, _03200_);
  or _63761_ (_12314_, _03200_, _03626_);
  nand _63762_ (_12315_, _03602_, _12314_);
  or _63763_ (_12316_, _12315_, _12313_);
  nand _63764_ (_12317_, _08163_, _04053_);
  and _63765_ (_12318_, _12317_, _12316_);
  or _63766_ (_12319_, _12318_, _04478_);
  and _63767_ (_12320_, _06718_, _05215_);
  nand _63768_ (_12321_, _08162_, _04478_);
  or _63769_ (_12322_, _12321_, _12320_);
  and _63770_ (_12323_, _12322_, _12319_);
  or _63771_ (_12324_, _12323_, _04476_);
  and _63772_ (_12325_, _05271_, \oc8051_golden_model_1.PSW [7]);
  nor _63773_ (_12326_, _12325_, _12269_);
  nand _63774_ (_12327_, _12326_, _04476_);
  and _63775_ (_12328_, _12327_, _04853_);
  and _63776_ (_12329_, _12328_, _12324_);
  and _63777_ (_12330_, _03223_, _03155_);
  or _63778_ (_12331_, _06040_, _12330_);
  or _63779_ (_12332_, _12331_, _12329_);
  and _63780_ (_12333_, _12332_, _12275_);
  or _63781_ (_12334_, _12333_, _06045_);
  or _63782_ (_12335_, _06718_, _06051_);
  and _63783_ (_12336_, _12335_, _06050_);
  and _63784_ (_12337_, _12336_, _12334_);
  nor _63785_ (_12338_, _06087_, _05026_);
  and _63786_ (_12339_, _06200_, \oc8051_golden_model_1.DPH [2]);
  and _63787_ (_12340_, _06206_, \oc8051_golden_model_1.TH1 [2]);
  nor _63788_ (_12341_, _12340_, _12339_);
  and _63789_ (_12342_, _06214_, \oc8051_golden_model_1.P2INREG [2]);
  not _63790_ (_12343_, _12342_);
  and _63791_ (_12344_, _06220_, \oc8051_golden_model_1.TMOD [2]);
  and _63792_ (_12345_, _06225_, \oc8051_golden_model_1.TL0 [2]);
  nor _63793_ (_12346_, _12345_, _12344_);
  and _63794_ (_12347_, _12346_, _12343_);
  and _63795_ (_12348_, _06230_, \oc8051_golden_model_1.IE [2]);
  not _63796_ (_12349_, _12348_);
  and _63797_ (_12350_, _06236_, \oc8051_golden_model_1.SCON [2]);
  and _63798_ (_12351_, _06238_, \oc8051_golden_model_1.SBUF [2]);
  nor _63799_ (_12352_, _12351_, _12350_);
  and _63800_ (_12353_, _12352_, _12349_);
  and _63801_ (_12354_, _06242_, \oc8051_golden_model_1.P0INREG [2]);
  not _63802_ (_12355_, _12354_);
  and _63803_ (_12356_, _06245_, \oc8051_golden_model_1.P1INREG [2]);
  and _63804_ (_12357_, _06249_, \oc8051_golden_model_1.P3INREG [2]);
  nor _63805_ (_12358_, _12357_, _12356_);
  and _63806_ (_12359_, _12358_, _12355_);
  and _63807_ (_12360_, _12359_, _12353_);
  and _63808_ (_12361_, _12360_, _12347_);
  and _63809_ (_12362_, _12361_, _12341_);
  and _63810_ (_12363_, _06256_, \oc8051_golden_model_1.TH0 [2]);
  and _63811_ (_12364_, _06258_, \oc8051_golden_model_1.TL1 [2]);
  nor _63812_ (_12365_, _12364_, _12363_);
  and _63813_ (_12366_, _06263_, \oc8051_golden_model_1.PCON [2]);
  and _63814_ (_12367_, _06265_, \oc8051_golden_model_1.TCON [2]);
  nor _63815_ (_12368_, _12367_, _12366_);
  and _63816_ (_12369_, _12368_, _12365_);
  and _63817_ (_12370_, _06269_, \oc8051_golden_model_1.IP [2]);
  and _63818_ (_12371_, _06273_, \oc8051_golden_model_1.B [2]);
  nor _63819_ (_12372_, _12371_, _12370_);
  and _63820_ (_12373_, _06276_, \oc8051_golden_model_1.PSW [2]);
  and _63821_ (_12374_, _06278_, \oc8051_golden_model_1.ACC [2]);
  nor _63822_ (_12375_, _12374_, _12373_);
  and _63823_ (_12376_, _12375_, _12372_);
  and _63824_ (_12377_, _06283_, \oc8051_golden_model_1.SP [2]);
  and _63825_ (_12378_, _06285_, \oc8051_golden_model_1.DPL [2]);
  nor _63826_ (_12379_, _12378_, _12377_);
  and _63827_ (_12380_, _12379_, _12376_);
  and _63828_ (_12381_, _12380_, _12369_);
  and _63829_ (_12382_, _12381_, _12362_);
  not _63830_ (_12383_, _12382_);
  nor _63831_ (_12384_, _12383_, _12338_);
  nor _63832_ (_12385_, _12384_, _06050_);
  or _63833_ (_12386_, _12385_, _06055_);
  or _63834_ (_12387_, _12386_, _12337_);
  and _63835_ (_12388_, _06055_, _03877_);
  nor _63836_ (_12389_, _12388_, _03439_);
  and _63837_ (_12390_, _12389_, _12387_);
  and _63838_ (_12391_, _06261_, _03439_);
  or _63839_ (_12392_, _12391_, _03189_);
  or _63840_ (_12393_, _12392_, _12390_);
  and _63841_ (_12394_, _03189_, _03626_);
  nor _63842_ (_12395_, _12394_, _04500_);
  and _63843_ (_12396_, _12395_, _12393_);
  or _63844_ (_12397_, _12396_, _12274_);
  and _63845_ (_12398_, _12397_, _05772_);
  nor _63846_ (_12399_, _05664_, _07506_);
  and _63847_ (_12400_, _05664_, _07506_);
  nor _63848_ (_12401_, _12400_, _12399_);
  and _63849_ (_12402_, _12401_, _04502_);
  or _63850_ (_12403_, _12402_, _04506_);
  or _63851_ (_12404_, _12403_, _12398_);
  or _63852_ (_12405_, _12271_, _04507_);
  and _63853_ (_12406_, _12405_, _04498_);
  and _63854_ (_12407_, _12406_, _12404_);
  and _63855_ (_12408_, _12399_, _04497_);
  or _63856_ (_12409_, _12408_, _03192_);
  or _63857_ (_12410_, _12409_, _12407_);
  and _63858_ (_12411_, _03192_, _03626_);
  nor _63859_ (_12412_, _12411_, _04516_);
  and _63860_ (_12413_, _12412_, _12410_);
  and _63861_ (_12414_, _12272_, _06324_);
  nor _63862_ (_12415_, _12414_, _04519_);
  or _63863_ (_12416_, _12415_, _12413_);
  nand _63864_ (_12417_, _12400_, _04518_);
  and _63865_ (_12418_, _12417_, _06328_);
  and _63866_ (_12419_, _12418_, _12416_);
  and _63867_ (_12420_, _03179_, _03155_);
  or _63868_ (_12421_, _10820_, _12420_);
  or _63869_ (_12422_, _12421_, _12419_);
  or _63870_ (_12423_, _12286_, _12013_);
  and _63871_ (_12424_, _12423_, _06343_);
  and _63872_ (_12425_, _12424_, _12422_);
  and _63873_ (_12426_, _06479_, _06569_);
  nor _63874_ (_12427_, _06479_, _06569_);
  or _63875_ (_12428_, _12427_, _12426_);
  and _63876_ (_12429_, _12428_, _04527_);
  or _63877_ (_12430_, _12429_, _12425_);
  and _63878_ (_12431_, _12430_, _06342_);
  nor _63879_ (_12432_, _12282_, _06342_);
  or _63880_ (_12433_, _12432_, _03641_);
  or _63881_ (_12434_, _12433_, _12431_);
  nand _63882_ (_12435_, _10188_, _03641_);
  and _63883_ (_12436_, _12435_, _03161_);
  and _63884_ (_12437_, _12436_, _12434_);
  and _63885_ (_12438_, _03160_, _03155_);
  or _63886_ (_12439_, _03435_, _12438_);
  or _63887_ (_12440_, _12439_, _12437_);
  and _63888_ (_12441_, _12440_, _12270_);
  or _63889_ (_12442_, _12441_, _12034_);
  and _63890_ (_12443_, _11572_, _03165_);
  not _63891_ (_12444_, _12443_);
  nor _63892_ (_12445_, _06692_, _07865_);
  nor _63893_ (_12446_, _12445_, _07866_);
  or _63894_ (_12447_, _12446_, _10843_);
  and _63895_ (_12448_, _12447_, _12444_);
  and _63896_ (_12449_, _12448_, _12442_);
  or _63897_ (_12450_, _12267_, _04212_);
  and _63898_ (_12451_, _12450_, _04540_);
  or _63899_ (_12452_, _12451_, _12449_);
  and _63900_ (_12453_, _12452_, _12268_);
  or _63901_ (_12454_, _12453_, _04544_);
  and _63902_ (_12455_, _05664_, _12250_);
  nor _63903_ (_12456_, _12455_, _05666_);
  or _63904_ (_12457_, _12456_, _06711_);
  and _63905_ (_12458_, _12457_, _04794_);
  and _63906_ (_12459_, _12458_, _12454_);
  or _63907_ (_12460_, _12459_, _11868_);
  or _63908_ (_12461_, _11867_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _63909_ (_12462_, _12461_, _12049_);
  and _63910_ (_12463_, _12462_, _12460_);
  not _63911_ (_12464_, _09989_);
  nor _63912_ (_12465_, _12464_, _03641_);
  and _63913_ (_12466_, _10142_, _03641_);
  or _63914_ (_12467_, _12466_, _12465_);
  and _63915_ (_12468_, _12467_, _12048_);
  or _63916_ (_40563_, _12468_, _12463_);
  nor _63917_ (_12469_, _11867_, _04798_);
  nor _63918_ (_12470_, _07866_, _07864_);
  nor _63919_ (_12471_, _12470_, _06694_);
  and _63920_ (_12472_, _12471_, _06712_);
  or _63921_ (_12473_, _12472_, _04721_);
  and _63922_ (_12474_, _03280_, _03179_);
  nand _63923_ (_12475_, _04843_, _06040_);
  nor _63924_ (_12476_, _12284_, _04843_);
  or _63925_ (_12477_, _12476_, _05825_);
  or _63926_ (_12478_, _12477_, _05831_);
  and _63927_ (_12479_, _03923_, _03280_);
  nor _63928_ (_12480_, _03923_, _07500_);
  or _63929_ (_12481_, _12480_, _05833_);
  or _63930_ (_12482_, _12481_, _12479_);
  and _63931_ (_12483_, _12482_, _12478_);
  and _63932_ (_12484_, _12483_, _04866_);
  and _63933_ (_12485_, _12280_, _05521_);
  nor _63934_ (_12486_, _12485_, _05944_);
  nor _63935_ (_12487_, _12486_, _04866_);
  or _63936_ (_12488_, _12487_, _12484_);
  or _63937_ (_12489_, _12488_, _04443_);
  nand _63938_ (_12490_, _11671_, _10739_);
  or _63939_ (_12491_, _12490_, _05820_);
  and _63940_ (_12492_, _12491_, _12489_);
  or _63941_ (_12493_, _12492_, _04746_);
  nor _63942_ (_12494_, _03280_, _03203_);
  nor _63943_ (_12495_, _12494_, _04454_);
  and _63944_ (_12496_, _12495_, _12493_);
  and _63945_ (_12497_, _07864_, _04454_);
  or _63946_ (_12498_, _12497_, _04462_);
  or _63947_ (_12499_, _12498_, _12496_);
  nor _63948_ (_12500_, _11671_, _05265_);
  or _63949_ (_12501_, _12500_, _05778_);
  and _63950_ (_12502_, _12501_, _12499_);
  or _63951_ (_12503_, _12502_, _03511_);
  nand _63952_ (_12504_, _08143_, _03511_);
  and _63953_ (_12505_, _12504_, _03509_);
  and _63954_ (_12506_, _12505_, _12503_);
  not _63955_ (_12507_, _11672_);
  and _63956_ (_12508_, _12490_, _12507_);
  and _63957_ (_12509_, _12508_, _03508_);
  or _63958_ (_12510_, _12509_, _12506_);
  and _63959_ (_12511_, _12510_, _03200_);
  or _63960_ (_12512_, _03675_, _03200_);
  nand _63961_ (_12513_, _03602_, _12512_);
  or _63962_ (_12514_, _12513_, _12511_);
  nand _63963_ (_12515_, _08143_, _04053_);
  and _63964_ (_12516_, _12515_, _12514_);
  or _63965_ (_12517_, _12516_, _04478_);
  and _63966_ (_12518_, _06717_, _05215_);
  nand _63967_ (_12519_, _08142_, _04478_);
  or _63968_ (_12520_, _12519_, _12518_);
  and _63969_ (_12521_, _12520_, _12517_);
  or _63970_ (_12522_, _12521_, _04476_);
  and _63971_ (_12523_, _05265_, \oc8051_golden_model_1.PSW [7]);
  nor _63972_ (_12524_, _10764_, _05265_);
  nor _63973_ (_12525_, _12524_, _12523_);
  nand _63974_ (_12526_, _12525_, _04476_);
  and _63975_ (_12527_, _12526_, _04853_);
  and _63976_ (_12528_, _12527_, _12522_);
  and _63977_ (_12529_, _03280_, _03223_);
  or _63978_ (_12530_, _06040_, _12529_);
  or _63979_ (_12531_, _12530_, _12528_);
  and _63980_ (_12532_, _12531_, _12475_);
  or _63981_ (_12533_, _12532_, _06045_);
  or _63982_ (_12534_, _06717_, _06051_);
  and _63983_ (_12535_, _12534_, _06050_);
  and _63984_ (_12536_, _12535_, _12533_);
  nor _63985_ (_12537_, _06087_, _04843_);
  and _63986_ (_12538_, _06200_, \oc8051_golden_model_1.DPH [3]);
  and _63987_ (_12539_, _06206_, \oc8051_golden_model_1.TH1 [3]);
  nor _63988_ (_12540_, _12539_, _12538_);
  and _63989_ (_12541_, _06214_, \oc8051_golden_model_1.P2INREG [3]);
  not _63990_ (_12542_, _12541_);
  and _63991_ (_12543_, _06220_, \oc8051_golden_model_1.TMOD [3]);
  and _63992_ (_12544_, _06225_, \oc8051_golden_model_1.TL0 [3]);
  nor _63993_ (_12545_, _12544_, _12543_);
  and _63994_ (_12546_, _12545_, _12542_);
  and _63995_ (_12547_, _06230_, \oc8051_golden_model_1.IE [3]);
  not _63996_ (_12548_, _12547_);
  and _63997_ (_12549_, _06236_, \oc8051_golden_model_1.SCON [3]);
  and _63998_ (_12550_, _06238_, \oc8051_golden_model_1.SBUF [3]);
  nor _63999_ (_12551_, _12550_, _12549_);
  and _64000_ (_12552_, _12551_, _12548_);
  and _64001_ (_12553_, _06242_, \oc8051_golden_model_1.P0INREG [3]);
  not _64002_ (_12554_, _12553_);
  and _64003_ (_12555_, _06245_, \oc8051_golden_model_1.P1INREG [3]);
  and _64004_ (_12556_, _06249_, \oc8051_golden_model_1.P3INREG [3]);
  nor _64005_ (_12557_, _12556_, _12555_);
  and _64006_ (_12558_, _12557_, _12554_);
  and _64007_ (_12559_, _12558_, _12552_);
  and _64008_ (_12560_, _12559_, _12546_);
  and _64009_ (_12561_, _12560_, _12540_);
  and _64010_ (_12562_, _06256_, \oc8051_golden_model_1.TH0 [3]);
  and _64011_ (_12563_, _06258_, \oc8051_golden_model_1.TL1 [3]);
  nor _64012_ (_12564_, _12563_, _12562_);
  and _64013_ (_12565_, _06263_, \oc8051_golden_model_1.PCON [3]);
  and _64014_ (_12566_, _06265_, \oc8051_golden_model_1.TCON [3]);
  nor _64015_ (_12567_, _12566_, _12565_);
  and _64016_ (_12568_, _12567_, _12564_);
  and _64017_ (_12569_, _06269_, \oc8051_golden_model_1.IP [3]);
  and _64018_ (_12570_, _06273_, \oc8051_golden_model_1.B [3]);
  nor _64019_ (_12571_, _12570_, _12569_);
  and _64020_ (_12572_, _06276_, \oc8051_golden_model_1.PSW [3]);
  and _64021_ (_12573_, _06278_, \oc8051_golden_model_1.ACC [3]);
  nor _64022_ (_12574_, _12573_, _12572_);
  and _64023_ (_12575_, _12574_, _12571_);
  and _64024_ (_12576_, _06283_, \oc8051_golden_model_1.SP [3]);
  and _64025_ (_12577_, _06285_, \oc8051_golden_model_1.DPL [3]);
  nor _64026_ (_12578_, _12577_, _12576_);
  and _64027_ (_12579_, _12578_, _12575_);
  and _64028_ (_12580_, _12579_, _12568_);
  and _64029_ (_12581_, _12580_, _12561_);
  not _64030_ (_12582_, _12581_);
  nor _64031_ (_12583_, _12582_, _12537_);
  nor _64032_ (_12584_, _12583_, _06050_);
  or _64033_ (_12585_, _12584_, _06055_);
  or _64034_ (_12586_, _12585_, _12536_);
  and _64035_ (_12587_, _06055_, _03432_);
  nor _64036_ (_12588_, _12587_, _03439_);
  and _64037_ (_12589_, _12588_, _12586_);
  and _64038_ (_12590_, _06217_, _03439_);
  or _64039_ (_12591_, _12590_, _03189_);
  or _64040_ (_12592_, _12591_, _12589_);
  and _64041_ (_12593_, _03675_, _03189_);
  nor _64042_ (_12594_, _12593_, _04500_);
  and _64043_ (_12595_, _12594_, _12592_);
  nor _64044_ (_12596_, _05520_, _03742_);
  and _64045_ (_12597_, _05520_, _03742_);
  nor _64046_ (_12598_, _12597_, _12596_);
  and _64047_ (_12599_, _12598_, _04500_);
  or _64048_ (_12600_, _12599_, _12595_);
  and _64049_ (_12601_, _12600_, _05772_);
  nor _64050_ (_12602_, _05520_, _07500_);
  and _64051_ (_12603_, _05520_, _07500_);
  nor _64052_ (_12604_, _12603_, _12602_);
  and _64053_ (_12605_, _12604_, _04502_);
  or _64054_ (_12606_, _12605_, _04506_);
  or _64055_ (_12607_, _12606_, _12601_);
  or _64056_ (_12608_, _12596_, _04507_);
  and _64057_ (_12609_, _12608_, _04498_);
  and _64058_ (_12610_, _12609_, _12607_);
  and _64059_ (_12611_, _12602_, _04497_);
  or _64060_ (_12612_, _12611_, _03192_);
  or _64061_ (_12613_, _12612_, _12610_);
  and _64062_ (_12614_, _03675_, _03192_);
  nor _64063_ (_12615_, _12614_, _04516_);
  and _64064_ (_12616_, _12615_, _12613_);
  and _64065_ (_12617_, _12597_, _06324_);
  nor _64066_ (_12618_, _12617_, _04519_);
  or _64067_ (_12619_, _12618_, _12616_);
  nand _64068_ (_12620_, _12603_, _04518_);
  and _64069_ (_12621_, _12620_, _06328_);
  and _64070_ (_12622_, _12621_, _12619_);
  or _64071_ (_12623_, _12622_, _12474_);
  and _64072_ (_12624_, _12623_, _12013_);
  and _64073_ (_12625_, _12477_, _10820_);
  or _64074_ (_12626_, _12625_, _04527_);
  or _64075_ (_12627_, _12626_, _12624_);
  nor _64076_ (_12628_, _12426_, _06524_);
  or _64077_ (_12629_, _06571_, _06343_);
  or _64078_ (_12630_, _12629_, _12628_);
  and _64079_ (_12631_, _12630_, _06342_);
  and _64080_ (_12632_, _12631_, _12627_);
  nor _64081_ (_12633_, _12486_, _06342_);
  or _64082_ (_12634_, _12633_, _03641_);
  or _64083_ (_12635_, _12634_, _12632_);
  nand _64084_ (_12636_, _10183_, _03641_);
  and _64085_ (_12637_, _12636_, _03161_);
  and _64086_ (_12638_, _12637_, _12635_);
  and _64087_ (_12639_, _03280_, _03160_);
  or _64088_ (_12640_, _03435_, _12639_);
  or _64089_ (_12641_, _12640_, _12638_);
  or _64090_ (_12642_, _12524_, _03436_);
  or _64091_ (_12643_, _04759_, _04205_);
  nor _64092_ (_12644_, _12643_, _04766_);
  and _64093_ (_12645_, _12644_, _12642_);
  and _64094_ (_12646_, _12645_, _12641_);
  not _64095_ (_12647_, _12644_);
  and _64096_ (_12648_, _12647_, _12471_);
  or _64097_ (_12649_, _12648_, _04209_);
  or _64098_ (_12650_, _12649_, _12646_);
  and _64099_ (_12651_, _12650_, _12473_);
  or _64100_ (_12652_, _08068_, _06717_);
  nor _64101_ (_12653_, _06720_, _06712_);
  and _64102_ (_12654_, _12653_, _12652_);
  or _64103_ (_12655_, _12654_, _04544_);
  or _64104_ (_12656_, _12655_, _12651_);
  nor _64105_ (_12657_, _05666_, _05521_);
  nor _64106_ (_12658_, _12657_, _05667_);
  or _64107_ (_12659_, _12658_, _06711_);
  and _64108_ (_12660_, _12659_, _04794_);
  and _64109_ (_12661_, _12660_, _12656_);
  and _64110_ (_12662_, _12661_, _11866_);
  or _64111_ (_12663_, _12662_, _12469_);
  and _64112_ (_12664_, _12663_, _12049_);
  nor _64113_ (_12665_, _05116_, _42967_);
  and _64114_ (_12666_, _12665_, _41755_);
  nor _64115_ (_12667_, _05116_, _03502_);
  and _64116_ (_12668_, _12667_, _42963_);
  and _64117_ (_12669_, _12668_, _41755_);
  nor _64118_ (_12670_, _05116_, \oc8051_golden_model_1.SP [1]);
  and _64119_ (_12671_, _12670_, _42963_);
  and _64120_ (_12672_, _12671_, _41755_);
  nor _64121_ (_12673_, _12672_, _12669_);
  not _64122_ (_12674_, _05110_);
  or _64123_ (_12675_, _05116_, _12674_);
  or _64124_ (_12676_, _12675_, _42967_);
  or _64125_ (_12677_, _12676_, rst);
  not _64126_ (_12678_, _05113_);
  or _64127_ (_12679_, _05116_, _12678_);
  or _64128_ (_12680_, _12679_, _42967_);
  or _64129_ (_12681_, _12680_, rst);
  and _64130_ (_12682_, _12681_, _12677_);
  and _64131_ (_12683_, _12682_, _12673_);
  and _64132_ (_12684_, _12683_, _12666_);
  not _64133_ (_12685_, _05116_);
  and _64134_ (_12686_, _09984_, _10832_);
  and _64135_ (_12687_, _10147_, _03641_);
  or _64136_ (_12688_, _12687_, _12686_);
  and _64137_ (_12689_, _12688_, _12685_);
  and _64138_ (_12690_, _12689_, _42963_);
  and _64139_ (_12691_, _12690_, _41755_);
  and _64140_ (_12692_, _12691_, _12684_);
  or _64141_ (_40565_, _12692_, _12664_);
  nor _64142_ (_12693_, _06720_, _06722_);
  nor _64143_ (_12694_, _12693_, _08046_);
  and _64144_ (_12695_, _12694_, _12443_);
  or _64145_ (_12696_, _06694_, _07848_);
  and _64146_ (_12697_, _06694_, _07848_);
  nor _64147_ (_12698_, _10843_, _12697_);
  and _64148_ (_12699_, _12698_, _12696_);
  and _64149_ (_12700_, _06571_, _06661_);
  nor _64150_ (_12701_, _06571_, _06661_);
  or _64151_ (_12703_, _12701_, _12700_);
  and _64152_ (_12704_, _12703_, _04527_);
  nor _64153_ (_12705_, _05825_, _05712_);
  and _64154_ (_12706_, _05825_, _05712_);
  or _64155_ (_12707_, _12706_, _12705_);
  or _64156_ (_12708_, _12707_, _04709_);
  nor _64157_ (_12709_, _06195_, _05760_);
  and _64158_ (_12710_, _06195_, _05760_);
  nor _64159_ (_12711_, _12710_, _12709_);
  and _64160_ (_12712_, _12711_, _04500_);
  nand _64161_ (_12713_, _05712_, _06040_);
  nor _64162_ (_12714_, _10677_, _10654_);
  and _64163_ (_12715_, _10654_, \oc8051_golden_model_1.PSW [7]);
  nor _64164_ (_12716_, _12715_, _12714_);
  nor _64165_ (_12717_, _12716_, _04901_);
  nor _64166_ (_12718_, _10654_, _11634_);
  or _64167_ (_12719_, _12718_, _05778_);
  or _64168_ (_12720_, _12707_, _05831_);
  and _64169_ (_12721_, _10015_, _03923_);
  nor _64170_ (_12722_, _03923_, _07405_);
  or _64171_ (_12724_, _12722_, _12721_);
  or _64172_ (_12725_, _12724_, _05833_);
  and _64173_ (_12726_, _12725_, _12720_);
  or _64174_ (_12727_, _12726_, _04438_);
  or _64175_ (_12728_, _06722_, _05847_);
  and _64176_ (_12729_, _12728_, _12727_);
  and _64177_ (_12730_, _12729_, _04866_);
  and _64178_ (_12731_, _05944_, _05760_);
  nor _64179_ (_12732_, _05944_, _05760_);
  nor _64180_ (_12733_, _12732_, _12731_);
  nor _64181_ (_12734_, _12733_, _04866_);
  or _64182_ (_12735_, _12734_, _12730_);
  and _64183_ (_12736_, _12735_, _05820_);
  nand _64184_ (_12737_, _10655_, _11634_);
  and _64185_ (_12738_, _12737_, _04443_);
  or _64186_ (_12739_, _12738_, _04746_);
  or _64187_ (_12740_, _12739_, _12736_);
  nor _64188_ (_12741_, _10015_, _03203_);
  nor _64189_ (_12742_, _12741_, _04454_);
  and _64190_ (_12743_, _12742_, _12740_);
  and _64191_ (_12744_, _07848_, _04454_);
  or _64192_ (_12745_, _12744_, _04462_);
  or _64193_ (_12746_, _12745_, _12743_);
  and _64194_ (_12747_, _12746_, _12719_);
  or _64195_ (_12748_, _12747_, _03511_);
  nand _64196_ (_12749_, _08222_, _03511_);
  and _64197_ (_12750_, _12749_, _03509_);
  and _64198_ (_12751_, _12750_, _12748_);
  not _64199_ (_12752_, _11635_);
  and _64200_ (_12753_, _12737_, _12752_);
  and _64201_ (_12754_, _12753_, _03508_);
  or _64202_ (_12755_, _12754_, _12751_);
  and _64203_ (_12756_, _12755_, _03200_);
  or _64204_ (_12757_, _10016_, _03200_);
  nand _64205_ (_12758_, _12757_, _03602_);
  or _64206_ (_12759_, _12758_, _12756_);
  nand _64207_ (_12760_, _08222_, _04053_);
  and _64208_ (_12761_, _12760_, _12759_);
  or _64209_ (_12762_, _12761_, _04478_);
  and _64210_ (_12763_, _06722_, _05215_);
  nand _64211_ (_12764_, _08221_, _04478_);
  or _64212_ (_12765_, _12764_, _12763_);
  and _64213_ (_12766_, _12765_, _04901_);
  and _64214_ (_12767_, _12766_, _12762_);
  or _64215_ (_12768_, _12767_, _12717_);
  and _64216_ (_12769_, _12768_, _04853_);
  and _64217_ (_12770_, _10015_, _03223_);
  or _64218_ (_12771_, _12770_, _06040_);
  or _64219_ (_12772_, _12771_, _12769_);
  and _64220_ (_12773_, _12772_, _12713_);
  or _64221_ (_12774_, _12773_, _06045_);
  or _64222_ (_12775_, _06722_, _06051_);
  and _64223_ (_12776_, _12775_, _06050_);
  and _64224_ (_12777_, _12776_, _12774_);
  nor _64225_ (_12778_, _06087_, _05712_);
  and _64226_ (_12779_, _06283_, \oc8051_golden_model_1.SP [4]);
  not _64227_ (_12780_, _12779_);
  and _64228_ (_12781_, _06230_, \oc8051_golden_model_1.IE [4]);
  not _64229_ (_12782_, _12781_);
  and _64230_ (_12783_, _06236_, \oc8051_golden_model_1.SCON [4]);
  and _64231_ (_12784_, _06238_, \oc8051_golden_model_1.SBUF [4]);
  nor _64232_ (_12785_, _12784_, _12783_);
  and _64233_ (_12786_, _12785_, _12782_);
  and _64234_ (_12787_, _06220_, \oc8051_golden_model_1.TMOD [4]);
  not _64235_ (_12788_, _12787_);
  and _64236_ (_12789_, _06245_, \oc8051_golden_model_1.P1INREG [4]);
  and _64237_ (_12790_, _06249_, \oc8051_golden_model_1.P3INREG [4]);
  nor _64238_ (_12791_, _12790_, _12789_);
  and _64239_ (_12792_, _12791_, _12788_);
  and _64240_ (_12793_, _12792_, _12786_);
  and _64241_ (_12794_, _12793_, _12780_);
  and _64242_ (_12795_, _06200_, \oc8051_golden_model_1.DPH [4]);
  and _64243_ (_12796_, _06206_, \oc8051_golden_model_1.TH1 [4]);
  nor _64244_ (_12797_, _12796_, _12795_);
  and _64245_ (_12798_, _06225_, \oc8051_golden_model_1.TL0 [4]);
  not _64246_ (_12799_, _12798_);
  and _64247_ (_12800_, _06242_, \oc8051_golden_model_1.P0INREG [4]);
  and _64248_ (_12801_, _06214_, \oc8051_golden_model_1.P2INREG [4]);
  nor _64249_ (_12802_, _12801_, _12800_);
  and _64250_ (_12803_, _12802_, _12799_);
  and _64251_ (_12804_, _12803_, _12797_);
  and _64252_ (_12805_, _12804_, _12794_);
  and _64253_ (_12806_, _06285_, \oc8051_golden_model_1.DPL [4]);
  not _64254_ (_12807_, _12806_);
  and _64255_ (_12808_, _06269_, \oc8051_golden_model_1.IP [4]);
  and _64256_ (_12809_, _06273_, \oc8051_golden_model_1.B [4]);
  nor _64257_ (_12810_, _12809_, _12808_);
  and _64258_ (_12811_, _06276_, \oc8051_golden_model_1.PSW [4]);
  and _64259_ (_12812_, _06278_, \oc8051_golden_model_1.ACC [4]);
  nor _64260_ (_12813_, _12812_, _12811_);
  and _64261_ (_12814_, _12813_, _12810_);
  and _64262_ (_12815_, _12814_, _12807_);
  and _64263_ (_12816_, _06229_, _06197_);
  and _64264_ (_12817_, _12816_, \oc8051_golden_model_1.TCON [4]);
  and _64265_ (_12818_, _06256_, \oc8051_golden_model_1.TH0 [4]);
  nor _64266_ (_12819_, _12818_, _12817_);
  and _64267_ (_12820_, _06263_, \oc8051_golden_model_1.PCON [4]);
  and _64268_ (_12821_, _06258_, \oc8051_golden_model_1.TL1 [4]);
  nor _64269_ (_12822_, _12821_, _12820_);
  and _64270_ (_12823_, _12822_, _12819_);
  and _64271_ (_12824_, _12823_, _12815_);
  and _64272_ (_12825_, _12824_, _12805_);
  not _64273_ (_12826_, _12825_);
  nor _64274_ (_12827_, _12826_, _12778_);
  nor _64275_ (_12828_, _12827_, _06050_);
  or _64276_ (_12829_, _12828_, _06055_);
  or _64277_ (_12830_, _12829_, _12777_);
  and _64278_ (_12831_, _06055_, _04249_);
  nor _64279_ (_12832_, _12831_, _03439_);
  and _64280_ (_12833_, _12832_, _12830_);
  and _64281_ (_12834_, _06233_, _03439_);
  or _64282_ (_12835_, _12834_, _03189_);
  or _64283_ (_12836_, _12835_, _12833_);
  and _64284_ (_12837_, _10016_, _03189_);
  nor _64285_ (_12838_, _12837_, _04500_);
  and _64286_ (_12839_, _12838_, _12836_);
  or _64287_ (_12840_, _12839_, _12712_);
  and _64288_ (_12841_, _12840_, _05772_);
  nor _64289_ (_12842_, _05760_, _07405_);
  and _64290_ (_12843_, _05760_, _07405_);
  nor _64291_ (_12844_, _12843_, _12842_);
  and _64292_ (_12845_, _12844_, _04502_);
  or _64293_ (_12846_, _12845_, _12841_);
  and _64294_ (_12847_, _12846_, _05771_);
  and _64295_ (_12848_, _12709_, _04506_);
  or _64296_ (_12849_, _12848_, _04497_);
  or _64297_ (_12850_, _12849_, _12847_);
  or _64298_ (_12851_, _12842_, _04498_);
  and _64299_ (_12852_, _12851_, _12850_);
  or _64300_ (_12853_, _12852_, _03192_);
  and _64301_ (_12854_, _10016_, _03192_);
  nor _64302_ (_12855_, _12854_, _04516_);
  and _64303_ (_12856_, _12855_, _12853_);
  and _64304_ (_12857_, _12710_, _06324_);
  nor _64305_ (_12858_, _12857_, _04519_);
  or _64306_ (_12859_, _12858_, _12856_);
  nand _64307_ (_12860_, _12843_, _04518_);
  and _64308_ (_12861_, _12860_, _06328_);
  and _64309_ (_12862_, _12861_, _12859_);
  nand _64310_ (_12863_, _10015_, _03179_);
  nand _64311_ (_12864_, _12863_, _04709_);
  or _64312_ (_12865_, _12864_, _12862_);
  and _64313_ (_12866_, _12865_, _12708_);
  or _64314_ (_12867_, _12866_, _04681_);
  or _64315_ (_12868_, _12707_, _06335_);
  and _64316_ (_12869_, _12868_, _06343_);
  and _64317_ (_12870_, _12869_, _12867_);
  or _64318_ (_12871_, _12870_, _12704_);
  and _64319_ (_12872_, _12871_, _06342_);
  nor _64320_ (_12873_, _12733_, _06342_);
  or _64321_ (_12874_, _12873_, _03641_);
  or _64322_ (_12875_, _12874_, _12872_);
  nand _64323_ (_12876_, _10179_, _03641_);
  and _64324_ (_12877_, _12876_, _03161_);
  and _64325_ (_12878_, _12877_, _12875_);
  and _64326_ (_12879_, _10015_, _03160_);
  or _64327_ (_12880_, _12879_, _03435_);
  or _64328_ (_12881_, _12880_, _12878_);
  or _64329_ (_12882_, _12714_, _03436_);
  and _64330_ (_12883_, _12882_, _10843_);
  and _64331_ (_12884_, _12883_, _12881_);
  or _64332_ (_12885_, _12884_, _12699_);
  and _64333_ (_12886_, _12885_, _12444_);
  or _64334_ (_12887_, _12886_, _12695_);
  and _64335_ (_12888_, _12887_, _12265_);
  and _64336_ (_12889_, _12694_, _04212_);
  or _64337_ (_12890_, _12889_, _04544_);
  or _64338_ (_12891_, _12890_, _12888_);
  nor _64339_ (_12892_, _05761_, _05667_);
  nor _64340_ (_12893_, _12892_, _05762_);
  or _64341_ (_12894_, _12893_, _06711_);
  and _64342_ (_12895_, _12894_, _04794_);
  and _64343_ (_12896_, _12895_, _12891_);
  or _64344_ (_12897_, _12896_, _11868_);
  or _64345_ (_12898_, _11867_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _64346_ (_12899_, _12898_, _12049_);
  and _64347_ (_12900_, _12899_, _12897_);
  not _64348_ (_12901_, _09981_);
  nor _64349_ (_12902_, _12901_, _03641_);
  and _64350_ (_12903_, _10138_, _03641_);
  or _64351_ (_12904_, _12903_, _12902_);
  and _64352_ (_12905_, _12904_, _12048_);
  or _64353_ (_40566_, _12905_, _12900_);
  nor _64354_ (_12906_, _08046_, _06721_);
  nor _64355_ (_12907_, _12906_, _06724_);
  or _64356_ (_12908_, _12907_, _06712_);
  nand _64357_ (_12909_, _05422_, _06040_);
  nor _64358_ (_12910_, _10790_, _10766_);
  and _64359_ (_12911_, _10766_, \oc8051_golden_model_1.PSW [7]);
  nor _64360_ (_12912_, _12911_, _12910_);
  nor _64361_ (_12913_, _12912_, _04901_);
  nor _64362_ (_12914_, _10766_, _11682_);
  or _64363_ (_12915_, _12914_, _05778_);
  nor _64364_ (_12916_, _12706_, _05422_);
  or _64365_ (_12917_, _12916_, _05826_);
  and _64366_ (_12918_, _12917_, _05833_);
  nor _64367_ (_12919_, _03923_, _07399_);
  and _64368_ (_12920_, _10010_, _03923_);
  or _64369_ (_12921_, _12920_, _12919_);
  and _64370_ (_12922_, _12921_, _05831_);
  or _64371_ (_12923_, _12922_, _12918_);
  and _64372_ (_12924_, _12923_, _05847_);
  and _64373_ (_12925_, _06721_, _04438_);
  or _64374_ (_12926_, _12925_, _12924_);
  and _64375_ (_12927_, _12926_, _04866_);
  not _64376_ (_12928_, _05945_);
  or _64377_ (_12929_, _12731_, _05471_);
  and _64378_ (_12930_, _12929_, _12928_);
  nor _64379_ (_12931_, _12930_, _04866_);
  or _64380_ (_12932_, _12931_, _12927_);
  and _64381_ (_12933_, _12932_, _05820_);
  nand _64382_ (_12934_, _10767_, _11682_);
  and _64383_ (_12935_, _12934_, _04443_);
  or _64384_ (_12936_, _12935_, _04746_);
  or _64385_ (_12937_, _12936_, _12933_);
  nor _64386_ (_12938_, _10010_, _03203_);
  nor _64387_ (_12939_, _12938_, _04454_);
  and _64388_ (_12940_, _12939_, _12937_);
  and _64389_ (_12941_, _07847_, _04454_);
  or _64390_ (_12942_, _12941_, _04462_);
  or _64391_ (_12943_, _12942_, _12940_);
  and _64392_ (_12944_, _12943_, _12915_);
  or _64393_ (_12945_, _12944_, _03511_);
  nand _64394_ (_12946_, _08205_, _03511_);
  and _64395_ (_12947_, _12946_, _03509_);
  and _64396_ (_12948_, _12947_, _12945_);
  not _64397_ (_12949_, _11683_);
  and _64398_ (_12950_, _12934_, _12949_);
  and _64399_ (_12951_, _12950_, _03508_);
  or _64400_ (_12952_, _12951_, _12948_);
  and _64401_ (_12953_, _12952_, _03200_);
  or _64402_ (_12954_, _10011_, _03200_);
  nand _64403_ (_12955_, _12954_, _03602_);
  or _64404_ (_12956_, _12955_, _12953_);
  nand _64405_ (_12957_, _08205_, _04053_);
  and _64406_ (_12958_, _12957_, _12956_);
  or _64407_ (_12959_, _12958_, _04478_);
  and _64408_ (_12960_, _06721_, _05215_);
  nand _64409_ (_12961_, _08204_, _04478_);
  or _64410_ (_12962_, _12961_, _12960_);
  and _64411_ (_12963_, _12962_, _04901_);
  and _64412_ (_12964_, _12963_, _12959_);
  or _64413_ (_12965_, _12964_, _12913_);
  and _64414_ (_12966_, _12965_, _04853_);
  and _64415_ (_12967_, _10010_, _03223_);
  or _64416_ (_12968_, _12967_, _06040_);
  or _64417_ (_12969_, _12968_, _12966_);
  and _64418_ (_12970_, _12969_, _12909_);
  or _64419_ (_12971_, _12970_, _06045_);
  or _64420_ (_12972_, _06721_, _06051_);
  and _64421_ (_12973_, _12972_, _06050_);
  and _64422_ (_12974_, _12973_, _12971_);
  nor _64423_ (_12975_, _06087_, _05422_);
  and _64424_ (_12976_, _06269_, \oc8051_golden_model_1.IP [5]);
  and _64425_ (_12977_, _06276_, \oc8051_golden_model_1.PSW [5]);
  nor _64426_ (_12978_, _12977_, _12976_);
  and _64427_ (_12979_, _06278_, \oc8051_golden_model_1.ACC [5]);
  and _64428_ (_12980_, _06273_, \oc8051_golden_model_1.B [5]);
  nor _64429_ (_12981_, _12980_, _12979_);
  and _64430_ (_12982_, _12981_, _12978_);
  and _64431_ (_12983_, _06225_, \oc8051_golden_model_1.TL0 [5]);
  not _64432_ (_12984_, _12983_);
  and _64433_ (_12985_, _06245_, \oc8051_golden_model_1.P1INREG [5]);
  and _64434_ (_12986_, _06249_, \oc8051_golden_model_1.P3INREG [5]);
  nor _64435_ (_12987_, _12986_, _12985_);
  and _64436_ (_12988_, _12987_, _12984_);
  and _64437_ (_12989_, _06242_, \oc8051_golden_model_1.P0INREG [5]);
  and _64438_ (_12990_, _06214_, \oc8051_golden_model_1.P2INREG [5]);
  nor _64439_ (_12991_, _12990_, _12989_);
  and _64440_ (_12992_, _12991_, _12988_);
  and _64441_ (_12993_, _06283_, \oc8051_golden_model_1.SP [5]);
  not _64442_ (_12994_, _12993_);
  and _64443_ (_12995_, _06230_, \oc8051_golden_model_1.IE [5]);
  not _64444_ (_12996_, _12995_);
  and _64445_ (_12997_, _06236_, \oc8051_golden_model_1.SCON [5]);
  and _64446_ (_12998_, _06238_, \oc8051_golden_model_1.SBUF [5]);
  nor _64447_ (_12999_, _12998_, _12997_);
  and _64448_ (_13000_, _12999_, _12996_);
  and _64449_ (_13001_, _13000_, _12994_);
  and _64450_ (_13002_, _13001_, _12992_);
  and _64451_ (_13003_, _13002_, _12982_);
  and _64452_ (_13004_, _06256_, \oc8051_golden_model_1.TH0 [5]);
  and _64453_ (_13005_, _06258_, \oc8051_golden_model_1.TL1 [5]);
  nor _64454_ (_13006_, _13005_, _13004_);
  and _64455_ (_13007_, _06263_, \oc8051_golden_model_1.PCON [5]);
  and _64456_ (_13008_, _06265_, \oc8051_golden_model_1.TCON [5]);
  nor _64457_ (_13009_, _13008_, _13007_);
  and _64458_ (_13010_, _13009_, _13006_);
  and _64459_ (_13011_, _06220_, \oc8051_golden_model_1.TMOD [5]);
  and _64460_ (_13012_, _06206_, \oc8051_golden_model_1.TH1 [5]);
  nor _64461_ (_13013_, _13012_, _13011_);
  and _64462_ (_13014_, _06285_, \oc8051_golden_model_1.DPL [5]);
  and _64463_ (_13015_, _06200_, \oc8051_golden_model_1.DPH [5]);
  nor _64464_ (_13016_, _13015_, _13014_);
  and _64465_ (_13017_, _13016_, _13013_);
  and _64466_ (_13018_, _13017_, _13010_);
  and _64467_ (_13019_, _13018_, _13003_);
  not _64468_ (_13020_, _13019_);
  nor _64469_ (_13021_, _13020_, _12975_);
  nor _64470_ (_13022_, _13021_, _06050_);
  or _64471_ (_13023_, _13022_, _06055_);
  or _64472_ (_13024_, _13023_, _12974_);
  and _64473_ (_13025_, _06055_, _03834_);
  nor _64474_ (_13026_, _13025_, _03439_);
  and _64475_ (_13027_, _13026_, _13024_);
  and _64476_ (_13028_, _06211_, _03439_);
  or _64477_ (_13029_, _13028_, _03189_);
  or _64478_ (_13030_, _13029_, _13027_);
  and _64479_ (_13031_, _10011_, _03189_);
  nor _64480_ (_13032_, _13031_, _04500_);
  and _64481_ (_13033_, _13032_, _13030_);
  nor _64482_ (_13034_, _06164_, _05471_);
  and _64483_ (_13035_, _06164_, _05471_);
  nor _64484_ (_13036_, _13035_, _13034_);
  and _64485_ (_13037_, _13036_, _04500_);
  or _64486_ (_13038_, _13037_, _13033_);
  and _64487_ (_13039_, _13038_, _05772_);
  nor _64488_ (_13040_, _05471_, _07399_);
  and _64489_ (_13041_, _05471_, _07399_);
  nor _64490_ (_13042_, _13041_, _13040_);
  and _64491_ (_13043_, _13042_, _04502_);
  or _64492_ (_13044_, _13043_, _04506_);
  or _64493_ (_13045_, _13044_, _13039_);
  or _64494_ (_13046_, _13034_, _04507_);
  and _64495_ (_13047_, _13046_, _04498_);
  and _64496_ (_13048_, _13047_, _13045_);
  and _64497_ (_13049_, _13040_, _04497_);
  or _64498_ (_13050_, _13049_, _03192_);
  or _64499_ (_13051_, _13050_, _13048_);
  and _64500_ (_13052_, _10011_, _03192_);
  nor _64501_ (_13053_, _13052_, _04516_);
  and _64502_ (_13054_, _13053_, _13051_);
  and _64503_ (_13055_, _13035_, _06324_);
  nor _64504_ (_13056_, _13055_, _04519_);
  or _64505_ (_13057_, _13056_, _13054_);
  nand _64506_ (_13058_, _13041_, _04518_);
  and _64507_ (_13059_, _13058_, _06328_);
  and _64508_ (_13060_, _13059_, _13057_);
  and _64509_ (_13061_, _07777_, _03665_);
  nor _64510_ (_13062_, _13061_, _12061_);
  and _64511_ (_13063_, _10010_, _03179_);
  or _64512_ (_13064_, _13063_, _13062_);
  or _64513_ (_13065_, _13064_, _13060_);
  and _64514_ (_13066_, _12917_, _12227_);
  or _64515_ (_13067_, _13066_, _12013_);
  and _64516_ (_13068_, _13067_, _13065_);
  and _64517_ (_13069_, _12917_, _04194_);
  or _64518_ (_13070_, _13069_, _04527_);
  or _64519_ (_13071_, _13070_, _13068_);
  nor _64520_ (_13072_, _12700_, _06616_);
  or _64521_ (_13073_, _06663_, _06343_);
  or _64522_ (_13074_, _13073_, _13072_);
  and _64523_ (_13075_, _13074_, _06342_);
  and _64524_ (_13076_, _13075_, _13071_);
  nor _64525_ (_13077_, _12930_, _06342_);
  or _64526_ (_13078_, _13077_, _03641_);
  or _64527_ (_13079_, _13078_, _13076_);
  nand _64528_ (_13080_, _10174_, _03641_);
  and _64529_ (_13081_, _13080_, _03161_);
  and _64530_ (_13082_, _13081_, _13079_);
  and _64531_ (_13083_, _10010_, _03160_);
  or _64532_ (_13084_, _13083_, _03435_);
  or _64533_ (_13085_, _13084_, _13082_);
  or _64534_ (_13086_, _12910_, _03436_);
  and _64535_ (_13087_, _13086_, _10843_);
  and _64536_ (_13088_, _13087_, _13085_);
  or _64537_ (_13089_, _12697_, _07847_);
  nor _64538_ (_13090_, _10843_, _06697_);
  and _64539_ (_13091_, _13090_, _13089_);
  or _64540_ (_13092_, _13091_, _04540_);
  or _64541_ (_13093_, _13092_, _13088_);
  and _64542_ (_13094_, _13093_, _12908_);
  or _64543_ (_13095_, _13094_, _04544_);
  nor _64544_ (_13096_, _05762_, _05472_);
  nor _64545_ (_13097_, _13096_, _05763_);
  or _64546_ (_13098_, _13097_, _06711_);
  and _64547_ (_13099_, _13098_, _04794_);
  and _64548_ (_13100_, _13099_, _13095_);
  or _64549_ (_13101_, _13100_, _11868_);
  or _64550_ (_13102_, _11867_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _64551_ (_13103_, _13102_, _12049_);
  and _64552_ (_13104_, _13103_, _13101_);
  and _64553_ (_13105_, _09977_, _10832_);
  and _64554_ (_13106_, _10133_, _03641_);
  or _64555_ (_13107_, _13106_, _13105_);
  and _64556_ (_13108_, _13107_, _12685_);
  and _64557_ (_13109_, _13108_, _42963_);
  and _64558_ (_13110_, _13109_, _41755_);
  and _64559_ (_13111_, _13110_, _12684_);
  or _64560_ (_40567_, _13111_, _13104_);
  nor _64561_ (_13112_, _06724_, _06713_);
  nor _64562_ (_13113_, _13112_, _06725_);
  and _64563_ (_13114_, _13113_, _12443_);
  nor _64564_ (_13115_, _04967_, _04207_);
  not _64565_ (_13116_, _13115_);
  and _64566_ (_13117_, _06697_, _05327_);
  nor _64567_ (_13118_, _06697_, _05327_);
  or _64568_ (_13119_, _13118_, _13117_);
  and _64569_ (_13120_, _13119_, _13116_);
  nor _64570_ (_13121_, _05945_, _05376_);
  nor _64571_ (_13122_, _13121_, _05946_);
  nor _64572_ (_13123_, _13122_, _06342_);
  nor _64573_ (_13124_, _06663_, _06388_);
  or _64574_ (_13125_, _13124_, _06664_);
  and _64575_ (_13126_, _13125_, _04527_);
  nor _64576_ (_13127_, _05826_, _05327_);
  or _64577_ (_13128_, _13127_, _05827_);
  or _64578_ (_13129_, _13128_, _04709_);
  nor _64579_ (_13130_, _10709_, _11658_);
  or _64580_ (_13131_, _13130_, _05778_);
  nor _64581_ (_13132_, _03923_, _07346_);
  and _64582_ (_13133_, _10003_, _03923_);
  or _64583_ (_13134_, _13133_, _13132_);
  and _64584_ (_13135_, _13134_, _05831_);
  and _64585_ (_13136_, _13128_, _05833_);
  or _64586_ (_13137_, _13136_, _13135_);
  and _64587_ (_13138_, _13137_, _05847_);
  and _64588_ (_13139_, _06713_, _04438_);
  or _64589_ (_13140_, _13139_, _13138_);
  and _64590_ (_13141_, _13140_, _04866_);
  nor _64591_ (_13142_, _13122_, _04866_);
  or _64592_ (_13143_, _13142_, _13141_);
  and _64593_ (_13144_, _13143_, _05820_);
  nand _64594_ (_13145_, _10710_, _11658_);
  and _64595_ (_13146_, _13145_, _04443_);
  or _64596_ (_13147_, _13146_, _04746_);
  or _64597_ (_13148_, _13147_, _13144_);
  nor _64598_ (_13149_, _10003_, _03203_);
  nor _64599_ (_13150_, _13149_, _04454_);
  and _64600_ (_13151_, _13150_, _13148_);
  and _64601_ (_13152_, _07831_, _04454_);
  or _64602_ (_13153_, _13152_, _04462_);
  or _64603_ (_13154_, _13153_, _13151_);
  and _64604_ (_13155_, _13154_, _13131_);
  or _64605_ (_13156_, _13155_, _03511_);
  nand _64606_ (_13157_, _08125_, _03511_);
  and _64607_ (_13158_, _13157_, _03509_);
  and _64608_ (_13159_, _13158_, _13156_);
  not _64609_ (_13160_, _11659_);
  and _64610_ (_13161_, _13145_, _13160_);
  and _64611_ (_13162_, _13161_, _03508_);
  or _64612_ (_13163_, _13162_, _13159_);
  and _64613_ (_13164_, _13163_, _03200_);
  or _64614_ (_13165_, _10004_, _03200_);
  nand _64615_ (_13166_, _13165_, _03602_);
  or _64616_ (_13167_, _13166_, _13164_);
  nand _64617_ (_13168_, _08125_, _04053_);
  and _64618_ (_13169_, _13168_, _13167_);
  or _64619_ (_13170_, _13169_, _04478_);
  and _64620_ (_13171_, _06713_, _05215_);
  nand _64621_ (_13172_, _08124_, _04478_);
  or _64622_ (_13173_, _13172_, _13171_);
  and _64623_ (_13174_, _13173_, _04901_);
  and _64624_ (_13175_, _13174_, _13170_);
  nor _64625_ (_13176_, _10736_, _10709_);
  and _64626_ (_13177_, _10709_, \oc8051_golden_model_1.PSW [7]);
  nor _64627_ (_13178_, _13177_, _13176_);
  nor _64628_ (_13179_, _13178_, _04901_);
  or _64629_ (_13180_, _13179_, _03223_);
  or _64630_ (_13181_, _13180_, _13175_);
  and _64631_ (_13182_, _10004_, _03223_);
  nor _64632_ (_13183_, _13182_, _06040_);
  and _64633_ (_13184_, _13183_, _13181_);
  nor _64634_ (_13185_, _05327_, _06046_);
  or _64635_ (_13186_, _13185_, _06045_);
  or _64636_ (_13187_, _13186_, _13184_);
  or _64637_ (_13188_, _06713_, _06051_);
  and _64638_ (_13189_, _13188_, _06050_);
  and _64639_ (_13190_, _13189_, _13187_);
  nor _64640_ (_13191_, _06087_, _05327_);
  and _64641_ (_13192_, _06269_, \oc8051_golden_model_1.IP [6]);
  and _64642_ (_13193_, _06273_, \oc8051_golden_model_1.B [6]);
  nor _64643_ (_13194_, _13193_, _13192_);
  and _64644_ (_13195_, _06276_, \oc8051_golden_model_1.PSW [6]);
  and _64645_ (_13196_, _06278_, \oc8051_golden_model_1.ACC [6]);
  nor _64646_ (_13197_, _13196_, _13195_);
  and _64647_ (_13198_, _13197_, _13194_);
  and _64648_ (_13199_, _06225_, \oc8051_golden_model_1.TL0 [6]);
  not _64649_ (_13200_, _13199_);
  and _64650_ (_13201_, _06245_, \oc8051_golden_model_1.P1INREG [6]);
  and _64651_ (_13202_, _06249_, \oc8051_golden_model_1.P3INREG [6]);
  nor _64652_ (_13203_, _13202_, _13201_);
  and _64653_ (_13204_, _13203_, _13200_);
  and _64654_ (_13205_, _06242_, \oc8051_golden_model_1.P0INREG [6]);
  and _64655_ (_13206_, _06214_, \oc8051_golden_model_1.P2INREG [6]);
  nor _64656_ (_13207_, _13206_, _13205_);
  and _64657_ (_13208_, _13207_, _13204_);
  and _64658_ (_13209_, _06283_, \oc8051_golden_model_1.SP [6]);
  not _64659_ (_13210_, _13209_);
  and _64660_ (_13211_, _06230_, \oc8051_golden_model_1.IE [6]);
  not _64661_ (_13212_, _13211_);
  and _64662_ (_13213_, _06236_, \oc8051_golden_model_1.SCON [6]);
  and _64663_ (_13214_, _06238_, \oc8051_golden_model_1.SBUF [6]);
  nor _64664_ (_13215_, _13214_, _13213_);
  and _64665_ (_13216_, _13215_, _13212_);
  and _64666_ (_13217_, _13216_, _13210_);
  and _64667_ (_13218_, _13217_, _13208_);
  and _64668_ (_13219_, _13218_, _13198_);
  and _64669_ (_13220_, _06256_, \oc8051_golden_model_1.TH0 [6]);
  and _64670_ (_13221_, _06258_, \oc8051_golden_model_1.TL1 [6]);
  nor _64671_ (_13222_, _13221_, _13220_);
  and _64672_ (_13223_, _06263_, \oc8051_golden_model_1.PCON [6]);
  and _64673_ (_13224_, _06265_, \oc8051_golden_model_1.TCON [6]);
  nor _64674_ (_13225_, _13224_, _13223_);
  and _64675_ (_13226_, _13225_, _13222_);
  and _64676_ (_13227_, _06220_, \oc8051_golden_model_1.TMOD [6]);
  and _64677_ (_13228_, _06206_, \oc8051_golden_model_1.TH1 [6]);
  nor _64678_ (_13229_, _13228_, _13227_);
  and _64679_ (_13230_, _06285_, \oc8051_golden_model_1.DPL [6]);
  and _64680_ (_13231_, _06200_, \oc8051_golden_model_1.DPH [6]);
  nor _64681_ (_13232_, _13231_, _13230_);
  and _64682_ (_13233_, _13232_, _13229_);
  and _64683_ (_13234_, _13233_, _13226_);
  and _64684_ (_13235_, _13234_, _13219_);
  not _64685_ (_13236_, _13235_);
  nor _64686_ (_13237_, _13236_, _13191_);
  nor _64687_ (_13238_, _13237_, _06050_);
  or _64688_ (_13239_, _13238_, _06055_);
  or _64689_ (_13240_, _13239_, _13190_);
  and _64690_ (_13241_, _06055_, _03561_);
  nor _64691_ (_13242_, _13241_, _03439_);
  and _64692_ (_13243_, _13242_, _13240_);
  not _64693_ (_13244_, _06132_);
  and _64694_ (_13245_, _13244_, _03439_);
  or _64695_ (_13246_, _13245_, _03189_);
  or _64696_ (_13247_, _13246_, _13243_);
  and _64697_ (_13248_, _10004_, _03189_);
  nor _64698_ (_13249_, _13248_, _04500_);
  and _64699_ (_13250_, _13249_, _13247_);
  and _64700_ (_13251_, _06132_, _05376_);
  nor _64701_ (_13252_, _06132_, _05376_);
  nor _64702_ (_13253_, _13252_, _13251_);
  nor _64703_ (_13254_, _13253_, _04502_);
  nor _64704_ (_13255_, _13254_, _04503_);
  or _64705_ (_13256_, _13255_, _13250_);
  nor _64706_ (_13257_, _05376_, _07346_);
  and _64707_ (_13258_, _05376_, _07346_);
  nor _64708_ (_13259_, _13258_, _13257_);
  or _64709_ (_13260_, _13259_, _05772_);
  and _64710_ (_13261_, _13260_, _04507_);
  and _64711_ (_13262_, _13261_, _13256_);
  and _64712_ (_13263_, _13252_, _05770_);
  or _64713_ (_13264_, _13263_, _13262_);
  and _64714_ (_13265_, _13264_, _04498_);
  and _64715_ (_13266_, _13257_, _04497_);
  or _64716_ (_13267_, _13266_, _03192_);
  or _64717_ (_13268_, _13267_, _13265_);
  and _64718_ (_13269_, _10004_, _03192_);
  nor _64719_ (_13270_, _13269_, _04516_);
  and _64720_ (_13271_, _13270_, _13268_);
  and _64721_ (_13272_, _13251_, _06324_);
  nor _64722_ (_13273_, _13272_, _04519_);
  or _64723_ (_13274_, _13273_, _13271_);
  nand _64724_ (_13275_, _13258_, _04518_);
  and _64725_ (_13276_, _13275_, _06328_);
  and _64726_ (_13277_, _13276_, _13274_);
  nand _64727_ (_13278_, _10003_, _03179_);
  nand _64728_ (_13279_, _13278_, _04709_);
  or _64729_ (_13280_, _13279_, _13277_);
  and _64730_ (_13281_, _13280_, _13129_);
  or _64731_ (_13282_, _13281_, _04681_);
  or _64732_ (_13283_, _13128_, _06335_);
  and _64733_ (_13284_, _13283_, _06343_);
  and _64734_ (_13285_, _13284_, _13282_);
  or _64735_ (_13286_, _13285_, _13126_);
  and _64736_ (_13287_, _13286_, _06342_);
  or _64737_ (_13288_, _13287_, _13123_);
  and _64738_ (_13289_, _13288_, _10832_);
  and _64739_ (_13290_, _10165_, _03641_);
  or _64740_ (_13291_, _13290_, _03160_);
  or _64741_ (_13292_, _13291_, _13289_);
  and _64742_ (_13293_, _10004_, _03160_);
  nor _64743_ (_13294_, _13293_, _03435_);
  and _64744_ (_13295_, _13294_, _13292_);
  and _64745_ (_13296_, _03484_, _03165_);
  and _64746_ (_13297_, _13176_, _03435_);
  or _64747_ (_13298_, _13297_, _13296_);
  or _64748_ (_13299_, _13298_, _13295_);
  not _64749_ (_13300_, _13296_);
  or _64750_ (_13301_, _13119_, _13300_);
  and _64751_ (_13302_, _13301_, _13115_);
  and _64752_ (_13303_, _13302_, _13299_);
  or _64753_ (_13304_, _13303_, _13120_);
  and _64754_ (_13305_, _13304_, _12444_);
  or _64755_ (_13306_, _13305_, _13114_);
  and _64756_ (_13307_, _13306_, _12265_);
  and _64757_ (_13308_, _13113_, _04212_);
  or _64758_ (_13309_, _13308_, _04544_);
  or _64759_ (_13310_, _13309_, _13307_);
  nor _64760_ (_13311_, _05763_, _05377_);
  nor _64761_ (_13312_, _13311_, _05764_);
  or _64762_ (_13313_, _13312_, _06711_);
  and _64763_ (_13314_, _13313_, _04794_);
  and _64764_ (_13315_, _13314_, _13310_);
  or _64765_ (_13316_, _13315_, _11868_);
  or _64766_ (_13317_, _11867_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _64767_ (_13318_, _13317_, _12049_);
  and _64768_ (_13319_, _13318_, _13316_);
  and _64769_ (_13320_, _09971_, _10832_);
  and _64770_ (_13321_, _10126_, _03641_);
  or _64771_ (_13322_, _13321_, _13320_);
  and _64772_ (_13323_, _13322_, _12048_);
  or _64773_ (_40569_, _13323_, _13319_);
  or _64774_ (_13324_, _11868_, _06732_);
  or _64775_ (_13325_, _11867_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _64776_ (_13326_, _13325_, _12049_);
  and _64777_ (_13327_, _13326_, _13324_);
  and _64778_ (_13328_, _06756_, _12685_);
  and _64779_ (_13329_, _13328_, _42963_);
  and _64780_ (_13330_, _13329_, _41755_);
  and _64781_ (_13331_, _12684_, _13330_);
  or _64782_ (_40570_, _13331_, _13327_);
  nand _64783_ (_13332_, _12047_, _04845_);
  or _64784_ (_13333_, _13332_, _12055_);
  and _64785_ (_13334_, _11862_, _04700_);
  and _64786_ (_13335_, _13334_, _11865_);
  and _64787_ (_13336_, _13335_, _12043_);
  or _64788_ (_13337_, _13335_, _04369_);
  nand _64789_ (_13338_, _13337_, _13332_);
  or _64790_ (_13339_, _13338_, _13336_);
  and _64791_ (_40574_, _13339_, _13333_);
  not _64792_ (_13340_, _13335_);
  or _64793_ (_13341_, _13340_, _12255_);
  or _64794_ (_13342_, _13335_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _64795_ (_13343_, _13342_, _13332_);
  and _64796_ (_13344_, _13343_, _13341_);
  and _64797_ (_13345_, _12263_, _12685_);
  and _64798_ (_13346_, _13345_, _42963_);
  and _64799_ (_13347_, _13346_, _41755_);
  not _64800_ (_13348_, _12672_);
  and _64801_ (_13349_, _13348_, _12669_);
  and _64802_ (_13350_, _13349_, _12682_);
  and _64803_ (_13351_, _13350_, _13347_);
  or _64804_ (_40576_, _13351_, _13344_);
  or _64805_ (_13352_, _13340_, _12459_);
  or _64806_ (_13353_, _13335_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _64807_ (_13354_, _13353_, _13332_);
  and _64808_ (_13355_, _13354_, _13352_);
  and _64809_ (_13356_, _12467_, _12685_);
  and _64810_ (_13357_, _13356_, _42963_);
  and _64811_ (_13358_, _13357_, _41755_);
  and _64812_ (_13359_, _13350_, _13358_);
  or _64813_ (_40577_, _13359_, _13355_);
  or _64814_ (_13360_, _13340_, _12661_);
  or _64815_ (_13361_, _13335_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _64816_ (_13362_, _13361_, _13332_);
  and _64817_ (_13363_, _13362_, _13360_);
  and _64818_ (_13364_, _13350_, _12691_);
  or _64819_ (_40578_, _13364_, _13363_);
  or _64820_ (_13365_, _13340_, _12896_);
  or _64821_ (_13366_, _13335_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _64822_ (_13367_, _13366_, _13332_);
  and _64823_ (_13368_, _13367_, _13365_);
  and _64824_ (_13369_, _12904_, _12685_);
  and _64825_ (_13370_, _13369_, _42963_);
  and _64826_ (_13371_, _13370_, _41755_);
  and _64827_ (_13372_, _13350_, _13371_);
  or _64828_ (_40579_, _13372_, _13368_);
  or _64829_ (_13373_, _13340_, _13100_);
  or _64830_ (_13374_, _13335_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _64831_ (_13375_, _13374_, _13332_);
  and _64832_ (_13376_, _13375_, _13373_);
  and _64833_ (_13377_, _13350_, _13110_);
  or _64834_ (_40580_, _13377_, _13376_);
  or _64835_ (_13378_, _13340_, _13315_);
  or _64836_ (_13379_, _13335_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _64837_ (_13380_, _13379_, _13332_);
  and _64838_ (_13381_, _13380_, _13378_);
  and _64839_ (_13382_, _13322_, _12685_);
  and _64840_ (_13383_, _13382_, _42963_);
  and _64841_ (_13384_, _13383_, _41755_);
  and _64842_ (_13385_, _13350_, _13384_);
  or _64843_ (_40582_, _13385_, _13381_);
  or _64844_ (_13386_, _13340_, _06733_);
  or _64845_ (_13387_, _13335_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _64846_ (_13388_, _13387_, _13332_);
  and _64847_ (_13389_, _13388_, _13386_);
  and _64848_ (_13390_, _13350_, _13330_);
  or _64849_ (_40583_, _13390_, _13389_);
  not _64850_ (_13391_, _04796_);
  nor _64851_ (_13392_, _13391_, _04547_);
  and _64852_ (_13393_, _13392_, _11865_);
  not _64853_ (_13394_, _13393_);
  or _64854_ (_13395_, _13394_, _12043_);
  and _64855_ (_13396_, _05117_, _05110_);
  nor _64856_ (_13397_, _05118_, _13396_);
  and _64857_ (_13398_, _13397_, _05117_);
  and _64858_ (_13399_, _13398_, _05848_);
  not _64859_ (_13400_, _13399_);
  or _64860_ (_13401_, _13393_, \oc8051_golden_model_1.IRAM[2] [0]);
  and _64861_ (_13402_, _13401_, _13400_);
  and _64862_ (_13403_, _13402_, _13395_);
  and _64863_ (_13404_, _12055_, _05117_);
  and _64864_ (_13405_, _13399_, _13404_);
  or _64865_ (_40587_, _13405_, _13403_);
  or _64866_ (_13406_, _13394_, _12255_);
  and _64867_ (_13407_, _12047_, _05848_);
  not _64868_ (_13408_, _13407_);
  or _64869_ (_13409_, _13393_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _64870_ (_13410_, _13409_, _13408_);
  and _64871_ (_13411_, _13410_, _13406_);
  and _64872_ (_13412_, _12263_, _05117_);
  and _64873_ (_13413_, _13412_, _13407_);
  or _64874_ (_40588_, _13413_, _13411_);
  or _64875_ (_13414_, _13394_, _12459_);
  or _64876_ (_13415_, _13393_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _64877_ (_13416_, _13415_, _13408_);
  and _64878_ (_13417_, _13416_, _13414_);
  and _64879_ (_13418_, _12467_, _05117_);
  and _64880_ (_13419_, _13418_, _13407_);
  or _64881_ (_40589_, _13419_, _13417_);
  or _64882_ (_13420_, _13394_, _12661_);
  or _64883_ (_13421_, _13393_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _64884_ (_13422_, _13421_, _13400_);
  and _64885_ (_13423_, _13422_, _13420_);
  and _64886_ (_13424_, _12688_, _05117_);
  and _64887_ (_13425_, _13424_, _13399_);
  or _64888_ (_40591_, _13425_, _13423_);
  or _64889_ (_13426_, _13394_, _12896_);
  or _64890_ (_13427_, _13393_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _64891_ (_13428_, _13427_, _13408_);
  and _64892_ (_13429_, _13428_, _13426_);
  and _64893_ (_13430_, _12904_, _05117_);
  and _64894_ (_13431_, _13430_, _13407_);
  or _64895_ (_40592_, _13431_, _13429_);
  or _64896_ (_13432_, _13394_, _13100_);
  or _64897_ (_13433_, _13393_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _64898_ (_13434_, _13433_, _13408_);
  and _64899_ (_13435_, _13434_, _13432_);
  and _64900_ (_13436_, _13107_, _05117_);
  and _64901_ (_13437_, _13436_, _13407_);
  or _64902_ (_40593_, _13437_, _13435_);
  or _64903_ (_13438_, _13394_, _13315_);
  or _64904_ (_13439_, _13393_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _64905_ (_13440_, _13439_, _13408_);
  and _64906_ (_13441_, _13440_, _13438_);
  and _64907_ (_13442_, _13322_, _05117_);
  and _64908_ (_13443_, _13442_, _13407_);
  or _64909_ (_40594_, _13443_, _13441_);
  or _64910_ (_13444_, _13394_, _06733_);
  or _64911_ (_13445_, _13393_, \oc8051_golden_model_1.IRAM[2] [7]);
  and _64912_ (_13446_, _13445_, _13408_);
  and _64913_ (_13447_, _13446_, _13444_);
  and _64914_ (_13448_, _13407_, _06757_);
  or _64915_ (_40595_, _13448_, _13447_);
  and _64916_ (_13449_, _11865_, _04797_);
  or _64917_ (_13450_, _13449_, \oc8051_golden_model_1.IRAM[3] [0]);
  and _64918_ (_13451_, _12047_, _04550_);
  not _64919_ (_13452_, _13451_);
  not _64920_ (_13453_, _13449_);
  or _64921_ (_13454_, _13453_, _12043_);
  and _64922_ (_13455_, _13454_, _13452_);
  and _64923_ (_13456_, _13455_, _13450_);
  and _64924_ (_13457_, _13451_, _13404_);
  or _64925_ (_40599_, _13457_, _13456_);
  or _64926_ (_13458_, _13449_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _64927_ (_13459_, _13458_, _13452_);
  or _64928_ (_13460_, _13453_, _12255_);
  and _64929_ (_13461_, _13460_, _13459_);
  and _64930_ (_13462_, _12672_, _12669_);
  and _64931_ (_13463_, _12682_, _13462_);
  and _64932_ (_13464_, _13463_, _13347_);
  or _64933_ (_40601_, _13464_, _13461_);
  or _64934_ (_13465_, _13449_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _64935_ (_13466_, _13465_, _13452_);
  or _64936_ (_13467_, _13453_, _12459_);
  and _64937_ (_13468_, _13467_, _13466_);
  and _64938_ (_13469_, _13463_, _13358_);
  or _64939_ (_40602_, _13469_, _13468_);
  or _64940_ (_13470_, _13449_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _64941_ (_13471_, _13470_, _13452_);
  or _64942_ (_13472_, _13453_, _12661_);
  and _64943_ (_13473_, _13472_, _13471_);
  and _64944_ (_13474_, _13451_, _13424_);
  or _64945_ (_40603_, _13474_, _13473_);
  or _64946_ (_13475_, _13449_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _64947_ (_13476_, _13475_, _13452_);
  or _64948_ (_13477_, _13453_, _12896_);
  and _64949_ (_13478_, _13477_, _13476_);
  and _64950_ (_13479_, _13463_, _13371_);
  or _64951_ (_40604_, _13479_, _13478_);
  or _64952_ (_13480_, _13449_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _64953_ (_13481_, _13480_, _13452_);
  or _64954_ (_13482_, _13453_, _13100_);
  and _64955_ (_13483_, _13482_, _13481_);
  and _64956_ (_13484_, _13451_, _13436_);
  or _64957_ (_40605_, _13484_, _13483_);
  or _64958_ (_13485_, _13449_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _64959_ (_13486_, _13485_, _13452_);
  or _64960_ (_13487_, _13453_, _13315_);
  and _64961_ (_13488_, _13487_, _13486_);
  and _64962_ (_13489_, _13463_, _13384_);
  or _64963_ (_40607_, _13489_, _13488_);
  or _64964_ (_13490_, _13449_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _64965_ (_13491_, _13490_, _13452_);
  or _64966_ (_13492_, _13453_, _06733_);
  and _64967_ (_13493_, _13492_, _13491_);
  and _64968_ (_13494_, _13451_, _06757_);
  or _64969_ (_40608_, _13494_, _13493_);
  and _64970_ (_13495_, _05103_, _04964_);
  and _64971_ (_13496_, _13495_, _11863_);
  not _64972_ (_13497_, _13496_);
  or _64973_ (_13498_, _13497_, _12043_);
  or _64974_ (_13499_, _13496_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _64975_ (_13500_, _13396_, _12678_);
  and _64976_ (_13501_, _13500_, _04551_);
  not _64977_ (_13502_, _13501_);
  and _64978_ (_13503_, _13502_, _13499_);
  and _64979_ (_13504_, _13503_, _13498_);
  and _64980_ (_13505_, _13501_, _13404_);
  or _64981_ (_40612_, _13505_, _13504_);
  or _64982_ (_13506_, _13497_, _12255_);
  or _64983_ (_13507_, _13496_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _64984_ (_13508_, _13507_, _13502_);
  and _64985_ (_13509_, _13508_, _13506_);
  and _64986_ (_13510_, _13501_, _13412_);
  or _64987_ (_40613_, _13510_, _13509_);
  or _64988_ (_13511_, _13497_, _12459_);
  or _64989_ (_13512_, _13496_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _64990_ (_13513_, _13512_, _13502_);
  and _64991_ (_13514_, _13513_, _13511_);
  and _64992_ (_13515_, _13501_, _13418_);
  or _64993_ (_40614_, _13515_, _13514_);
  or _64994_ (_13516_, _13497_, _12661_);
  or _64995_ (_13517_, _13496_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _64996_ (_13518_, _13517_, _13502_);
  and _64997_ (_13519_, _13518_, _13516_);
  and _64998_ (_13520_, _13501_, _13424_);
  or _64999_ (_40616_, _13520_, _13519_);
  or _65000_ (_13521_, _13497_, _12896_);
  or _65001_ (_13522_, _13496_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _65002_ (_13523_, _13522_, _13502_);
  and _65003_ (_13524_, _13523_, _13521_);
  and _65004_ (_13525_, _13501_, _13430_);
  or _65005_ (_40617_, _13525_, _13524_);
  or _65006_ (_13526_, _13497_, _13100_);
  or _65007_ (_13527_, _13496_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _65008_ (_13528_, _13527_, _13502_);
  and _65009_ (_13529_, _13528_, _13526_);
  and _65010_ (_13530_, _13501_, _13436_);
  or _65011_ (_40618_, _13530_, _13529_);
  or _65012_ (_13531_, _13497_, _13315_);
  or _65013_ (_13532_, _13496_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _65014_ (_13533_, _13532_, _13502_);
  and _65015_ (_13534_, _13533_, _13531_);
  and _65016_ (_13535_, _13501_, _13442_);
  or _65017_ (_40619_, _13535_, _13534_);
  or _65018_ (_13536_, _13497_, _06733_);
  or _65019_ (_13537_, _13496_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _65020_ (_13538_, _13537_, _13502_);
  and _65021_ (_13539_, _13538_, _13536_);
  and _65022_ (_13540_, _13501_, _06757_);
  or _65023_ (_40620_, _13540_, _13539_);
  and _65024_ (_13541_, _13500_, _04845_);
  not _65025_ (_13542_, _13541_);
  or _65026_ (_13543_, _13542_, _13404_);
  and _65027_ (_13544_, _13495_, _13334_);
  and _65028_ (_13545_, _13544_, _12043_);
  nor _65029_ (_13546_, _13544_, _04388_);
  or _65030_ (_13547_, _13546_, _13541_);
  or _65031_ (_13548_, _13547_, _13545_);
  and _65032_ (_40624_, _13548_, _13543_);
  not _65033_ (_13549_, _13544_);
  or _65034_ (_13550_, _13549_, _12255_);
  or _65035_ (_13551_, _13544_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _65036_ (_13552_, _13551_, _13542_);
  and _65037_ (_13553_, _13552_, _13550_);
  and _65038_ (_13554_, _13541_, _13412_);
  or _65039_ (_40625_, _13554_, _13553_);
  or _65040_ (_13555_, _13549_, _12459_);
  or _65041_ (_13556_, _13544_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _65042_ (_13557_, _13556_, _13542_);
  and _65043_ (_13558_, _13557_, _13555_);
  and _65044_ (_13559_, _13541_, _13418_);
  or _65045_ (_40627_, _13559_, _13558_);
  or _65046_ (_13560_, _13549_, _12661_);
  or _65047_ (_13561_, _13544_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _65048_ (_13562_, _13561_, _13542_);
  and _65049_ (_13563_, _13562_, _13560_);
  and _65050_ (_13564_, _13541_, _13424_);
  or _65051_ (_40628_, _13564_, _13563_);
  or _65052_ (_13565_, _13549_, _12896_);
  or _65053_ (_13566_, _13544_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _65054_ (_13567_, _13566_, _13542_);
  and _65055_ (_13568_, _13567_, _13565_);
  and _65056_ (_13569_, _13541_, _13430_);
  or _65057_ (_40629_, _13569_, _13568_);
  or _65058_ (_13570_, _13549_, _13100_);
  or _65059_ (_13571_, _13544_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _65060_ (_13572_, _13571_, _13542_);
  and _65061_ (_13573_, _13572_, _13570_);
  and _65062_ (_13574_, _13541_, _13436_);
  or _65063_ (_40630_, _13574_, _13573_);
  or _65064_ (_13575_, _13549_, _13315_);
  or _65065_ (_13576_, _13544_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _65066_ (_13577_, _13576_, _13542_);
  and _65067_ (_13578_, _13577_, _13575_);
  and _65068_ (_13579_, _13541_, _13442_);
  or _65069_ (_40631_, _13579_, _13578_);
  or _65070_ (_13580_, _13549_, _06733_);
  or _65071_ (_13581_, _13544_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _65072_ (_13582_, _13581_, _13542_);
  and _65073_ (_13583_, _13582_, _13580_);
  and _65074_ (_13584_, _13541_, _06757_);
  or _65075_ (_40633_, _13584_, _13583_);
  and _65076_ (_13585_, _13495_, _13392_);
  not _65077_ (_13586_, _13585_);
  or _65078_ (_13587_, _13586_, _12043_);
  or _65079_ (_13588_, _13585_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _65080_ (_13589_, _13500_, _05848_);
  not _65081_ (_13590_, _13589_);
  and _65082_ (_13591_, _13590_, _13588_);
  and _65083_ (_13592_, _13591_, _13587_);
  and _65084_ (_13593_, _13589_, _13404_);
  or _65085_ (_40636_, _13593_, _13592_);
  or _65086_ (_13594_, _13586_, _12255_);
  or _65087_ (_13595_, _13585_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _65088_ (_13596_, _13595_, _13590_);
  and _65089_ (_13597_, _13596_, _13594_);
  and _65090_ (_13598_, _13589_, _13412_);
  or _65091_ (_40637_, _13598_, _13597_);
  or _65092_ (_13600_, _13586_, _12459_);
  or _65093_ (_13601_, _13585_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _65094_ (_13602_, _13601_, _13590_);
  and _65095_ (_13603_, _13602_, _13600_);
  and _65096_ (_13604_, _13589_, _13418_);
  or _65097_ (_40639_, _13604_, _13603_);
  or _65098_ (_13605_, _13586_, _12661_);
  or _65099_ (_13606_, _13585_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _65100_ (_13607_, _13606_, _13590_);
  and _65101_ (_13609_, _13607_, _13605_);
  and _65102_ (_13610_, _13589_, _13424_);
  or _65103_ (_40640_, _13610_, _13609_);
  or _65104_ (_13611_, _13586_, _12896_);
  or _65105_ (_13612_, _13585_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _65106_ (_13613_, _13612_, _13590_);
  and _65107_ (_13614_, _13613_, _13611_);
  and _65108_ (_13615_, _13589_, _13430_);
  or _65109_ (_40641_, _13615_, _13614_);
  or _65110_ (_13616_, _13586_, _13100_);
  or _65111_ (_13618_, _13585_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _65112_ (_13619_, _13618_, _13590_);
  and _65113_ (_13620_, _13619_, _13616_);
  and _65114_ (_13621_, _13589_, _13436_);
  or _65115_ (_40642_, _13621_, _13620_);
  or _65116_ (_13622_, _13586_, _13315_);
  or _65117_ (_13623_, _13585_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _65118_ (_13624_, _13623_, _13590_);
  and _65119_ (_13625_, _13624_, _13622_);
  and _65120_ (_13626_, _13589_, _13442_);
  or _65121_ (_40643_, _13626_, _13625_);
  or _65122_ (_13628_, _13586_, _06733_);
  or _65123_ (_13629_, _13585_, \oc8051_golden_model_1.IRAM[6] [7]);
  and _65124_ (_13630_, _13629_, _13590_);
  and _65125_ (_13631_, _13630_, _13628_);
  and _65126_ (_13632_, _13589_, _06757_);
  or _65127_ (_40645_, _13632_, _13631_);
  not _65128_ (_13633_, _04700_);
  and _65129_ (_13634_, _11862_, _13633_);
  and _65130_ (_13635_, _13495_, _13634_);
  not _65131_ (_13637_, _13635_);
  or _65132_ (_13638_, _13637_, _12043_);
  and _65133_ (_13639_, _13495_, _04797_);
  or _65134_ (_13640_, _13639_, \oc8051_golden_model_1.IRAM[7] [0]);
  and _65135_ (_13641_, _13500_, _04550_);
  not _65136_ (_13642_, _13641_);
  and _65137_ (_13643_, _13642_, _13640_);
  and _65138_ (_13644_, _13643_, _13638_);
  and _65139_ (_13645_, _13641_, _13404_);
  or _65140_ (_40648_, _13645_, _13644_);
  or _65141_ (_13647_, _13639_, \oc8051_golden_model_1.IRAM[7] [1]);
  and _65142_ (_13648_, _13647_, _13642_);
  not _65143_ (_13649_, _13639_);
  or _65144_ (_13650_, _13649_, _12255_);
  and _65145_ (_13651_, _13650_, _13648_);
  and _65146_ (_13652_, _13641_, _13412_);
  or _65147_ (_40650_, _13652_, _13651_);
  or _65148_ (_13653_, _13639_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _65149_ (_13654_, _13653_, _13642_);
  or _65150_ (_13655_, _13649_, _12459_);
  and _65151_ (_13657_, _13655_, _13654_);
  and _65152_ (_13658_, _13641_, _13418_);
  or _65153_ (_40651_, _13658_, _13657_);
  or _65154_ (_13659_, _13637_, _12661_);
  or _65155_ (_13660_, _13635_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _65156_ (_13661_, _13660_, _13642_);
  and _65157_ (_13662_, _13661_, _13659_);
  and _65158_ (_13663_, _13641_, _13424_);
  or _65159_ (_40652_, _13663_, _13662_);
  or _65160_ (_13664_, _13639_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _65161_ (_13666_, _13664_, _13642_);
  or _65162_ (_13667_, _13649_, _12896_);
  and _65163_ (_13668_, _13667_, _13666_);
  and _65164_ (_13669_, _13641_, _13430_);
  or _65165_ (_40653_, _13669_, _13668_);
  or _65166_ (_13670_, _13639_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _65167_ (_13671_, _13670_, _13642_);
  or _65168_ (_13672_, _13649_, _13100_);
  and _65169_ (_13673_, _13672_, _13671_);
  and _65170_ (_13674_, _13641_, _13436_);
  or _65171_ (_40654_, _13674_, _13673_);
  or _65172_ (_13676_, _13639_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _65173_ (_13677_, _13676_, _13642_);
  or _65174_ (_13678_, _13649_, _13315_);
  and _65175_ (_13679_, _13678_, _13677_);
  and _65176_ (_13680_, _13641_, _13442_);
  or _65177_ (_40656_, _13680_, _13679_);
  or _65178_ (_13681_, _13639_, \oc8051_golden_model_1.IRAM[7] [7]);
  and _65179_ (_13682_, _13681_, _13642_);
  or _65180_ (_13683_, _13649_, _06733_);
  and _65181_ (_13685_, _13683_, _13682_);
  and _65182_ (_13686_, _13641_, _06757_);
  or _65183_ (_40657_, _13686_, _13685_);
  and _65184_ (_13687_, _11864_, _05102_);
  and _65185_ (_13688_, _13687_, _11863_);
  not _65186_ (_13689_, _13688_);
  or _65187_ (_13690_, _13689_, _12043_);
  and _65188_ (_13691_, _05118_, _12674_);
  and _65189_ (_13692_, _13691_, _04551_);
  not _65190_ (_13693_, _13692_);
  or _65191_ (_13695_, _13688_, \oc8051_golden_model_1.IRAM[8] [0]);
  and _65192_ (_13696_, _13695_, _13693_);
  and _65193_ (_13697_, _13696_, _13690_);
  and _65194_ (_13698_, _13692_, _13404_);
  or _65195_ (_40661_, _13698_, _13697_);
  or _65196_ (_13699_, _13689_, _12255_);
  or _65197_ (_13700_, _13688_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _65198_ (_13701_, _13700_, _13693_);
  and _65199_ (_13702_, _13701_, _13699_);
  and _65200_ (_13703_, _13692_, _13412_);
  or _65201_ (_40662_, _13703_, _13702_);
  or _65202_ (_13705_, _13689_, _12459_);
  or _65203_ (_13706_, _13688_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _65204_ (_13707_, _13706_, _13693_);
  and _65205_ (_13708_, _13707_, _13705_);
  and _65206_ (_13709_, _13692_, _13418_);
  or _65207_ (_40663_, _13709_, _13708_);
  or _65208_ (_13710_, _13689_, _12661_);
  or _65209_ (_13711_, _13688_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _65210_ (_13712_, _13711_, _13693_);
  and _65211_ (_13714_, _13712_, _13710_);
  and _65212_ (_13715_, _13692_, _13424_);
  or _65213_ (_40665_, _13715_, _13714_);
  or _65214_ (_13716_, _13689_, _12896_);
  or _65215_ (_13717_, _13688_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _65216_ (_13718_, _13717_, _13693_);
  and _65217_ (_13719_, _13718_, _13716_);
  and _65218_ (_13720_, _13692_, _13430_);
  or _65219_ (_40666_, _13720_, _13719_);
  or _65220_ (_13721_, _13689_, _13100_);
  or _65221_ (_13723_, _13688_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _65222_ (_13724_, _13723_, _13693_);
  and _65223_ (_13725_, _13724_, _13721_);
  and _65224_ (_13726_, _13692_, _13436_);
  or _65225_ (_40667_, _13726_, _13725_);
  or _65226_ (_13727_, _13689_, _13315_);
  or _65227_ (_13728_, _13688_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _65228_ (_13729_, _13728_, _13693_);
  and _65229_ (_13730_, _13729_, _13727_);
  and _65230_ (_13731_, _13692_, _13442_);
  or _65231_ (_40668_, _13731_, _13730_);
  or _65232_ (_13732_, _13689_, _06733_);
  or _65233_ (_13733_, _13688_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _65234_ (_13734_, _13733_, _13693_);
  and _65235_ (_13735_, _13734_, _13732_);
  and _65236_ (_13736_, _13692_, _06757_);
  or _65237_ (_40669_, _13736_, _13735_);
  and _65238_ (_13737_, _13687_, _13334_);
  not _65239_ (_13738_, _13737_);
  nor _65240_ (_13739_, _13738_, _12043_);
  nor _65241_ (_13740_, _13737_, \oc8051_golden_model_1.IRAM[9] [0]);
  or _65242_ (_13741_, _13740_, _13739_);
  and _65243_ (_13742_, _13691_, _04845_);
  not _65244_ (_13743_, _13742_);
  nand _65245_ (_13744_, _13743_, _13741_);
  or _65246_ (_13745_, _13743_, _13404_);
  and _65247_ (_40673_, _13745_, _13744_);
  or _65248_ (_13746_, _13738_, _12255_);
  or _65249_ (_13747_, _13737_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _65250_ (_13748_, _13747_, _13743_);
  and _65251_ (_13749_, _13748_, _13746_);
  and _65252_ (_13750_, _13742_, _13412_);
  or _65253_ (_40674_, _13750_, _13749_);
  or _65254_ (_13751_, _13738_, _12459_);
  or _65255_ (_13752_, _13737_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _65256_ (_13753_, _13752_, _13743_);
  and _65257_ (_13754_, _13753_, _13751_);
  and _65258_ (_13755_, _13742_, _13418_);
  or _65259_ (_40676_, _13755_, _13754_);
  or _65260_ (_13756_, _13738_, _12661_);
  or _65261_ (_13757_, _13737_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _65262_ (_13758_, _13757_, _13743_);
  and _65263_ (_13759_, _13758_, _13756_);
  and _65264_ (_13760_, _13742_, _13424_);
  or _65265_ (_40677_, _13760_, _13759_);
  or _65266_ (_13761_, _13738_, _12896_);
  or _65267_ (_13762_, _13737_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _65268_ (_13763_, _13762_, _13743_);
  and _65269_ (_13764_, _13763_, _13761_);
  and _65270_ (_13765_, _13742_, _13430_);
  or _65271_ (_40678_, _13765_, _13764_);
  or _65272_ (_13766_, _13738_, _13100_);
  or _65273_ (_13767_, _13737_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _65274_ (_13768_, _13767_, _13743_);
  and _65275_ (_13769_, _13768_, _13766_);
  and _65276_ (_13770_, _13742_, _13436_);
  or _65277_ (_40679_, _13770_, _13769_);
  or _65278_ (_13771_, _13738_, _13315_);
  or _65279_ (_13772_, _13737_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _65280_ (_13773_, _13772_, _13743_);
  and _65281_ (_13774_, _13773_, _13771_);
  and _65282_ (_13775_, _13742_, _13442_);
  or _65283_ (_40680_, _13775_, _13774_);
  or _65284_ (_13776_, _13738_, _06733_);
  or _65285_ (_13777_, _13737_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _65286_ (_13778_, _13777_, _13743_);
  and _65287_ (_13779_, _13778_, _13776_);
  and _65288_ (_13780_, _13742_, _06757_);
  or _65289_ (_40682_, _13780_, _13779_);
  and _65290_ (_13781_, _13687_, _13392_);
  not _65291_ (_13782_, _13781_);
  or _65292_ (_13783_, _13782_, _12043_);
  or _65293_ (_13784_, _13781_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _65294_ (_13785_, _13691_, _05848_);
  not _65295_ (_13786_, _13785_);
  and _65296_ (_13787_, _13786_, _13784_);
  and _65297_ (_13788_, _13787_, _13783_);
  and _65298_ (_13789_, _13785_, _13404_);
  or _65299_ (_40685_, _13789_, _13788_);
  or _65300_ (_13790_, _13782_, _12255_);
  or _65301_ (_13791_, _13781_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _65302_ (_13792_, _13791_, _13786_);
  and _65303_ (_13793_, _13792_, _13790_);
  and _65304_ (_13794_, _13785_, _13412_);
  or _65305_ (_40686_, _13794_, _13793_);
  or _65306_ (_13795_, _13782_, _12459_);
  or _65307_ (_13796_, _13781_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _65308_ (_13797_, _13796_, _13786_);
  and _65309_ (_13798_, _13797_, _13795_);
  and _65310_ (_13799_, _13785_, _13418_);
  or _65311_ (_40688_, _13799_, _13798_);
  or _65312_ (_13800_, _13782_, _12661_);
  or _65313_ (_13801_, _13781_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _65314_ (_13802_, _13801_, _13786_);
  and _65315_ (_13803_, _13802_, _13800_);
  and _65316_ (_13804_, _13785_, _13424_);
  or _65317_ (_40689_, _13804_, _13803_);
  or _65318_ (_13805_, _13782_, _12896_);
  or _65319_ (_13806_, _13781_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _65320_ (_13807_, _13806_, _13786_);
  and _65321_ (_13808_, _13807_, _13805_);
  and _65322_ (_13809_, _13785_, _13430_);
  or _65323_ (_40690_, _13809_, _13808_);
  or _65324_ (_13810_, _13782_, _13100_);
  or _65325_ (_13811_, _13781_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _65326_ (_13812_, _13811_, _13786_);
  and _65327_ (_13813_, _13812_, _13810_);
  and _65328_ (_13814_, _13785_, _13436_);
  or _65329_ (_40691_, _13814_, _13813_);
  or _65330_ (_13815_, _13782_, _13315_);
  or _65331_ (_13816_, _13781_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _65332_ (_13817_, _13816_, _13786_);
  and _65333_ (_13818_, _13817_, _13815_);
  and _65334_ (_13819_, _13785_, _13442_);
  or _65335_ (_40692_, _13819_, _13818_);
  or _65336_ (_13820_, _13782_, _06733_);
  or _65337_ (_13821_, _13781_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _65338_ (_13822_, _13821_, _13786_);
  and _65339_ (_13823_, _13822_, _13820_);
  and _65340_ (_13824_, _13785_, _06757_);
  or _65341_ (_40694_, _13824_, _13823_);
  and _65342_ (_13825_, _13687_, _13634_);
  not _65343_ (_13826_, _13825_);
  or _65344_ (_13827_, _13826_, _12043_);
  or _65345_ (_13828_, _13825_, \oc8051_golden_model_1.IRAM[11] [0]);
  and _65346_ (_13829_, _13828_, _13827_);
  and _65347_ (_13830_, _13691_, _04550_);
  or _65348_ (_13831_, _13830_, _13829_);
  not _65349_ (_13832_, _13830_);
  or _65350_ (_13833_, _13832_, _13404_);
  and _65351_ (_40697_, _13833_, _13831_);
  and _65352_ (_13834_, _13687_, _04797_);
  or _65353_ (_13835_, _13834_, \oc8051_golden_model_1.IRAM[11] [1]);
  and _65354_ (_13836_, _13835_, _13832_);
  not _65355_ (_13837_, _13834_);
  or _65356_ (_13838_, _13837_, _12255_);
  and _65357_ (_13839_, _13838_, _13836_);
  and _65358_ (_13840_, _13830_, _13412_);
  or _65359_ (_40699_, _13840_, _13839_);
  or _65360_ (_13841_, _13834_, \oc8051_golden_model_1.IRAM[11] [2]);
  and _65361_ (_13842_, _13841_, _13832_);
  or _65362_ (_13843_, _13837_, _12459_);
  and _65363_ (_13844_, _13843_, _13842_);
  and _65364_ (_13845_, _13830_, _13418_);
  or _65365_ (_40700_, _13845_, _13844_);
  or _65366_ (_13846_, _13826_, _12661_);
  or _65367_ (_13847_, _13825_, \oc8051_golden_model_1.IRAM[11] [3]);
  and _65368_ (_13848_, _13847_, _13832_);
  and _65369_ (_13849_, _13848_, _13846_);
  and _65370_ (_13850_, _13830_, _13424_);
  or _65371_ (_40701_, _13850_, _13849_);
  or _65372_ (_13851_, _13834_, \oc8051_golden_model_1.IRAM[11] [4]);
  and _65373_ (_13852_, _13851_, _13832_);
  or _65374_ (_13853_, _13837_, _12896_);
  and _65375_ (_13854_, _13853_, _13852_);
  and _65376_ (_13855_, _13830_, _13430_);
  or _65377_ (_40702_, _13855_, _13854_);
  or _65378_ (_13856_, _13834_, \oc8051_golden_model_1.IRAM[11] [5]);
  and _65379_ (_13857_, _13856_, _13832_);
  or _65380_ (_13858_, _13837_, _13100_);
  and _65381_ (_13859_, _13858_, _13857_);
  and _65382_ (_13860_, _13830_, _13436_);
  or _65383_ (_40703_, _13860_, _13859_);
  or _65384_ (_13861_, _13834_, \oc8051_golden_model_1.IRAM[11] [6]);
  and _65385_ (_13862_, _13861_, _13832_);
  or _65386_ (_13863_, _13837_, _13315_);
  and _65387_ (_13864_, _13863_, _13862_);
  and _65388_ (_13865_, _13830_, _13442_);
  or _65389_ (_40705_, _13865_, _13864_);
  or _65390_ (_13866_, _13834_, \oc8051_golden_model_1.IRAM[11] [7]);
  and _65391_ (_13867_, _13866_, _13832_);
  or _65392_ (_13868_, _13837_, _06733_);
  and _65393_ (_13869_, _13868_, _13867_);
  and _65394_ (_13870_, _13830_, _06757_);
  or _65395_ (_40706_, _13870_, _13869_);
  and _65396_ (_13871_, _11863_, _05105_);
  nor _65397_ (_13872_, _13871_, \oc8051_golden_model_1.IRAM[12] [0]);
  not _65398_ (_13873_, _05102_);
  and _65399_ (_13874_, _11864_, _13873_);
  and _65400_ (_13875_, _11863_, _13874_);
  not _65401_ (_13876_, _13875_);
  nor _65402_ (_13877_, _13876_, _12043_);
  or _65403_ (_13878_, _13877_, _13872_);
  and _65404_ (_13879_, _05119_, _04551_);
  nor _65405_ (_13880_, _13879_, _13878_);
  and _65406_ (_13881_, _13879_, _13404_);
  or _65407_ (_40710_, _13881_, _13880_);
  not _65408_ (_13882_, _13879_);
  or _65409_ (_13883_, _13871_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _65410_ (_13884_, _13883_, _13882_);
  or _65411_ (_13885_, _13876_, _12255_);
  and _65412_ (_13886_, _13885_, _13884_);
  and _65413_ (_13887_, _13879_, _13412_);
  or _65414_ (_40711_, _13887_, _13886_);
  or _65415_ (_13888_, _13871_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _65416_ (_13889_, _13888_, _13882_);
  or _65417_ (_13890_, _13876_, _12459_);
  and _65418_ (_13891_, _13890_, _13889_);
  and _65419_ (_13892_, _13879_, _13418_);
  or _65420_ (_40712_, _13892_, _13891_);
  or _65421_ (_13893_, _13876_, _12661_);
  or _65422_ (_13894_, _13875_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _65423_ (_13895_, _13894_, _13882_);
  and _65424_ (_13896_, _13895_, _13893_);
  and _65425_ (_13897_, _13879_, _13424_);
  or _65426_ (_40713_, _13897_, _13896_);
  or _65427_ (_13898_, _13871_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _65428_ (_13899_, _13898_, _13882_);
  or _65429_ (_13900_, _13876_, _12896_);
  and _65430_ (_13901_, _13900_, _13899_);
  and _65431_ (_13902_, _13879_, _13430_);
  or _65432_ (_40714_, _13902_, _13901_);
  or _65433_ (_13903_, _13871_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _65434_ (_13904_, _13903_, _13882_);
  or _65435_ (_13905_, _13876_, _13100_);
  and _65436_ (_13906_, _13905_, _13904_);
  and _65437_ (_13907_, _13879_, _13436_);
  or _65438_ (_40716_, _13907_, _13906_);
  or _65439_ (_13908_, _13871_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _65440_ (_13909_, _13908_, _13882_);
  or _65441_ (_13910_, _13876_, _13315_);
  and _65442_ (_13911_, _13910_, _13909_);
  and _65443_ (_13912_, _13879_, _13442_);
  or _65444_ (_40717_, _13912_, _13911_);
  or _65445_ (_13913_, _13871_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _65446_ (_13914_, _13913_, _13882_);
  or _65447_ (_13915_, _13876_, _06733_);
  and _65448_ (_13916_, _13915_, _13914_);
  and _65449_ (_13917_, _13879_, _06757_);
  or _65450_ (_40718_, _13917_, _13916_);
  nand _65451_ (_13918_, _13334_, _13874_);
  or _65452_ (_13919_, _13918_, _12043_);
  and _65453_ (_13920_, _13334_, _05105_);
  or _65454_ (_13921_, _13920_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _65455_ (_13922_, _05119_, _04845_);
  not _65456_ (_13923_, _13922_);
  and _65457_ (_13924_, _13923_, _13921_);
  and _65458_ (_13925_, _13924_, _13919_);
  and _65459_ (_13926_, _13922_, _13404_);
  or _65460_ (_40722_, _13926_, _13925_);
  or _65461_ (_13927_, _13920_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _65462_ (_13928_, _13927_, _13923_);
  or _65463_ (_13929_, _13918_, _12255_);
  and _65464_ (_13930_, _13929_, _13928_);
  and _65465_ (_13931_, _13922_, _13412_);
  or _65466_ (_40723_, _13931_, _13930_);
  or _65467_ (_13932_, _13920_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _65468_ (_13933_, _13932_, _13923_);
  or _65469_ (_13934_, _13918_, _12459_);
  and _65470_ (_13935_, _13934_, _13933_);
  and _65471_ (_13936_, _13922_, _13418_);
  or _65472_ (_40724_, _13936_, _13935_);
  or _65473_ (_13937_, _13920_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _65474_ (_13938_, _13937_, _13923_);
  or _65475_ (_13939_, _13918_, _12661_);
  and _65476_ (_13940_, _13939_, _13938_);
  and _65477_ (_13941_, _13922_, _13424_);
  or _65478_ (_40725_, _13941_, _13940_);
  or _65479_ (_13942_, _13920_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _65480_ (_13943_, _13942_, _13923_);
  or _65481_ (_13944_, _13918_, _12896_);
  and _65482_ (_13945_, _13944_, _13943_);
  and _65483_ (_13946_, _13922_, _13430_);
  or _65484_ (_40727_, _13946_, _13945_);
  or _65485_ (_13947_, _13920_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _65486_ (_13948_, _13947_, _13923_);
  or _65487_ (_13949_, _13918_, _13100_);
  and _65488_ (_13950_, _13949_, _13948_);
  and _65489_ (_13951_, _13922_, _13436_);
  or _65490_ (_40728_, _13951_, _13950_);
  or _65491_ (_13952_, _13920_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _65492_ (_13953_, _13952_, _13923_);
  or _65493_ (_13954_, _13918_, _13315_);
  and _65494_ (_13955_, _13954_, _13953_);
  and _65495_ (_13956_, _13922_, _13442_);
  or _65496_ (_40729_, _13956_, _13955_);
  or _65497_ (_13957_, _13920_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _65498_ (_13958_, _13957_, _13923_);
  or _65499_ (_13959_, _13918_, _06733_);
  and _65500_ (_13960_, _13959_, _13958_);
  and _65501_ (_13961_, _13922_, _06757_);
  or _65502_ (_40730_, _13961_, _13960_);
  and _65503_ (_13962_, _13392_, _13874_);
  not _65504_ (_13963_, _13962_);
  or _65505_ (_13964_, _13963_, _12043_);
  and _65506_ (_13965_, _05848_, _05119_);
  not _65507_ (_13966_, _13965_);
  or _65508_ (_13967_, _13962_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _65509_ (_13968_, _13967_, _13966_);
  and _65510_ (_13969_, _13968_, _13964_);
  and _65511_ (_13970_, _13965_, _13404_);
  or _65512_ (_40734_, _13970_, _13969_);
  or _65513_ (_13971_, _13962_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _65514_ (_13972_, _13971_, _13966_);
  or _65515_ (_13973_, _13963_, _12255_);
  and _65516_ (_13974_, _13973_, _13972_);
  and _65517_ (_13975_, _13965_, _13412_);
  or _65518_ (_40735_, _13975_, _13974_);
  or _65519_ (_13976_, _13962_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _65520_ (_13977_, _13976_, _13966_);
  or _65521_ (_13978_, _13963_, _12459_);
  and _65522_ (_13979_, _13978_, _13977_);
  and _65523_ (_13980_, _13965_, _13418_);
  or _65524_ (_40736_, _13980_, _13979_);
  or _65525_ (_13981_, _13963_, _12661_);
  or _65526_ (_13982_, _13962_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _65527_ (_13983_, _13982_, _13966_);
  and _65528_ (_13984_, _13983_, _13981_);
  and _65529_ (_13985_, _13965_, _13424_);
  or _65530_ (_40737_, _13985_, _13984_);
  or _65531_ (_13986_, _13962_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _65532_ (_13987_, _13986_, _13966_);
  or _65533_ (_13988_, _13963_, _12896_);
  and _65534_ (_13989_, _13988_, _13987_);
  and _65535_ (_13990_, _13965_, _13430_);
  or _65536_ (_40739_, _13990_, _13989_);
  or _65537_ (_13991_, _13962_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _65538_ (_13992_, _13991_, _13966_);
  or _65539_ (_13993_, _13963_, _13100_);
  and _65540_ (_13994_, _13993_, _13992_);
  and _65541_ (_13995_, _13965_, _13436_);
  or _65542_ (_40740_, _13995_, _13994_);
  or _65543_ (_13996_, _13962_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _65544_ (_13997_, _13996_, _13966_);
  or _65545_ (_13998_, _13963_, _13315_);
  and _65546_ (_13999_, _13998_, _13997_);
  and _65547_ (_14000_, _13965_, _13442_);
  or _65548_ (_40741_, _14000_, _13999_);
  or _65549_ (_14001_, _13962_, \oc8051_golden_model_1.IRAM[14] [7]);
  and _65550_ (_14002_, _14001_, _13966_);
  or _65551_ (_14003_, _13963_, _06733_);
  and _65552_ (_14004_, _14003_, _14002_);
  and _65553_ (_14005_, _13965_, _06757_);
  or _65554_ (_40742_, _14005_, _14004_);
  and _65555_ (_14006_, _13874_, _13634_);
  not _65556_ (_14007_, _14006_);
  or _65557_ (_14008_, _12043_, _14007_);
  or _65558_ (_14009_, _14006_, \oc8051_golden_model_1.IRAM[15] [0]);
  and _65559_ (_14010_, _14009_, _14008_);
  or _65560_ (_14011_, _14010_, _05120_);
  or _65561_ (_14012_, _13404_, _05121_);
  and _65562_ (_40746_, _14012_, _14011_);
  or _65563_ (_14013_, _05106_, \oc8051_golden_model_1.IRAM[15] [1]);
  and _65564_ (_14014_, _14013_, _05121_);
  or _65565_ (_14015_, _12255_, _05123_);
  and _65566_ (_14016_, _14015_, _14014_);
  and _65567_ (_14017_, _13412_, _05120_);
  or _65568_ (_40747_, _14017_, _14016_);
  or _65569_ (_14018_, _05106_, \oc8051_golden_model_1.IRAM[15] [2]);
  and _65570_ (_14019_, _14018_, _05121_);
  or _65571_ (_14020_, _12459_, _05123_);
  and _65572_ (_14021_, _14020_, _14019_);
  and _65573_ (_14022_, _13418_, _05120_);
  or _65574_ (_40748_, _14022_, _14021_);
  or _65575_ (_14023_, _12661_, _14007_);
  or _65576_ (_14024_, _14006_, \oc8051_golden_model_1.IRAM[15] [3]);
  and _65577_ (_14025_, _14024_, _05121_);
  and _65578_ (_14026_, _14025_, _14023_);
  and _65579_ (_14027_, _13424_, _05120_);
  or _65580_ (_40749_, _14027_, _14026_);
  or _65581_ (_14028_, _05106_, \oc8051_golden_model_1.IRAM[15] [4]);
  and _65582_ (_14029_, _14028_, _05121_);
  or _65583_ (_14030_, _12896_, _05123_);
  and _65584_ (_14031_, _14030_, _14029_);
  and _65585_ (_14032_, _13430_, _05120_);
  or _65586_ (_40751_, _14032_, _14031_);
  or _65587_ (_14033_, _05106_, \oc8051_golden_model_1.IRAM[15] [5]);
  and _65588_ (_14034_, _14033_, _05121_);
  or _65589_ (_14035_, _13100_, _05123_);
  and _65590_ (_14036_, _14035_, _14034_);
  and _65591_ (_14037_, _13436_, _05120_);
  or _65592_ (_40752_, _14037_, _14036_);
  or _65593_ (_14038_, _05106_, \oc8051_golden_model_1.IRAM[15] [6]);
  and _65594_ (_14039_, _14038_, _05121_);
  or _65595_ (_14040_, _13315_, _05123_);
  and _65596_ (_14041_, _14040_, _14039_);
  and _65597_ (_14042_, _13442_, _05120_);
  or _65598_ (_40753_, _14042_, _14041_);
  nor _65599_ (_14043_, _42963_, _07340_);
  nor _65600_ (_14044_, _05221_, _07340_);
  and _65601_ (_14045_, _11995_, _05221_);
  or _65602_ (_14046_, _14045_, _14044_);
  and _65603_ (_14047_, _14046_, _03769_);
  and _65604_ (_14048_, _05221_, _06202_);
  or _65605_ (_14049_, _14048_, _14044_);
  or _65606_ (_14050_, _14049_, _03438_);
  and _65607_ (_14051_, _05221_, _04419_);
  or _65608_ (_14052_, _14051_, _14044_);
  or _65609_ (_14053_, _14052_, _06039_);
  and _65610_ (_14054_, _05941_, _05221_);
  or _65611_ (_14055_, _14054_, _14044_);
  and _65612_ (_14056_, _14055_, _03570_);
  nor _65613_ (_14057_, _04426_, _07340_);
  and _65614_ (_14058_, _05221_, \oc8051_golden_model_1.ACC [0]);
  or _65615_ (_14059_, _14058_, _14044_);
  and _65616_ (_14060_, _14059_, _04426_);
  or _65617_ (_14061_, _14060_, _14057_);
  and _65618_ (_14062_, _14061_, _04444_);
  or _65619_ (_14063_, _14062_, _03516_);
  or _65620_ (_14064_, _14063_, _14056_);
  and _65621_ (_14065_, _11887_, _05785_);
  nor _65622_ (_14066_, _05785_, _07340_);
  or _65623_ (_14067_, _14066_, _14065_);
  or _65624_ (_14068_, _14067_, _03517_);
  and _65625_ (_14069_, _14068_, _14064_);
  or _65626_ (_14070_, _14069_, _03568_);
  or _65627_ (_14071_, _14052_, _03983_);
  and _65628_ (_14072_, _14071_, _14070_);
  or _65629_ (_14073_, _14072_, _03575_);
  or _65630_ (_14074_, _14059_, _03583_);
  and _65631_ (_14075_, _14074_, _03513_);
  and _65632_ (_14076_, _14075_, _14073_);
  and _65633_ (_14077_, _14044_, _03512_);
  or _65634_ (_14078_, _14077_, _03505_);
  or _65635_ (_14079_, _14078_, _14076_);
  or _65636_ (_14080_, _14055_, _03506_);
  and _65637_ (_14081_, _14080_, _14079_);
  or _65638_ (_14082_, _14081_, _06794_);
  nor _65639_ (_14083_, _07287_, _07285_);
  nor _65640_ (_14084_, _14083_, _07288_);
  or _65641_ (_14085_, _14084_, _06800_);
  and _65642_ (_14086_, _14085_, _03500_);
  and _65643_ (_14087_, _14086_, _14082_);
  nor _65644_ (_14088_, _11916_, _07315_);
  or _65645_ (_14089_, _14088_, _14066_);
  and _65646_ (_14090_, _14089_, _03499_);
  or _65647_ (_14091_, _14090_, _07314_);
  or _65648_ (_14092_, _14091_, _14087_);
  and _65649_ (_14093_, _14092_, _14053_);
  or _65650_ (_14094_, _14093_, _03479_);
  and _65651_ (_14095_, _06715_, _05221_);
  or _65652_ (_14096_, _14044_, _06044_);
  or _65653_ (_14097_, _14096_, _14095_);
  and _65654_ (_14098_, _14097_, _14094_);
  or _65655_ (_14099_, _14098_, _03221_);
  nor _65656_ (_14100_, _11975_, _06762_);
  or _65657_ (_14101_, _14044_, _03474_);
  or _65658_ (_14102_, _14101_, _14100_);
  and _65659_ (_14103_, _14102_, _07677_);
  and _65660_ (_14104_, _14103_, _14099_);
  nand _65661_ (_14105_, _07675_, _03321_);
  nor _65662_ (_14106_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor _65663_ (_14107_, _14106_, _07266_);
  or _65664_ (_14108_, _07675_, _14107_);
  and _65665_ (_14109_, _14108_, _07328_);
  and _65666_ (_14110_, _14109_, _14105_);
  or _65667_ (_14111_, _14110_, _03437_);
  or _65668_ (_14112_, _14111_, _14104_);
  and _65669_ (_14113_, _14112_, _14050_);
  or _65670_ (_14114_, _14113_, _03636_);
  and _65671_ (_14115_, _11990_, _05221_);
  or _65672_ (_14116_, _14115_, _14044_);
  or _65673_ (_14117_, _14116_, _04499_);
  and _65674_ (_14118_, _14117_, _04501_);
  and _65675_ (_14119_, _14118_, _14114_);
  or _65676_ (_14120_, _14119_, _14047_);
  and _65677_ (_14121_, _14120_, _05769_);
  nand _65678_ (_14122_, _14049_, _03754_);
  nor _65679_ (_14123_, _14122_, _14054_);
  or _65680_ (_14124_, _14123_, _14121_);
  and _65681_ (_14125_, _14124_, _03753_);
  or _65682_ (_14126_, _14044_, _05617_);
  and _65683_ (_14127_, _14059_, _03752_);
  and _65684_ (_14128_, _14127_, _14126_);
  or _65685_ (_14129_, _14128_, _03758_);
  or _65686_ (_14130_, _14129_, _14125_);
  nor _65687_ (_14131_, _11988_, _06762_);
  or _65688_ (_14132_, _14044_, _03759_);
  or _65689_ (_14133_, _14132_, _14131_);
  and _65690_ (_14134_, _14133_, _04517_);
  and _65691_ (_14135_, _14134_, _14130_);
  nor _65692_ (_14136_, _11870_, _06762_);
  or _65693_ (_14137_, _14136_, _14044_);
  and _65694_ (_14138_, _14137_, _03760_);
  or _65695_ (_14139_, _14138_, _03790_);
  or _65696_ (_14140_, _14139_, _14135_);
  or _65697_ (_14141_, _14055_, _04192_);
  and _65698_ (_14142_, _14141_, _03152_);
  and _65699_ (_14143_, _14142_, _14140_);
  and _65700_ (_14144_, _14044_, _03151_);
  or _65701_ (_14145_, _14144_, _03520_);
  or _65702_ (_14146_, _14145_, _14143_);
  or _65703_ (_14147_, _14055_, _03521_);
  and _65704_ (_14148_, _14147_, _42963_);
  and _65705_ (_14149_, _14148_, _14146_);
  or _65706_ (_14150_, _14149_, _14043_);
  and _65707_ (_43194_, _14150_, _41755_);
  nor _65708_ (_14151_, _42963_, _07334_);
  or _65709_ (_14152_, _05221_, \oc8051_golden_model_1.B [1]);
  and _65710_ (_14153_, _12252_, _05221_);
  not _65711_ (_14154_, _14153_);
  and _65712_ (_14155_, _14154_, _14152_);
  or _65713_ (_14156_, _14155_, _04444_);
  nand _65714_ (_14157_, _05221_, _03233_);
  and _65715_ (_14158_, _14157_, _14152_);
  and _65716_ (_14159_, _14158_, _04426_);
  nor _65717_ (_14160_, _04426_, _07334_);
  or _65718_ (_14161_, _14160_, _03570_);
  or _65719_ (_14162_, _14161_, _14159_);
  and _65720_ (_14163_, _14162_, _03517_);
  and _65721_ (_14164_, _14163_, _14156_);
  not _65722_ (_14165_, _03576_);
  and _65723_ (_14166_, _12083_, _05785_);
  nor _65724_ (_14167_, _05785_, _07334_);
  or _65725_ (_14168_, _14167_, _03568_);
  or _65726_ (_14169_, _14168_, _14166_);
  and _65727_ (_14170_, _14169_, _14165_);
  or _65728_ (_14171_, _14170_, _14164_);
  nor _65729_ (_14172_, _05221_, _07334_);
  nor _65730_ (_14173_, _06762_, _04603_);
  or _65731_ (_14174_, _14173_, _14172_);
  or _65732_ (_14175_, _14174_, _03983_);
  and _65733_ (_14176_, _14175_, _14171_);
  or _65734_ (_14177_, _14176_, _03575_);
  or _65735_ (_14178_, _14158_, _03583_);
  and _65736_ (_14179_, _14178_, _03513_);
  and _65737_ (_14180_, _14179_, _14177_);
  and _65738_ (_14181_, _12069_, _05785_);
  or _65739_ (_14182_, _14181_, _14167_);
  and _65740_ (_14183_, _14182_, _03512_);
  or _65741_ (_14184_, _14183_, _14180_);
  and _65742_ (_14185_, _14184_, _03506_);
  and _65743_ (_14186_, _14166_, _12098_);
  or _65744_ (_14187_, _14186_, _14167_);
  and _65745_ (_14188_, _14187_, _03505_);
  or _65746_ (_14189_, _14188_, _06794_);
  or _65747_ (_14190_, _14189_, _14185_);
  nor _65748_ (_14191_, _07290_, _07233_);
  nor _65749_ (_14192_, _14191_, _07291_);
  or _65750_ (_14193_, _14192_, _06800_);
  and _65751_ (_14194_, _14193_, _03500_);
  and _65752_ (_14195_, _14194_, _14190_);
  nor _65753_ (_14196_, _12116_, _07315_);
  or _65754_ (_14197_, _14196_, _14167_);
  and _65755_ (_14198_, _14197_, _03499_);
  or _65756_ (_14199_, _14198_, _07314_);
  or _65757_ (_14200_, _14199_, _14195_);
  or _65758_ (_14201_, _14174_, _06039_);
  and _65759_ (_14202_, _14201_, _14200_);
  or _65760_ (_14203_, _14202_, _03479_);
  and _65761_ (_14204_, _06714_, _05221_);
  or _65762_ (_14205_, _14172_, _06044_);
  or _65763_ (_14206_, _14205_, _14204_);
  and _65764_ (_14207_, _14206_, _03474_);
  and _65765_ (_14208_, _14207_, _14203_);
  nand _65766_ (_14209_, _12176_, _05221_);
  and _65767_ (_14210_, _14152_, _03221_);
  and _65768_ (_14211_, _14210_, _14209_);
  or _65769_ (_14212_, _14211_, _07328_);
  or _65770_ (_14213_, _14212_, _14208_);
  and _65771_ (_14214_, _07675_, _07641_);
  nor _65772_ (_14215_, _07670_, _07669_);
  or _65773_ (_14216_, _14215_, _07671_);
  nor _65774_ (_14217_, _14216_, _07675_);
  or _65775_ (_14218_, _14217_, _14214_);
  or _65776_ (_14219_, _14218_, _07677_);
  and _65777_ (_14220_, _14219_, _03438_);
  and _65778_ (_14221_, _14220_, _14213_);
  nand _65779_ (_14222_, _05221_, _04317_);
  and _65780_ (_14223_, _14152_, _03437_);
  and _65781_ (_14224_, _14223_, _14222_);
  or _65782_ (_14225_, _14224_, _14221_);
  and _65783_ (_14226_, _14225_, _04499_);
  or _65784_ (_14227_, _12191_, _06762_);
  and _65785_ (_14228_, _14152_, _03636_);
  and _65786_ (_14229_, _14228_, _14227_);
  or _65787_ (_14230_, _14229_, _14226_);
  and _65788_ (_14231_, _14230_, _04501_);
  or _65789_ (_14232_, _12197_, _06762_);
  and _65790_ (_14233_, _14152_, _03769_);
  and _65791_ (_14234_, _14233_, _14232_);
  or _65792_ (_14235_, _14234_, _14231_);
  and _65793_ (_14236_, _14235_, _05769_);
  or _65794_ (_14237_, _12190_, _06762_);
  and _65795_ (_14238_, _14237_, _03754_);
  and _65796_ (_14239_, _14238_, _14152_);
  or _65797_ (_14240_, _14239_, _14236_);
  and _65798_ (_14241_, _14240_, _03753_);
  or _65799_ (_14242_, _14172_, _05569_);
  and _65800_ (_14243_, _14158_, _03752_);
  and _65801_ (_14244_, _14243_, _14242_);
  or _65802_ (_14245_, _14244_, _14241_);
  and _65803_ (_14246_, _14245_, _03759_);
  or _65804_ (_14247_, _14222_, _05569_);
  and _65805_ (_14248_, _14152_, _03758_);
  and _65806_ (_14249_, _14248_, _14247_);
  or _65807_ (_14250_, _14249_, _14246_);
  and _65808_ (_14251_, _14250_, _04517_);
  nand _65809_ (_14252_, _12196_, _05221_);
  and _65810_ (_14253_, _14252_, _03760_);
  and _65811_ (_14254_, _14253_, _14152_);
  or _65812_ (_14255_, _14254_, _03790_);
  or _65813_ (_14256_, _14255_, _14251_);
  or _65814_ (_14257_, _14155_, _04192_);
  and _65815_ (_14258_, _14257_, _03152_);
  and _65816_ (_14259_, _14258_, _14256_);
  and _65817_ (_14260_, _14182_, _03151_);
  or _65818_ (_14261_, _14260_, _03520_);
  or _65819_ (_14262_, _14261_, _14259_);
  or _65820_ (_14263_, _14172_, _03521_);
  or _65821_ (_14264_, _14263_, _14153_);
  and _65822_ (_14265_, _14264_, _42963_);
  and _65823_ (_14266_, _14265_, _14262_);
  or _65824_ (_14267_, _14266_, _14151_);
  and _65825_ (_43195_, _14267_, _41755_);
  nor _65826_ (_14268_, _42963_, _07388_);
  nor _65827_ (_14269_, _05221_, _07388_);
  and _65828_ (_14270_, _12401_, _05221_);
  or _65829_ (_14271_, _14270_, _14269_);
  and _65830_ (_14272_, _14271_, _03769_);
  and _65831_ (_14273_, _05221_, _06261_);
  or _65832_ (_14274_, _14273_, _14269_);
  or _65833_ (_14275_, _14274_, _03438_);
  nor _65834_ (_14276_, _06762_, _05026_);
  or _65835_ (_14277_, _14276_, _14269_);
  or _65836_ (_14278_, _14277_, _06039_);
  and _65837_ (_14279_, _12278_, _05785_);
  and _65838_ (_14280_, _14279_, _12309_);
  nor _65839_ (_14281_, _05785_, _07388_);
  or _65840_ (_14282_, _14281_, _03506_);
  or _65841_ (_14283_, _14282_, _14280_);
  or _65842_ (_14284_, _14277_, _03983_);
  nor _65843_ (_14285_, _12282_, _06762_);
  or _65844_ (_14286_, _14285_, _14269_);
  or _65845_ (_14287_, _14286_, _04444_);
  and _65846_ (_14288_, _05221_, \oc8051_golden_model_1.ACC [2]);
  or _65847_ (_14289_, _14288_, _14269_);
  and _65848_ (_14290_, _14289_, _04426_);
  nor _65849_ (_14291_, _04426_, _07388_);
  or _65850_ (_14292_, _14291_, _03570_);
  or _65851_ (_14293_, _14292_, _14290_);
  and _65852_ (_14294_, _14293_, _03517_);
  and _65853_ (_14295_, _14294_, _14287_);
  or _65854_ (_14296_, _14281_, _14279_);
  and _65855_ (_14297_, _14296_, _03516_);
  or _65856_ (_14298_, _14297_, _03568_);
  or _65857_ (_14299_, _14298_, _14295_);
  and _65858_ (_14300_, _14299_, _14284_);
  or _65859_ (_14301_, _14300_, _03575_);
  or _65860_ (_14302_, _14289_, _03583_);
  and _65861_ (_14303_, _14302_, _03513_);
  and _65862_ (_14304_, _14303_, _14301_);
  and _65863_ (_14305_, _12276_, _05785_);
  or _65864_ (_14306_, _14305_, _14281_);
  and _65865_ (_14307_, _14306_, _03512_);
  or _65866_ (_14308_, _14307_, _03505_);
  or _65867_ (_14309_, _14308_, _14304_);
  and _65868_ (_14310_, _14309_, _14283_);
  or _65869_ (_14311_, _14310_, _06794_);
  or _65870_ (_14312_, _07292_, _07188_);
  and _65871_ (_14313_, _14312_, _07293_);
  or _65872_ (_14314_, _14313_, _06800_);
  and _65873_ (_14315_, _14314_, _03500_);
  and _65874_ (_14316_, _14315_, _14311_);
  nor _65875_ (_14317_, _12326_, _07315_);
  or _65876_ (_14318_, _14317_, _14281_);
  and _65877_ (_14319_, _14318_, _03499_);
  or _65878_ (_14320_, _14319_, _07314_);
  or _65879_ (_14321_, _14320_, _14316_);
  and _65880_ (_14322_, _14321_, _14278_);
  or _65881_ (_14323_, _14322_, _03479_);
  and _65882_ (_14324_, _06718_, _05221_);
  or _65883_ (_14325_, _14269_, _06044_);
  or _65884_ (_14326_, _14325_, _14324_);
  and _65885_ (_14327_, _14326_, _14323_);
  or _65886_ (_14328_, _14327_, _03221_);
  nor _65887_ (_14329_, _12384_, _06762_);
  or _65888_ (_14330_, _14269_, _03474_);
  or _65889_ (_14331_, _14330_, _14329_);
  and _65890_ (_14332_, _14331_, _07677_);
  and _65891_ (_14333_, _14332_, _14328_);
  nor _65892_ (_14334_, _07671_, _07642_);
  not _65893_ (_14335_, _14334_);
  and _65894_ (_14336_, _14335_, _07634_);
  nor _65895_ (_14337_, _14335_, _07634_);
  nor _65896_ (_14338_, _14337_, _14336_);
  or _65897_ (_14339_, _14338_, _07675_);
  not _65898_ (_14340_, _07675_);
  or _65899_ (_14341_, _14340_, _07631_);
  and _65900_ (_14342_, _14341_, _07328_);
  and _65901_ (_14343_, _14342_, _14339_);
  or _65902_ (_14344_, _14343_, _03437_);
  or _65903_ (_14345_, _14344_, _14333_);
  and _65904_ (_14346_, _14345_, _14275_);
  or _65905_ (_14347_, _14346_, _03636_);
  and _65906_ (_14348_, _12273_, _05221_);
  or _65907_ (_14349_, _14348_, _14269_);
  or _65908_ (_14350_, _14349_, _04499_);
  and _65909_ (_14351_, _14350_, _04501_);
  and _65910_ (_14352_, _14351_, _14347_);
  or _65911_ (_14353_, _14352_, _14272_);
  and _65912_ (_14354_, _14353_, _05769_);
  or _65913_ (_14355_, _14269_, _05665_);
  and _65914_ (_14356_, _14355_, _03754_);
  and _65915_ (_14357_, _14356_, _14274_);
  or _65916_ (_14358_, _14357_, _14354_);
  and _65917_ (_14359_, _14358_, _03753_);
  and _65918_ (_14360_, _14289_, _03752_);
  and _65919_ (_14361_, _14360_, _14355_);
  or _65920_ (_14362_, _14361_, _03758_);
  or _65921_ (_14363_, _14362_, _14359_);
  nor _65922_ (_14364_, _12272_, _06762_);
  or _65923_ (_14365_, _14269_, _03759_);
  or _65924_ (_14366_, _14365_, _14364_);
  and _65925_ (_14367_, _14366_, _04517_);
  and _65926_ (_14368_, _14367_, _14363_);
  nor _65927_ (_14369_, _12400_, _06762_);
  or _65928_ (_14370_, _14369_, _14269_);
  and _65929_ (_14371_, _14370_, _03760_);
  or _65930_ (_14372_, _14371_, _03790_);
  or _65931_ (_14373_, _14372_, _14368_);
  or _65932_ (_14374_, _14286_, _04192_);
  and _65933_ (_14375_, _14374_, _03152_);
  and _65934_ (_14376_, _14375_, _14373_);
  and _65935_ (_14377_, _14306_, _03151_);
  or _65936_ (_14378_, _14377_, _03520_);
  or _65937_ (_14379_, _14378_, _14376_);
  and _65938_ (_14380_, _12456_, _05221_);
  or _65939_ (_14381_, _14269_, _03521_);
  or _65940_ (_14382_, _14381_, _14380_);
  and _65941_ (_14383_, _14382_, _42963_);
  and _65942_ (_14384_, _14383_, _14379_);
  or _65943_ (_14385_, _14384_, _14268_);
  and _65944_ (_43196_, _14385_, _41755_);
  nor _65945_ (_14386_, _42963_, _07374_);
  nor _65946_ (_14387_, _05221_, _07374_);
  and _65947_ (_14388_, _12604_, _05221_);
  or _65948_ (_14389_, _14388_, _14387_);
  and _65949_ (_14390_, _14389_, _03769_);
  and _65950_ (_14391_, _05221_, _06217_);
  or _65951_ (_14392_, _14391_, _14387_);
  or _65952_ (_14393_, _14392_, _03438_);
  nor _65953_ (_14394_, _06762_, _04843_);
  or _65954_ (_14395_, _14394_, _14387_);
  or _65955_ (_14396_, _14395_, _06039_);
  nor _65956_ (_14397_, _05785_, _07374_);
  and _65957_ (_14398_, _12490_, _05785_);
  or _65958_ (_14399_, _14398_, _14397_);
  or _65959_ (_14400_, _14397_, _12507_);
  and _65960_ (_14401_, _14400_, _14399_);
  or _65961_ (_14402_, _14401_, _03506_);
  nor _65962_ (_14403_, _12486_, _06762_);
  or _65963_ (_14404_, _14403_, _14387_);
  or _65964_ (_14405_, _14404_, _04444_);
  and _65965_ (_14406_, _05221_, \oc8051_golden_model_1.ACC [3]);
  or _65966_ (_14407_, _14406_, _14387_);
  and _65967_ (_14408_, _14407_, _04426_);
  nor _65968_ (_14409_, _04426_, _07374_);
  or _65969_ (_14410_, _14409_, _03570_);
  or _65970_ (_14411_, _14410_, _14408_);
  and _65971_ (_14412_, _14411_, _03517_);
  and _65972_ (_14413_, _14412_, _14405_);
  and _65973_ (_14414_, _14399_, _03516_);
  or _65974_ (_14415_, _14414_, _03568_);
  or _65975_ (_14416_, _14415_, _14413_);
  or _65976_ (_14417_, _14395_, _03983_);
  and _65977_ (_14418_, _14417_, _14416_);
  or _65978_ (_14419_, _14418_, _03575_);
  or _65979_ (_14420_, _14407_, _03583_);
  and _65980_ (_14421_, _14420_, _03513_);
  and _65981_ (_14422_, _14421_, _14419_);
  and _65982_ (_14423_, _12500_, _05785_);
  or _65983_ (_14424_, _14423_, _14397_);
  and _65984_ (_14425_, _14424_, _03512_);
  or _65985_ (_14426_, _14425_, _03505_);
  or _65986_ (_14427_, _14426_, _14422_);
  and _65987_ (_14428_, _14427_, _14402_);
  or _65988_ (_14429_, _14428_, _06794_);
  nor _65989_ (_14430_, _07295_, _07130_);
  nor _65990_ (_14431_, _14430_, _07296_);
  or _65991_ (_14432_, _14431_, _06800_);
  and _65992_ (_14433_, _14432_, _03500_);
  and _65993_ (_14434_, _14433_, _14429_);
  nor _65994_ (_14435_, _12525_, _07315_);
  or _65995_ (_14436_, _14435_, _14397_);
  and _65996_ (_14437_, _14436_, _03499_);
  or _65997_ (_14438_, _14437_, _07314_);
  or _65998_ (_14439_, _14438_, _14434_);
  and _65999_ (_14440_, _14439_, _14396_);
  or _66000_ (_14441_, _14440_, _03479_);
  and _66001_ (_14442_, _06717_, _05221_);
  or _66002_ (_14443_, _14387_, _06044_);
  or _66003_ (_14444_, _14443_, _14442_);
  and _66004_ (_14445_, _14444_, _14441_);
  or _66005_ (_14446_, _14445_, _03221_);
  nor _66006_ (_14447_, _12583_, _06762_);
  or _66007_ (_14448_, _14387_, _03474_);
  or _66008_ (_14449_, _14448_, _14447_);
  and _66009_ (_14450_, _14449_, _07677_);
  and _66010_ (_14451_, _14450_, _14446_);
  nor _66011_ (_14452_, _14336_, _07633_);
  nor _66012_ (_14453_, _14452_, _07626_);
  and _66013_ (_14454_, _14452_, _07626_);
  or _66014_ (_14455_, _14454_, _14453_);
  or _66015_ (_14456_, _14455_, _07675_);
  or _66016_ (_14457_, _14340_, _07623_);
  and _66017_ (_14458_, _14457_, _07328_);
  and _66018_ (_14459_, _14458_, _14456_);
  or _66019_ (_14460_, _14459_, _03437_);
  or _66020_ (_14461_, _14460_, _14451_);
  and _66021_ (_14462_, _14461_, _14393_);
  or _66022_ (_14463_, _14462_, _03636_);
  and _66023_ (_14464_, _12598_, _05221_);
  or _66024_ (_14465_, _14464_, _14387_);
  or _66025_ (_14466_, _14465_, _04499_);
  and _66026_ (_14467_, _14466_, _04501_);
  and _66027_ (_14468_, _14467_, _14463_);
  or _66028_ (_14469_, _14468_, _14390_);
  and _66029_ (_14470_, _14469_, _05769_);
  or _66030_ (_14471_, _14387_, _05521_);
  and _66031_ (_14472_, _14471_, _03754_);
  and _66032_ (_14473_, _14472_, _14392_);
  or _66033_ (_14474_, _14473_, _14470_);
  and _66034_ (_14475_, _14474_, _03753_);
  and _66035_ (_14476_, _14407_, _03752_);
  and _66036_ (_14477_, _14476_, _14471_);
  or _66037_ (_14478_, _14477_, _03758_);
  or _66038_ (_14479_, _14478_, _14475_);
  nor _66039_ (_14480_, _12597_, _06762_);
  or _66040_ (_14481_, _14387_, _03759_);
  or _66041_ (_14482_, _14481_, _14480_);
  and _66042_ (_14483_, _14482_, _04517_);
  and _66043_ (_14484_, _14483_, _14479_);
  nor _66044_ (_14485_, _12603_, _06762_);
  or _66045_ (_14486_, _14485_, _14387_);
  and _66046_ (_14487_, _14486_, _03760_);
  or _66047_ (_14488_, _14487_, _03790_);
  or _66048_ (_14489_, _14488_, _14484_);
  or _66049_ (_14490_, _14404_, _04192_);
  and _66050_ (_14491_, _14490_, _03152_);
  and _66051_ (_14492_, _14491_, _14489_);
  and _66052_ (_14493_, _14424_, _03151_);
  or _66053_ (_14494_, _14493_, _03520_);
  or _66054_ (_14495_, _14494_, _14492_);
  and _66055_ (_14496_, _12658_, _05221_);
  or _66056_ (_14497_, _14387_, _03521_);
  or _66057_ (_14498_, _14497_, _14496_);
  and _66058_ (_14499_, _14498_, _42963_);
  and _66059_ (_14500_, _14499_, _14495_);
  or _66060_ (_14501_, _14500_, _14386_);
  and _66061_ (_43198_, _14501_, _41755_);
  nor _66062_ (_14502_, _42963_, _07472_);
  nor _66063_ (_14503_, _05221_, _07472_);
  and _66064_ (_14504_, _12844_, _05221_);
  or _66065_ (_14505_, _14504_, _14503_);
  and _66066_ (_14506_, _14505_, _03769_);
  and _66067_ (_14507_, _06233_, _05221_);
  or _66068_ (_14508_, _14507_, _14503_);
  or _66069_ (_14509_, _14508_, _03438_);
  nor _66070_ (_14510_, _12827_, _06762_);
  or _66071_ (_14511_, _14510_, _14503_);
  and _66072_ (_14512_, _14511_, _03221_);
  nor _66073_ (_14513_, _05785_, _07472_);
  and _66074_ (_14514_, _12718_, _05785_);
  or _66075_ (_14515_, _14514_, _14513_);
  and _66076_ (_14516_, _14515_, _03512_);
  nor _66077_ (_14517_, _12733_, _06762_);
  or _66078_ (_14518_, _14517_, _14503_);
  or _66079_ (_14519_, _14518_, _04444_);
  and _66080_ (_14520_, _05221_, \oc8051_golden_model_1.ACC [4]);
  or _66081_ (_14521_, _14520_, _14503_);
  and _66082_ (_14522_, _14521_, _04426_);
  nor _66083_ (_14523_, _04426_, _07472_);
  or _66084_ (_14524_, _14523_, _03570_);
  or _66085_ (_14525_, _14524_, _14522_);
  and _66086_ (_14526_, _14525_, _03517_);
  and _66087_ (_14527_, _14526_, _14519_);
  and _66088_ (_14528_, _12737_, _05785_);
  or _66089_ (_14529_, _14528_, _14513_);
  and _66090_ (_14530_, _14529_, _03516_);
  or _66091_ (_14531_, _14530_, _03568_);
  or _66092_ (_14532_, _14531_, _14527_);
  nor _66093_ (_14533_, _05712_, _06762_);
  or _66094_ (_14534_, _14533_, _14503_);
  or _66095_ (_14535_, _14534_, _03983_);
  and _66096_ (_14536_, _14535_, _14532_);
  or _66097_ (_14537_, _14536_, _03575_);
  or _66098_ (_14538_, _14521_, _03583_);
  and _66099_ (_14539_, _14538_, _03513_);
  and _66100_ (_14540_, _14539_, _14537_);
  or _66101_ (_14541_, _14540_, _14516_);
  and _66102_ (_14542_, _14541_, _03506_);
  or _66103_ (_14543_, _14513_, _12752_);
  and _66104_ (_14544_, _14543_, _03505_);
  and _66105_ (_14545_, _14544_, _14529_);
  or _66106_ (_14546_, _14545_, _06794_);
  or _66107_ (_14547_, _14546_, _14542_);
  or _66108_ (_14548_, _07299_, _07297_);
  and _66109_ (_14549_, _14548_, _07300_);
  or _66110_ (_14550_, _14549_, _06800_);
  and _66111_ (_14551_, _14550_, _03500_);
  and _66112_ (_14552_, _14551_, _14547_);
  nor _66113_ (_14553_, _12716_, _07315_);
  or _66114_ (_14554_, _14553_, _14513_);
  and _66115_ (_14555_, _14554_, _03499_);
  or _66116_ (_14556_, _14555_, _07314_);
  or _66117_ (_14557_, _14556_, _14552_);
  or _66118_ (_14558_, _14534_, _06039_);
  and _66119_ (_14559_, _14558_, _14557_);
  or _66120_ (_14560_, _14559_, _03479_);
  and _66121_ (_14561_, _06722_, _05221_);
  or _66122_ (_14562_, _14503_, _06044_);
  or _66123_ (_14563_, _14562_, _14561_);
  and _66124_ (_14564_, _14563_, _03474_);
  and _66125_ (_14565_, _14564_, _14560_);
  or _66126_ (_14566_, _14565_, _14512_);
  and _66127_ (_14567_, _14566_, _07677_);
  or _66128_ (_14568_, _14340_, _07615_);
  nor _66129_ (_14569_, _14452_, _07625_);
  or _66130_ (_14570_, _14569_, _07624_);
  nand _66131_ (_14571_, _14570_, _07662_);
  or _66132_ (_14572_, _14570_, _07662_);
  and _66133_ (_14573_, _14572_, _14571_);
  or _66134_ (_14574_, _14573_, _07675_);
  and _66135_ (_14575_, _14574_, _07328_);
  and _66136_ (_14576_, _14575_, _14568_);
  or _66137_ (_14577_, _14576_, _03437_);
  or _66138_ (_14578_, _14577_, _14567_);
  and _66139_ (_14579_, _14578_, _14509_);
  or _66140_ (_14580_, _14579_, _03636_);
  and _66141_ (_14581_, _12711_, _05221_);
  or _66142_ (_14582_, _14581_, _14503_);
  or _66143_ (_14583_, _14582_, _04499_);
  and _66144_ (_14584_, _14583_, _04501_);
  and _66145_ (_14585_, _14584_, _14580_);
  or _66146_ (_14586_, _14585_, _14506_);
  and _66147_ (_14587_, _14586_, _05769_);
  or _66148_ (_14588_, _14503_, _05761_);
  and _66149_ (_14589_, _14588_, _03754_);
  and _66150_ (_14590_, _14589_, _14508_);
  or _66151_ (_14591_, _14590_, _14587_);
  and _66152_ (_14592_, _14591_, _03753_);
  and _66153_ (_14593_, _14521_, _03752_);
  and _66154_ (_14594_, _14593_, _14588_);
  or _66155_ (_14595_, _14594_, _03758_);
  or _66156_ (_14596_, _14595_, _14592_);
  nor _66157_ (_14597_, _12710_, _06762_);
  or _66158_ (_14598_, _14503_, _03759_);
  or _66159_ (_14599_, _14598_, _14597_);
  and _66160_ (_14600_, _14599_, _04517_);
  and _66161_ (_14601_, _14600_, _14596_);
  nor _66162_ (_14602_, _12843_, _06762_);
  or _66163_ (_14603_, _14602_, _14503_);
  and _66164_ (_14604_, _14603_, _03760_);
  or _66165_ (_14605_, _14604_, _03790_);
  or _66166_ (_14606_, _14605_, _14601_);
  or _66167_ (_14607_, _14518_, _04192_);
  and _66168_ (_14608_, _14607_, _03152_);
  and _66169_ (_14609_, _14608_, _14606_);
  and _66170_ (_14610_, _14515_, _03151_);
  or _66171_ (_14611_, _14610_, _03520_);
  or _66172_ (_14612_, _14611_, _14609_);
  and _66173_ (_14613_, _12893_, _05221_);
  or _66174_ (_14614_, _14503_, _03521_);
  or _66175_ (_14615_, _14614_, _14613_);
  and _66176_ (_14616_, _14615_, _42963_);
  and _66177_ (_14617_, _14616_, _14612_);
  or _66178_ (_14618_, _14617_, _14502_);
  and _66179_ (_43199_, _14618_, _41755_);
  nor _66180_ (_14619_, _42963_, _07460_);
  nor _66181_ (_14620_, _05221_, _07460_);
  and _66182_ (_14621_, _13042_, _05221_);
  or _66183_ (_14622_, _14621_, _14620_);
  and _66184_ (_14623_, _14622_, _03769_);
  nor _66185_ (_14624_, _13021_, _06762_);
  or _66186_ (_14625_, _14624_, _14620_);
  and _66187_ (_14626_, _14625_, _03221_);
  nor _66188_ (_14627_, _05422_, _06762_);
  or _66189_ (_14628_, _14627_, _14620_);
  or _66190_ (_14629_, _14628_, _06039_);
  nor _66191_ (_14630_, _05785_, _07460_);
  and _66192_ (_14631_, _12914_, _05785_);
  or _66193_ (_14632_, _14631_, _14630_);
  and _66194_ (_14633_, _14632_, _03512_);
  nor _66195_ (_14634_, _12930_, _06762_);
  or _66196_ (_14635_, _14634_, _14620_);
  or _66197_ (_14636_, _14635_, _04444_);
  and _66198_ (_14637_, _05221_, \oc8051_golden_model_1.ACC [5]);
  or _66199_ (_14638_, _14637_, _14620_);
  and _66200_ (_14639_, _14638_, _04426_);
  nor _66201_ (_14640_, _04426_, _07460_);
  or _66202_ (_14641_, _14640_, _03570_);
  or _66203_ (_14642_, _14641_, _14639_);
  and _66204_ (_14643_, _14642_, _03517_);
  and _66205_ (_14644_, _14643_, _14636_);
  and _66206_ (_14645_, _12934_, _05785_);
  or _66207_ (_14646_, _14645_, _14630_);
  and _66208_ (_14647_, _14646_, _03516_);
  or _66209_ (_14648_, _14647_, _03568_);
  or _66210_ (_14649_, _14648_, _14644_);
  or _66211_ (_14650_, _14628_, _03983_);
  and _66212_ (_14651_, _14650_, _14649_);
  or _66213_ (_14652_, _14651_, _03575_);
  or _66214_ (_14653_, _14638_, _03583_);
  and _66215_ (_14654_, _14653_, _03513_);
  and _66216_ (_14655_, _14654_, _14652_);
  or _66217_ (_14656_, _14655_, _14633_);
  and _66218_ (_14657_, _14656_, _03506_);
  or _66219_ (_14658_, _14630_, _12949_);
  and _66220_ (_14659_, _14658_, _03505_);
  and _66221_ (_14660_, _14659_, _14646_);
  or _66222_ (_14661_, _14660_, _06794_);
  or _66223_ (_14662_, _14661_, _14657_);
  or _66224_ (_14663_, _07004_, _07003_);
  not _66225_ (_14664_, _14663_);
  nor _66226_ (_14665_, _14664_, _07301_);
  and _66227_ (_14666_, _14664_, _07301_);
  or _66228_ (_14667_, _14666_, _14665_);
  or _66229_ (_14668_, _14667_, _06800_);
  and _66230_ (_14669_, _14668_, _03500_);
  and _66231_ (_14670_, _14669_, _14662_);
  nor _66232_ (_14671_, _12912_, _07315_);
  or _66233_ (_14672_, _14671_, _14630_);
  and _66234_ (_14673_, _14672_, _03499_);
  or _66235_ (_14674_, _14673_, _07314_);
  or _66236_ (_14675_, _14674_, _14670_);
  and _66237_ (_14676_, _14675_, _14629_);
  or _66238_ (_14677_, _14676_, _03479_);
  and _66239_ (_14678_, _06721_, _05221_);
  or _66240_ (_14679_, _14620_, _06044_);
  or _66241_ (_14680_, _14679_, _14678_);
  and _66242_ (_14681_, _14680_, _03474_);
  and _66243_ (_14682_, _14681_, _14677_);
  or _66244_ (_14683_, _14682_, _14626_);
  and _66245_ (_14684_, _14683_, _07677_);
  and _66246_ (_14685_, _07607_, _07328_);
  and _66247_ (_14686_, _14685_, _07675_);
  not _66248_ (_14687_, _07653_);
  and _66249_ (_14688_, _14571_, _14687_);
  nor _66250_ (_14689_, _14688_, _07663_);
  and _66251_ (_14690_, _14688_, _07663_);
  or _66252_ (_14691_, _14690_, _14689_);
  nor _66253_ (_14692_, _07675_, _07677_);
  and _66254_ (_14693_, _14692_, _14691_);
  or _66255_ (_14694_, _14693_, _14686_);
  or _66256_ (_14695_, _14694_, _03437_);
  or _66257_ (_14696_, _14695_, _14684_);
  and _66258_ (_14697_, _06211_, _05221_);
  or _66259_ (_14698_, _14697_, _14620_);
  or _66260_ (_14699_, _14698_, _03438_);
  and _66261_ (_14700_, _14699_, _14696_);
  or _66262_ (_14701_, _14700_, _03636_);
  and _66263_ (_14702_, _13036_, _05221_);
  or _66264_ (_14703_, _14702_, _14620_);
  or _66265_ (_14704_, _14703_, _04499_);
  and _66266_ (_14705_, _14704_, _04501_);
  and _66267_ (_14706_, _14705_, _14701_);
  or _66268_ (_14707_, _14706_, _14623_);
  and _66269_ (_14708_, _14707_, _05769_);
  or _66270_ (_14709_, _14620_, _05472_);
  and _66271_ (_14710_, _14709_, _03754_);
  and _66272_ (_14711_, _14710_, _14698_);
  or _66273_ (_14712_, _14711_, _14708_);
  and _66274_ (_14713_, _14712_, _03753_);
  and _66275_ (_14714_, _14638_, _03752_);
  and _66276_ (_14715_, _14714_, _14709_);
  or _66277_ (_14716_, _14715_, _03758_);
  or _66278_ (_14717_, _14716_, _14713_);
  nor _66279_ (_14718_, _13035_, _06762_);
  or _66280_ (_14719_, _14620_, _03759_);
  or _66281_ (_14720_, _14719_, _14718_);
  and _66282_ (_14721_, _14720_, _04517_);
  and _66283_ (_14722_, _14721_, _14717_);
  nor _66284_ (_14723_, _13041_, _06762_);
  or _66285_ (_14724_, _14723_, _14620_);
  and _66286_ (_14725_, _14724_, _03760_);
  or _66287_ (_14726_, _14725_, _03790_);
  or _66288_ (_14727_, _14726_, _14722_);
  or _66289_ (_14728_, _14635_, _04192_);
  and _66290_ (_14729_, _14728_, _03152_);
  and _66291_ (_14730_, _14729_, _14727_);
  and _66292_ (_14731_, _14632_, _03151_);
  or _66293_ (_14732_, _14731_, _03520_);
  or _66294_ (_14733_, _14732_, _14730_);
  and _66295_ (_14734_, _13097_, _05221_);
  or _66296_ (_14735_, _14620_, _03521_);
  or _66297_ (_14736_, _14735_, _14734_);
  and _66298_ (_14737_, _14736_, _42963_);
  and _66299_ (_14738_, _14737_, _14733_);
  or _66300_ (_14739_, _14738_, _14619_);
  and _66301_ (_43200_, _14739_, _41755_);
  nor _66302_ (_14740_, _42963_, _07592_);
  nor _66303_ (_14741_, _05221_, _07592_);
  and _66304_ (_14742_, _13259_, _05221_);
  or _66305_ (_14743_, _14742_, _14741_);
  and _66306_ (_14744_, _14743_, _03769_);
  and _66307_ (_14745_, _13244_, _05221_);
  or _66308_ (_14746_, _14745_, _14741_);
  or _66309_ (_14747_, _14746_, _03438_);
  nor _66310_ (_14748_, _13237_, _06762_);
  or _66311_ (_14749_, _14748_, _14741_);
  and _66312_ (_14750_, _14749_, _03221_);
  nor _66313_ (_14751_, _05327_, _06762_);
  or _66314_ (_14752_, _14751_, _14741_);
  or _66315_ (_14753_, _14752_, _06039_);
  nor _66316_ (_14754_, _05785_, _07592_);
  and _66317_ (_14755_, _13130_, _05785_);
  or _66318_ (_14756_, _14755_, _14754_);
  and _66319_ (_14757_, _14756_, _03512_);
  nor _66320_ (_14758_, _13122_, _06762_);
  or _66321_ (_14759_, _14758_, _14741_);
  or _66322_ (_14760_, _14759_, _04444_);
  and _66323_ (_14761_, _05221_, \oc8051_golden_model_1.ACC [6]);
  or _66324_ (_14762_, _14761_, _14741_);
  and _66325_ (_14763_, _14762_, _04426_);
  nor _66326_ (_14764_, _04426_, _07592_);
  or _66327_ (_14765_, _14764_, _03570_);
  or _66328_ (_14766_, _14765_, _14763_);
  and _66329_ (_14767_, _14766_, _03517_);
  and _66330_ (_14768_, _14767_, _14760_);
  and _66331_ (_14769_, _13145_, _05785_);
  or _66332_ (_14770_, _14769_, _14754_);
  and _66333_ (_14771_, _14770_, _03516_);
  or _66334_ (_14772_, _14771_, _03568_);
  or _66335_ (_14773_, _14772_, _14768_);
  or _66336_ (_14774_, _14752_, _03983_);
  and _66337_ (_14775_, _14774_, _14773_);
  or _66338_ (_14776_, _14775_, _03575_);
  or _66339_ (_14777_, _14762_, _03583_);
  and _66340_ (_14778_, _14777_, _03513_);
  and _66341_ (_14779_, _14778_, _14776_);
  or _66342_ (_14780_, _14779_, _14757_);
  and _66343_ (_14781_, _14780_, _03506_);
  or _66344_ (_14782_, _14754_, _13160_);
  and _66345_ (_14783_, _14782_, _03505_);
  and _66346_ (_14784_, _14783_, _14770_);
  or _66347_ (_14785_, _14784_, _06794_);
  or _66348_ (_14786_, _14785_, _14781_);
  nor _66349_ (_14787_, _07307_, _07303_);
  nor _66350_ (_14788_, _14787_, _07308_);
  or _66351_ (_14789_, _14788_, _06800_);
  and _66352_ (_14790_, _14789_, _03500_);
  and _66353_ (_14791_, _14790_, _14786_);
  nor _66354_ (_14792_, _13178_, _07315_);
  or _66355_ (_14793_, _14792_, _14754_);
  and _66356_ (_14794_, _14793_, _03499_);
  or _66357_ (_14795_, _14794_, _07314_);
  or _66358_ (_14796_, _14795_, _14791_);
  and _66359_ (_14797_, _14796_, _14753_);
  or _66360_ (_14798_, _14797_, _03479_);
  and _66361_ (_14799_, _06713_, _05221_);
  or _66362_ (_14800_, _14741_, _06044_);
  or _66363_ (_14801_, _14800_, _14799_);
  and _66364_ (_14802_, _14801_, _03474_);
  and _66365_ (_14803_, _14802_, _14798_);
  or _66366_ (_14804_, _14803_, _14750_);
  and _66367_ (_14805_, _14804_, _07677_);
  or _66368_ (_14806_, _14340_, _07598_);
  nor _66369_ (_14807_, _14688_, _07608_);
  or _66370_ (_14808_, _14807_, _07609_);
  or _66371_ (_14809_, _14808_, _07665_);
  nand _66372_ (_14810_, _14808_, _07665_);
  and _66373_ (_14811_, _14810_, _14809_);
  or _66374_ (_14812_, _14811_, _07675_);
  and _66375_ (_14813_, _14812_, _07328_);
  and _66376_ (_14814_, _14813_, _14806_);
  or _66377_ (_14815_, _14814_, _03437_);
  or _66378_ (_14816_, _14815_, _14805_);
  and _66379_ (_14817_, _14816_, _14747_);
  or _66380_ (_14818_, _14817_, _03636_);
  and _66381_ (_14819_, _13253_, _05221_);
  or _66382_ (_14820_, _14819_, _14741_);
  or _66383_ (_14821_, _14820_, _04499_);
  and _66384_ (_14822_, _14821_, _04501_);
  and _66385_ (_14823_, _14822_, _14818_);
  or _66386_ (_14824_, _14823_, _14744_);
  and _66387_ (_14825_, _14824_, _05769_);
  or _66388_ (_14826_, _14741_, _05377_);
  and _66389_ (_14827_, _14826_, _03754_);
  and _66390_ (_14828_, _14827_, _14746_);
  or _66391_ (_14829_, _14828_, _14825_);
  and _66392_ (_14830_, _14829_, _03753_);
  and _66393_ (_14831_, _14762_, _03752_);
  and _66394_ (_14832_, _14831_, _14826_);
  or _66395_ (_14833_, _14832_, _03758_);
  or _66396_ (_14834_, _14833_, _14830_);
  nor _66397_ (_14835_, _13251_, _06762_);
  or _66398_ (_14836_, _14741_, _03759_);
  or _66399_ (_14837_, _14836_, _14835_);
  and _66400_ (_14838_, _14837_, _04517_);
  and _66401_ (_14839_, _14838_, _14834_);
  nor _66402_ (_14840_, _13258_, _06762_);
  or _66403_ (_14841_, _14840_, _14741_);
  and _66404_ (_14842_, _14841_, _03760_);
  or _66405_ (_14843_, _14842_, _03790_);
  or _66406_ (_14844_, _14843_, _14839_);
  or _66407_ (_14845_, _14759_, _04192_);
  and _66408_ (_14846_, _14845_, _03152_);
  and _66409_ (_14847_, _14846_, _14844_);
  and _66410_ (_14848_, _14756_, _03151_);
  or _66411_ (_14849_, _14848_, _03520_);
  or _66412_ (_14850_, _14849_, _14847_);
  and _66413_ (_14851_, _13312_, _05221_);
  or _66414_ (_14852_, _14741_, _03521_);
  or _66415_ (_14853_, _14852_, _14851_);
  and _66416_ (_14854_, _14853_, _42963_);
  and _66417_ (_14855_, _14854_, _14850_);
  or _66418_ (_14856_, _14855_, _14740_);
  and _66419_ (_43201_, _14856_, _41755_);
  nor _66420_ (_14857_, _42963_, _03321_);
  nand _66421_ (_14858_, _07729_, _05834_);
  nor _66422_ (_14859_, _08334_, _03321_);
  nor _66423_ (_14860_, _14859_, _08335_);
  nand _66424_ (_14861_, _08523_, _14860_);
  nor _66425_ (_14862_, _07890_, _03321_);
  nor _66426_ (_14863_, _14862_, _08016_);
  nand _66427_ (_14864_, _14863_, _04155_);
  nand _66428_ (_14865_, _08477_, _10394_);
  and _66429_ (_14866_, _04439_, _03321_);
  nand _66430_ (_14867_, _08456_, _14866_);
  or _66431_ (_14868_, _11994_, _07911_);
  and _66432_ (_14869_, _14868_, _07910_);
  nand _66433_ (_14870_, _03191_, _03147_);
  not _66434_ (_14871_, _14870_);
  and _66435_ (_14872_, _14871_, _07806_);
  nor _66436_ (_14873_, _05227_, _03321_);
  and _66437_ (_14874_, _11990_, _05227_);
  nor _66438_ (_14875_, _14874_, _14873_);
  nand _66439_ (_14876_, _14875_, _03636_);
  and _66440_ (_14877_, _06478_, _03321_);
  nor _66441_ (_14878_, _14877_, _07757_);
  or _66442_ (_14879_, _14878_, _04126_);
  nand _66443_ (_14880_, _03471_, _03231_);
  nor _66444_ (_14881_, _11975_, _07918_);
  nor _66445_ (_14882_, _14881_, _14873_);
  nor _66446_ (_14883_, _14882_, _03474_);
  and _66447_ (_14884_, _05227_, _04419_);
  nor _66448_ (_14885_, _14884_, _14873_);
  nand _66449_ (_14886_, _14885_, _07314_);
  nand _66450_ (_14887_, _14860_, _08108_);
  or _66451_ (_14888_, _07927_, _04419_);
  nor _66452_ (_14889_, _07935_, _04438_);
  or _66453_ (_14890_, _14889_, _06715_);
  and _66454_ (_14891_, _07933_, _04419_);
  or _66455_ (_14892_, _04012_, \oc8051_golden_model_1.ACC [0]);
  nand _66456_ (_14893_, _04012_, \oc8051_golden_model_1.ACC [0]);
  nand _66457_ (_14894_, _14893_, _14892_);
  nor _66458_ (_14895_, _14894_, _07933_);
  or _66459_ (_14896_, _14895_, _07935_);
  or _66460_ (_14897_, _14896_, _14891_);
  and _66461_ (_14898_, _14897_, _03208_);
  or _66462_ (_14899_, _14898_, _04438_);
  and _66463_ (_14900_, _14899_, _04444_);
  and _66464_ (_14901_, _14900_, _14890_);
  and _66465_ (_14902_, _05941_, _05227_);
  nor _66466_ (_14903_, _14902_, _14873_);
  nor _66467_ (_14904_, _14903_, _04444_);
  or _66468_ (_14905_, _14904_, _03516_);
  or _66469_ (_14906_, _14905_, _14901_);
  nor _66470_ (_14907_, _05792_, _03321_);
  and _66471_ (_14908_, _11887_, _05792_);
  nor _66472_ (_14909_, _14908_, _14907_);
  nand _66473_ (_14910_, _14909_, _03516_);
  and _66474_ (_14911_, _14910_, _03983_);
  and _66475_ (_14912_, _14911_, _14906_);
  nor _66476_ (_14913_, _14885_, _03983_);
  or _66477_ (_14914_, _14913_, _07928_);
  or _66478_ (_14915_, _14914_, _14912_);
  and _66479_ (_14916_, _14915_, _14888_);
  or _66480_ (_14917_, _14916_, _04458_);
  or _66481_ (_14918_, _06715_, _07987_);
  and _66482_ (_14919_, _14918_, _03583_);
  and _66483_ (_14920_, _14919_, _14917_);
  nor _66484_ (_14921_, _08191_, _03583_);
  or _66485_ (_14922_, _14921_, _07991_);
  or _66486_ (_14923_, _14922_, _14920_);
  nand _66487_ (_14924_, _07991_, _07405_);
  and _66488_ (_14925_, _14924_, _14923_);
  or _66489_ (_14926_, _14925_, _03512_);
  or _66490_ (_14927_, _14873_, _03513_);
  and _66491_ (_14928_, _14927_, _03506_);
  and _66492_ (_14929_, _14928_, _14926_);
  nor _66493_ (_14930_, _14903_, _03506_);
  or _66494_ (_14931_, _14930_, _06794_);
  or _66495_ (_14932_, _14931_, _14929_);
  nand _66496_ (_14933_, _14863_, _11705_);
  not _66497_ (_14934_, _07266_);
  and _66498_ (_14935_, _14934_, _06794_);
  nor _66499_ (_14936_, _14935_, _11700_);
  and _66500_ (_14937_, _14936_, _14933_);
  and _66501_ (_14938_, _14937_, _14932_);
  nor _66502_ (_14939_, _14863_, _07922_);
  or _66503_ (_14940_, _14939_, _08035_);
  or _66504_ (_14941_, _14940_, _14938_);
  nor _66505_ (_14942_, _08087_, _03321_);
  nor _66506_ (_14943_, _14942_, _08088_);
  nand _66507_ (_14944_, _14943_, _08035_);
  and _66508_ (_14945_, _14944_, _03619_);
  and _66509_ (_14946_, _14945_, _14941_);
  nor _66510_ (_14947_, _08268_, _03321_);
  nor _66511_ (_14948_, _14947_, _08269_);
  nand _66512_ (_14949_, _14948_, _08109_);
  and _66513_ (_14950_, _14949_, _10431_);
  or _66514_ (_14951_, _14950_, _14946_);
  and _66515_ (_14952_, _14951_, _14887_);
  or _66516_ (_14953_, _14952_, _03311_);
  nand _66517_ (_14954_, _03471_, _03311_);
  and _66518_ (_14955_, _14954_, _03500_);
  and _66519_ (_14956_, _14955_, _14953_);
  nor _66520_ (_14957_, _11916_, _08358_);
  nor _66521_ (_14958_, _14957_, _14907_);
  nor _66522_ (_14959_, _14958_, _03500_);
  or _66523_ (_14960_, _14959_, _07314_);
  or _66524_ (_14961_, _14960_, _14956_);
  and _66525_ (_14962_, _14961_, _14886_);
  or _66526_ (_14963_, _14962_, _03479_);
  and _66527_ (_14964_, _06715_, _05227_);
  nor _66528_ (_14965_, _14964_, _14873_);
  nand _66529_ (_14966_, _14965_, _03479_);
  and _66530_ (_14967_, _14966_, _03474_);
  and _66531_ (_14968_, _14967_, _14963_);
  or _66532_ (_14969_, _14968_, _14883_);
  and _66533_ (_14970_, _14969_, _07677_);
  or _66534_ (_14971_, _14692_, _03231_);
  or _66535_ (_14972_, _14971_, _14970_);
  and _66536_ (_14973_, _14972_, _14880_);
  or _66537_ (_14974_, _14973_, _03437_);
  and _66538_ (_14975_, _05227_, _06202_);
  nor _66539_ (_14976_, _14975_, _14873_);
  nand _66540_ (_14977_, _14976_, _03437_);
  and _66541_ (_14978_, _14977_, _08386_);
  and _66542_ (_14979_, _14978_, _14974_);
  nor _66543_ (_14980_, _08386_, _03471_);
  or _66544_ (_14981_, _14980_, _08392_);
  or _66545_ (_14982_, _14981_, _14979_);
  nor _66546_ (_14983_, _14866_, _07806_);
  and _66547_ (_14984_, _08396_, _14983_);
  or _66548_ (_14985_, _14984_, _08397_);
  and _66549_ (_14986_, _14985_, _14982_);
  and _66550_ (_14987_, _08401_, _14983_);
  or _66551_ (_14988_, _14987_, _04128_);
  or _66552_ (_14989_, _14988_, _14986_);
  and _66553_ (_14990_, _11572_, _03193_);
  not _66554_ (_14991_, _14990_);
  not _66555_ (_14992_, _04128_);
  or _66556_ (_14993_, _14983_, _14992_);
  and _66557_ (_14994_, _14993_, _14991_);
  and _66558_ (_14995_, _14994_, _14989_);
  or _66559_ (_14996_, _14878_, _03043_);
  and _66560_ (_14997_, _14996_, _08405_);
  or _66561_ (_14998_, _14997_, _14995_);
  and _66562_ (_14999_, _14998_, _14879_);
  or _66563_ (_15000_, _14999_, _03767_);
  or _66564_ (_15001_, _11995_, _03768_);
  and _66565_ (_15002_, _15001_, _08416_);
  and _66566_ (_15003_, _15002_, _15000_);
  and _66567_ (_15004_, _08415_, _10395_);
  or _66568_ (_15005_, _15004_, _03636_);
  or _66569_ (_15006_, _15005_, _15003_);
  and _66570_ (_15007_, _15006_, _14876_);
  or _66571_ (_15008_, _15007_, _03769_);
  or _66572_ (_15009_, _14873_, _04501_);
  and _66573_ (_15010_, _15009_, _14870_);
  and _66574_ (_15011_, _15010_, _15008_);
  or _66575_ (_15012_, _15011_, _14872_);
  and _66576_ (_15013_, _15012_, _08446_);
  and _66577_ (_15014_, _08445_, _07757_);
  or _66578_ (_15015_, _15014_, _03755_);
  or _66579_ (_15016_, _15015_, _15013_);
  and _66580_ (_15017_, _15016_, _14869_);
  and _66581_ (_15018_, _08666_, _07909_);
  or _66582_ (_15019_, _15018_, _15017_);
  and _66583_ (_15020_, _15019_, _05769_);
  nor _66584_ (_15021_, _14976_, _14902_);
  and _66585_ (_15022_, _15021_, _04504_);
  or _66586_ (_15023_, _15022_, _08456_);
  or _66587_ (_15024_, _15023_, _15020_);
  and _66588_ (_15025_, _15024_, _14867_);
  nor _66589_ (_15026_, _08465_, _08455_);
  not _66590_ (_15027_, _15026_);
  or _66591_ (_15028_, _15027_, _15025_);
  not _66592_ (_15029_, _04161_);
  nand _66593_ (_15030_, _15027_, _14866_);
  and _66594_ (_15031_, _15030_, _15029_);
  and _66595_ (_15032_, _15031_, _15028_);
  nor _66596_ (_15033_, _14866_, _15029_);
  or _66597_ (_15034_, _15033_, _08469_);
  or _66598_ (_15035_, _15034_, _15032_);
  nand _66599_ (_15036_, _08469_, _14877_);
  and _66600_ (_15037_, _15036_, _08473_);
  and _66601_ (_15038_, _15037_, _15035_);
  nand _66602_ (_15039_, _11870_, _08480_);
  and _66603_ (_15040_, _15039_, _08479_);
  or _66604_ (_15041_, _15040_, _15038_);
  and _66605_ (_15042_, _15041_, _14865_);
  or _66606_ (_15043_, _15042_, _03758_);
  nor _66607_ (_15044_, _13061_, _04156_);
  nor _66608_ (_15045_, _11988_, _07918_);
  nor _66609_ (_15046_, _15045_, _14873_);
  and _66610_ (_15047_, _15046_, _03758_);
  nor _66611_ (_15048_, _15047_, _15044_);
  and _66612_ (_15049_, _15048_, _15043_);
  not _66613_ (_15050_, _14863_);
  and _66614_ (_15051_, _15044_, _15050_);
  or _66615_ (_15052_, _15051_, _04155_);
  or _66616_ (_15053_, _15052_, _15049_);
  and _66617_ (_15054_, _15053_, _14864_);
  or _66618_ (_15055_, _15054_, _07825_);
  nand _66619_ (_15056_, _07825_, _14943_);
  and _66620_ (_15057_, _15056_, _03766_);
  and _66621_ (_15058_, _15057_, _15055_);
  nand _66622_ (_15059_, _08557_, _14948_);
  and _66623_ (_15060_, _15059_, _08525_);
  or _66624_ (_15061_, _15060_, _15058_);
  and _66625_ (_15062_, _15061_, _14861_);
  or _66626_ (_15063_, _15062_, _08555_);
  nand _66627_ (_15064_, _08555_, _07888_);
  and _66628_ (_15065_, _15064_, _07775_);
  and _66629_ (_15066_, _15065_, _07779_);
  and _66630_ (_15067_, _15066_, _15063_);
  and _66631_ (_15068_, _11572_, _03171_);
  not _66632_ (_15069_, _07780_);
  and _66633_ (_15070_, _14983_, _15069_);
  or _66634_ (_15071_, _15070_, _15068_);
  or _66635_ (_15072_, _15071_, _15067_);
  and _66636_ (_15073_, _04004_, _03171_);
  not _66637_ (_15074_, _15073_);
  not _66638_ (_15075_, _15068_);
  or _66639_ (_15076_, _15075_, _14878_);
  and _66640_ (_15077_, _15076_, _15074_);
  and _66641_ (_15078_, _15077_, _15072_);
  and _66642_ (_15079_, _14878_, _15073_);
  or _66643_ (_15080_, _15079_, _03524_);
  or _66644_ (_15081_, _15080_, _15078_);
  nand _66645_ (_15082_, _10375_, _03524_);
  and _66646_ (_15083_, _15082_, _08598_);
  and _66647_ (_15084_, _15083_, _15081_);
  and _66648_ (_15085_, _08597_, _10395_);
  or _66649_ (_15086_, _15085_, _07729_);
  or _66650_ (_15087_, _15086_, _15084_);
  and _66651_ (_15088_, _15087_, _14858_);
  or _66652_ (_15089_, _15088_, _03790_);
  nand _66653_ (_15090_, _14903_, _03790_);
  and _66654_ (_15091_, _15090_, _08688_);
  and _66655_ (_15092_, _15091_, _15089_);
  nor _66656_ (_15093_, _08692_, _03321_);
  nor _66657_ (_15094_, _15093_, _10828_);
  or _66658_ (_15095_, _15094_, _15092_);
  nand _66659_ (_15096_, _08692_, _03233_);
  and _66660_ (_15097_, _15096_, _03152_);
  and _66661_ (_15098_, _15097_, _15095_);
  and _66662_ (_15099_, _14873_, _03151_);
  or _66663_ (_15100_, _15099_, _03520_);
  or _66664_ (_15101_, _15100_, _15098_);
  nand _66665_ (_15102_, _14903_, _03520_);
  and _66666_ (_15103_, _15102_, _08710_);
  and _66667_ (_15104_, _15103_, _15101_);
  nor _66668_ (_15105_, _08716_, _03321_);
  nor _66669_ (_15106_, _15105_, _10851_);
  or _66670_ (_15107_, _15106_, _15104_);
  nand _66671_ (_15108_, _08716_, _03233_);
  and _66672_ (_15109_, _15108_, _42963_);
  and _66673_ (_15110_, _15109_, _15107_);
  or _66674_ (_15111_, _15110_, _14857_);
  and _66675_ (_43203_, _15111_, _41755_);
  nor _66676_ (_15112_, _42963_, _03233_);
  nand _66677_ (_15113_, _07729_, _03321_);
  and _66678_ (_15114_, _08627_, _08625_);
  nor _66679_ (_15115_, _15114_, _08628_);
  or _66680_ (_15116_, _15115_, _03526_);
  and _66681_ (_15117_, _15116_, _08598_);
  and _66682_ (_15118_, _08536_, _08534_);
  nor _66683_ (_15119_, _15118_, _08537_);
  and _66684_ (_15120_, _15119_, _03765_);
  nand _66685_ (_15121_, _08477_, _08664_);
  nand _66686_ (_15122_, _08458_, _07804_);
  or _66687_ (_15123_, _12195_, _07911_);
  and _66688_ (_15124_, _15123_, _07910_);
  and _66689_ (_15125_, _14871_, _07803_);
  nor _66690_ (_15126_, _05227_, _03233_);
  and _66691_ (_15127_, _12191_, _05227_);
  nor _66692_ (_15128_, _15127_, _15126_);
  nand _66693_ (_15129_, _15128_, _03636_);
  nand _66694_ (_15130_, _04284_, _03231_);
  nor _66695_ (_15131_, _07918_, _04603_);
  nor _66696_ (_15132_, _15131_, _15126_);
  nand _66697_ (_15133_, _15132_, _07314_);
  and _66698_ (_15134_, \oc8051_golden_model_1.PSW [7], _03321_);
  and _66699_ (_15135_, _07888_, \oc8051_golden_model_1.ACC [0]);
  not _66700_ (_15136_, _15135_);
  and _66701_ (_15137_, _15136_, _06715_);
  nor _66702_ (_15138_, _15137_, _15134_);
  and _66703_ (_15139_, _15138_, _07756_);
  nor _66704_ (_15140_, _15138_, _07756_);
  or _66705_ (_15141_, _15140_, _15139_);
  or _66706_ (_15142_, _15141_, _08037_);
  nand _66707_ (_15143_, _07928_, _04603_);
  nand _66708_ (_15144_, _07933_, _04603_);
  nor _66709_ (_15145_, _04012_, _03233_);
  and _66710_ (_15146_, _04012_, _03233_);
  or _66711_ (_15147_, _15146_, _15145_);
  or _66712_ (_15148_, _15147_, _07933_);
  and _66713_ (_15149_, _15148_, _07936_);
  and _66714_ (_15150_, _15149_, _15144_);
  and _66715_ (_15151_, _15150_, _05847_);
  or _66716_ (_15152_, _15151_, _06714_);
  or _66717_ (_15153_, _15150_, _07935_);
  and _66718_ (_15154_, _15153_, _03208_);
  or _66719_ (_15155_, _15154_, _04438_);
  and _66720_ (_15156_, _15155_, _04444_);
  and _66721_ (_15157_, _15156_, _15152_);
  nor _66722_ (_15158_, _05227_, \oc8051_golden_model_1.ACC [1]);
  and _66723_ (_15159_, _12252_, _05227_);
  nor _66724_ (_15160_, _15159_, _15158_);
  and _66725_ (_15161_, _15160_, _03570_);
  or _66726_ (_15162_, _15161_, _07948_);
  or _66727_ (_15163_, _15162_, _15157_);
  nor _66728_ (_15164_, _07955_, \oc8051_golden_model_1.PSW [6]);
  nor _66729_ (_15165_, _15164_, \oc8051_golden_model_1.ACC [1]);
  and _66730_ (_15166_, _15164_, \oc8051_golden_model_1.ACC [1]);
  nor _66731_ (_15167_, _15166_, _15165_);
  nand _66732_ (_15168_, _15167_, _07948_);
  and _66733_ (_15169_, _15168_, _03576_);
  and _66734_ (_15170_, _15169_, _15163_);
  nor _66735_ (_15171_, _05792_, _03233_);
  and _66736_ (_15172_, _12083_, _05792_);
  nor _66737_ (_15173_, _15172_, _15171_);
  nor _66738_ (_15174_, _15173_, _03517_);
  nor _66739_ (_15175_, _15132_, _03983_);
  or _66740_ (_15176_, _15175_, _07928_);
  or _66741_ (_15177_, _15176_, _15174_);
  or _66742_ (_15178_, _15177_, _15170_);
  and _66743_ (_15179_, _15178_, _15143_);
  or _66744_ (_15180_, _15179_, _04458_);
  or _66745_ (_15181_, _06714_, _07987_);
  and _66746_ (_15182_, _15181_, _03583_);
  and _66747_ (_15183_, _15182_, _15180_);
  nor _66748_ (_15184_, _08177_, _03583_);
  or _66749_ (_15185_, _15184_, _07991_);
  or _66750_ (_15186_, _15185_, _15183_);
  nand _66751_ (_15187_, _07991_, _07399_);
  and _66752_ (_15188_, _15187_, _15186_);
  or _66753_ (_15189_, _15188_, _03512_);
  and _66754_ (_15190_, _12069_, _05792_);
  nor _66755_ (_15191_, _15190_, _15171_);
  nand _66756_ (_15192_, _15191_, _03512_);
  and _66757_ (_15193_, _15192_, _03506_);
  and _66758_ (_15194_, _15193_, _15189_);
  and _66759_ (_15195_, _15172_, _12098_);
  nor _66760_ (_15196_, _15195_, _15171_);
  nor _66761_ (_15197_, _15196_, _03506_);
  or _66762_ (_15198_, _15197_, _06794_);
  or _66763_ (_15199_, _15198_, _15194_);
  and _66764_ (_15200_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor _66765_ (_15201_, _15200_, _07637_);
  nor _66766_ (_15202_, _15201_, _07267_);
  or _66767_ (_15203_, _15202_, _06800_);
  and _66768_ (_15204_, _15203_, _07922_);
  and _66769_ (_15205_, _15204_, _15199_);
  and _66770_ (_15206_, _15136_, _04419_);
  nor _66771_ (_15207_, _15206_, _15134_);
  and _66772_ (_15208_, _15207_, _07805_);
  nor _66773_ (_15209_, _15207_, _07805_);
  or _66774_ (_15210_, _15209_, _15208_);
  and _66775_ (_15211_, _15210_, _07923_);
  or _66776_ (_15212_, _15211_, _08035_);
  or _66777_ (_15213_, _15212_, _15205_);
  and _66778_ (_15214_, _15213_, _15142_);
  or _66779_ (_15215_, _15214_, _03614_);
  nor _66780_ (_15216_, _08191_, _15135_);
  nor _66781_ (_15217_, _15216_, _15134_);
  and _66782_ (_15218_, _15217_, _08625_);
  nor _66783_ (_15219_, _15217_, _08625_);
  or _66784_ (_15220_, _15219_, _15218_);
  nand _66785_ (_15221_, _15220_, _03614_);
  and _66786_ (_15222_, _15221_, _08109_);
  and _66787_ (_15223_, _15222_, _15215_);
  nor _66788_ (_15224_, _15135_, _03471_);
  nor _66789_ (_15225_, _15224_, _15134_);
  and _66790_ (_15226_, _15225_, _08665_);
  nor _66791_ (_15227_, _15225_, _08665_);
  nor _66792_ (_15228_, _15227_, _15226_);
  nor _66793_ (_15229_, _15228_, _08109_);
  or _66794_ (_15230_, _15229_, _03311_);
  or _66795_ (_15231_, _15230_, _15223_);
  nand _66796_ (_15232_, _04284_, _03311_);
  and _66797_ (_15233_, _15232_, _03500_);
  and _66798_ (_15234_, _15233_, _15231_);
  nor _66799_ (_15235_, _12116_, _08358_);
  nor _66800_ (_15236_, _15235_, _15171_);
  nor _66801_ (_15237_, _15236_, _03500_);
  or _66802_ (_15238_, _15237_, _07314_);
  or _66803_ (_15239_, _15238_, _15234_);
  and _66804_ (_15240_, _15239_, _15133_);
  or _66805_ (_15241_, _15240_, _03479_);
  and _66806_ (_15242_, _06714_, _05227_);
  nor _66807_ (_15243_, _15242_, _15126_);
  nand _66808_ (_15244_, _15243_, _03479_);
  and _66809_ (_15245_, _15244_, _03474_);
  and _66810_ (_15246_, _15245_, _15241_);
  nor _66811_ (_15247_, _12176_, _07918_);
  nor _66812_ (_15248_, _15247_, _15126_);
  nor _66813_ (_15249_, _15248_, _03474_);
  or _66814_ (_15250_, _15249_, _07328_);
  or _66815_ (_15251_, _15250_, _15246_);
  nand _66816_ (_15252_, _07585_, _07328_);
  and _66817_ (_15253_, _15252_, _15251_);
  or _66818_ (_15254_, _15253_, _03231_);
  and _66819_ (_15255_, _15254_, _15130_);
  or _66820_ (_15256_, _15255_, _03437_);
  and _66821_ (_15257_, _05227_, _04317_);
  nor _66822_ (_15258_, _15257_, _15158_);
  or _66823_ (_15259_, _15258_, _03438_);
  and _66824_ (_15260_, _15259_, _08386_);
  and _66825_ (_15261_, _15260_, _15256_);
  nor _66826_ (_15262_, _08386_, _04284_);
  or _66827_ (_15263_, _15262_, _08392_);
  or _66828_ (_15264_, _15263_, _15261_);
  or _66829_ (_15265_, _07805_, _03936_);
  and _66830_ (_15266_, _15265_, _08396_);
  and _66831_ (_15267_, _15266_, _15264_);
  and _66832_ (_15268_, _03664_, _03193_);
  not _66833_ (_15269_, _15268_);
  and _66834_ (_15270_, _08396_, _15269_);
  nor _66835_ (_15271_, _07805_, _15268_);
  nor _66836_ (_15272_, _15271_, _15270_);
  or _66837_ (_15273_, _15272_, _04129_);
  or _66838_ (_15274_, _15273_, _15267_);
  or _66839_ (_15275_, _07805_, _14992_);
  and _66840_ (_15276_, _15275_, _08406_);
  and _66841_ (_15277_, _15276_, _15274_);
  and _66842_ (_15278_, _08405_, _07756_);
  or _66843_ (_15279_, _15278_, _03767_);
  or _66844_ (_15280_, _15279_, _15277_);
  or _66845_ (_15281_, _12197_, _03768_);
  and _66846_ (_15282_, _15281_, _08416_);
  and _66847_ (_15283_, _15282_, _15280_);
  and _66848_ (_15284_, _08415_, _08665_);
  or _66849_ (_15285_, _15284_, _03636_);
  or _66850_ (_15286_, _15285_, _15283_);
  and _66851_ (_15287_, _15286_, _15129_);
  or _66852_ (_15288_, _15287_, _03769_);
  or _66853_ (_15289_, _15126_, _04501_);
  and _66854_ (_15290_, _15289_, _14870_);
  and _66855_ (_15291_, _15290_, _15288_);
  or _66856_ (_15292_, _15291_, _15125_);
  and _66857_ (_15293_, _15292_, _08446_);
  and _66858_ (_15294_, _08445_, _07754_);
  or _66859_ (_15295_, _15294_, _03755_);
  or _66860_ (_15296_, _15295_, _15293_);
  and _66861_ (_15297_, _15296_, _15124_);
  and _66862_ (_15298_, _08663_, _07909_);
  or _66863_ (_15299_, _15298_, _15297_);
  and _66864_ (_15300_, _15299_, _05769_);
  and _66865_ (_15301_, _12190_, _05227_);
  nor _66866_ (_15302_, _15301_, _15126_);
  nor _66867_ (_15303_, _15302_, _04505_);
  or _66868_ (_15304_, _15303_, _08458_);
  or _66869_ (_15305_, _15304_, _15300_);
  and _66870_ (_15306_, _15305_, _15122_);
  or _66871_ (_15307_, _15306_, _08465_);
  nand _66872_ (_15308_, _08465_, _07804_);
  and _66873_ (_15309_, _15308_, _15029_);
  and _66874_ (_15310_, _15309_, _15307_);
  nor _66875_ (_15311_, _07804_, _15029_);
  or _66876_ (_15312_, _15311_, _08469_);
  or _66877_ (_15313_, _15312_, _15310_);
  nand _66878_ (_15314_, _08469_, _07755_);
  and _66879_ (_15315_, _15314_, _08473_);
  and _66880_ (_15316_, _15315_, _15313_);
  nand _66881_ (_15317_, _12196_, _08480_);
  and _66882_ (_15318_, _15317_, _08479_);
  or _66883_ (_15319_, _15318_, _15316_);
  and _66884_ (_15320_, _15319_, _15121_);
  or _66885_ (_15321_, _15320_, _03758_);
  nor _66886_ (_15322_, _12189_, _07918_);
  or _66887_ (_15323_, _15322_, _15126_);
  or _66888_ (_15324_, _15323_, _03759_);
  and _66889_ (_15325_, _15324_, _07830_);
  and _66890_ (_15326_, _15325_, _15321_);
  and _66891_ (_15327_, _07892_, _07887_);
  nor _66892_ (_15328_, _15327_, _07893_);
  and _66893_ (_15329_, _15328_, _08490_);
  or _66894_ (_15330_, _15329_, _07825_);
  or _66895_ (_15331_, _15330_, _15326_);
  and _66896_ (_15332_, _08504_, _08502_);
  nor _66897_ (_15333_, _15332_, _08505_);
  or _66898_ (_15334_, _15333_, _08495_);
  and _66899_ (_15335_, _15334_, _03766_);
  and _66900_ (_15336_, _15335_, _15331_);
  or _66901_ (_15337_, _15336_, _15120_);
  and _66902_ (_15338_, _15337_, _08557_);
  and _66903_ (_15339_, _08566_, _08564_);
  nor _66904_ (_15340_, _15339_, _08567_);
  and _66905_ (_15341_, _15340_, _08523_);
  or _66906_ (_15342_, _15341_, _08555_);
  or _66907_ (_15343_, _15342_, _15338_);
  nand _66908_ (_15344_, _08555_, _03321_);
  and _66909_ (_15345_, _15344_, _07780_);
  and _66910_ (_15346_, _15345_, _15343_);
  nor _66911_ (_15347_, _07806_, _07805_);
  nor _66912_ (_15348_, _15347_, _07807_);
  and _66913_ (_15349_, _15348_, _15069_);
  or _66914_ (_15350_, _15349_, _07731_);
  or _66915_ (_15351_, _15350_, _15346_);
  nor _66916_ (_15352_, _07757_, _07756_);
  nor _66917_ (_15353_, _15352_, _07758_);
  or _66918_ (_15354_, _15353_, _07732_);
  and _66919_ (_15355_, _15354_, _15351_);
  or _66920_ (_15356_, _15355_, _03524_);
  and _66921_ (_15357_, _15356_, _15117_);
  nor _66922_ (_15358_, _08666_, _08665_);
  nor _66923_ (_15359_, _15358_, _08667_);
  and _66924_ (_15360_, _15359_, _08597_);
  or _66925_ (_15361_, _15360_, _07729_);
  or _66926_ (_15362_, _15361_, _15357_);
  and _66927_ (_15363_, _15362_, _15113_);
  or _66928_ (_15364_, _15363_, _03790_);
  or _66929_ (_15365_, _15160_, _04192_);
  and _66930_ (_15366_, _15365_, _08688_);
  and _66931_ (_15367_, _15366_, _15364_);
  nor _66932_ (_15368_, _08717_, _08693_);
  and _66933_ (_15369_, _15368_, _11839_);
  nor _66934_ (_15370_, _15369_, _10828_);
  or _66935_ (_15371_, _15370_, _15367_);
  nand _66936_ (_15372_, _08692_, _07506_);
  and _66937_ (_15373_, _15372_, _03152_);
  and _66938_ (_15374_, _15373_, _15371_);
  nor _66939_ (_15375_, _15191_, _03152_);
  or _66940_ (_15376_, _15375_, _03520_);
  or _66941_ (_15377_, _15376_, _15374_);
  nor _66942_ (_15378_, _15159_, _15126_);
  nand _66943_ (_15379_, _15378_, _03520_);
  and _66944_ (_15380_, _15379_, _08710_);
  and _66945_ (_15381_, _15380_, _15377_);
  and _66946_ (_15382_, _15368_, _08709_);
  or _66947_ (_15383_, _15382_, _08716_);
  or _66948_ (_15384_, _15383_, _15381_);
  nand _66949_ (_15385_, _08716_, _07506_);
  and _66950_ (_15386_, _15385_, _42963_);
  and _66951_ (_15387_, _15386_, _15384_);
  or _66952_ (_15388_, _15387_, _15112_);
  and _66953_ (_43204_, _15388_, _41755_);
  nor _66954_ (_15389_, _42963_, _07506_);
  nand _66955_ (_15390_, _07729_, _03233_);
  and _66956_ (_15391_, _08629_, _08621_);
  nor _66957_ (_15392_, _15391_, _08630_);
  or _66958_ (_15393_, _15392_, _03526_);
  and _66959_ (_15394_, _15393_, _08598_);
  and _66960_ (_15395_, _08506_, _08079_);
  nor _66961_ (_15396_, _15395_, _08507_);
  or _66962_ (_15397_, _15396_, _08495_);
  nand _66963_ (_15398_, _08477_, _08660_);
  and _66964_ (_15399_, _14871_, _07799_);
  nor _66965_ (_15400_, _05227_, _07506_);
  and _66966_ (_15401_, _12273_, _05227_);
  nor _66967_ (_15402_, _15401_, _15400_);
  nand _66968_ (_15403_, _15402_, _03636_);
  or _66969_ (_15404_, _07752_, _04126_);
  nand _66970_ (_15405_, _03877_, _03231_);
  nor _66971_ (_15406_, _07918_, _05026_);
  nor _66972_ (_15407_, _15406_, _15400_);
  nand _66973_ (_15408_, _15407_, _07314_);
  nand _66974_ (_15409_, _07928_, _05026_);
  or _66975_ (_15410_, _14889_, _06718_);
  nor _66976_ (_15411_, _10288_, _05026_);
  and _66977_ (_15412_, _04012_, _07506_);
  nor _66978_ (_15413_, _04012_, _07506_);
  nor _66979_ (_15414_, _15413_, _15412_);
  nor _66980_ (_15415_, _15414_, _07933_);
  or _66981_ (_15416_, _15415_, _07935_);
  or _66982_ (_15417_, _15416_, _15411_);
  and _66983_ (_15418_, _15417_, _03208_);
  or _66984_ (_15419_, _15418_, _04438_);
  and _66985_ (_15420_, _15419_, _04444_);
  and _66986_ (_15421_, _15420_, _15410_);
  not _66987_ (_15422_, _15400_);
  or _66988_ (_15423_, _12282_, _07918_);
  and _66989_ (_15424_, _15423_, _15422_);
  nor _66990_ (_15425_, _15424_, _04444_);
  or _66991_ (_15426_, _15425_, _07948_);
  or _66992_ (_15427_, _15426_, _15421_);
  nand _66993_ (_15428_, _15164_, \oc8051_golden_model_1.ACC [2]);
  and _66994_ (_15429_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor _66995_ (_15430_, _15429_, _07954_);
  or _66996_ (_15431_, _15430_, _15164_);
  and _66997_ (_15432_, _15431_, _15428_);
  nand _66998_ (_15433_, _15432_, _07948_);
  and _66999_ (_15434_, _15433_, _03576_);
  and _67000_ (_15435_, _15434_, _15427_);
  nor _67001_ (_15436_, _05792_, _07506_);
  and _67002_ (_15437_, _12278_, _05792_);
  nor _67003_ (_15438_, _15437_, _15436_);
  nor _67004_ (_15439_, _15438_, _03517_);
  nor _67005_ (_15440_, _15407_, _03983_);
  or _67006_ (_15441_, _15440_, _07928_);
  or _67007_ (_15442_, _15441_, _15439_);
  or _67008_ (_15443_, _15442_, _15435_);
  and _67009_ (_15444_, _15443_, _15409_);
  or _67010_ (_15445_, _15444_, _04458_);
  or _67011_ (_15446_, _06718_, _07987_);
  and _67012_ (_15447_, _15446_, _03583_);
  and _67013_ (_15448_, _15447_, _15445_);
  nor _67014_ (_15449_, _08163_, _03583_);
  or _67015_ (_15450_, _15449_, _07991_);
  or _67016_ (_15451_, _15450_, _15448_);
  nand _67017_ (_15452_, _07991_, _07346_);
  and _67018_ (_15453_, _15452_, _15451_);
  or _67019_ (_15454_, _15453_, _03512_);
  and _67020_ (_15455_, _12276_, _05792_);
  nor _67021_ (_15456_, _15455_, _15436_);
  nand _67022_ (_15457_, _15456_, _03512_);
  and _67023_ (_15458_, _15457_, _03506_);
  and _67024_ (_15459_, _15458_, _15454_);
  and _67025_ (_15460_, _15437_, _12309_);
  nor _67026_ (_15461_, _15460_, _15436_);
  nor _67027_ (_15462_, _15461_, _03506_);
  or _67028_ (_15463_, _15462_, _06794_);
  or _67029_ (_15464_, _15463_, _15459_);
  nor _67030_ (_15465_, _07269_, _07267_);
  nor _67031_ (_15466_, _15465_, _07270_);
  or _67032_ (_15467_, _15466_, _06800_);
  and _67033_ (_15468_, _15467_, _15464_);
  or _67034_ (_15469_, _15468_, _07923_);
  and _67035_ (_15470_, _04603_, \oc8051_golden_model_1.ACC [1]);
  and _67036_ (_15471_, _04419_, _03321_);
  nor _67037_ (_15472_, _15471_, _07805_);
  nor _67038_ (_15473_, _15472_, _15470_);
  nor _67039_ (_15474_, _15473_, _07801_);
  and _67040_ (_15475_, _15473_, _07801_);
  nor _67041_ (_15476_, _15475_, _15474_);
  nor _67042_ (_15477_, _14983_, _07805_);
  not _67043_ (_15478_, _15477_);
  or _67044_ (_15479_, _15478_, _15476_);
  and _67045_ (_15480_, _15479_, \oc8051_golden_model_1.PSW [7]);
  nor _67046_ (_15481_, _15476_, \oc8051_golden_model_1.PSW [7]);
  or _67047_ (_15482_, _15481_, _15480_);
  nand _67048_ (_15483_, _15478_, _15476_);
  and _67049_ (_15484_, _15483_, _15482_);
  nand _67050_ (_15485_, _15484_, _07923_);
  and _67051_ (_15486_, _15485_, _15469_);
  or _67052_ (_15487_, _15486_, _08035_);
  and _67053_ (_15488_, _06433_, \oc8051_golden_model_1.ACC [1]);
  and _67054_ (_15489_, _06715_, _03321_);
  nor _67055_ (_15490_, _15489_, _07756_);
  nor _67056_ (_15491_, _15490_, _15488_);
  nor _67057_ (_15492_, _15491_, _07752_);
  and _67058_ (_15493_, _15491_, _07752_);
  nor _67059_ (_15494_, _15493_, _15492_);
  nor _67060_ (_15495_, _14878_, _07756_);
  not _67061_ (_15497_, _15495_);
  or _67062_ (_15498_, _15497_, _15494_);
  and _67063_ (_15499_, _15498_, \oc8051_golden_model_1.PSW [7]);
  nor _67064_ (_15500_, _15494_, \oc8051_golden_model_1.PSW [7]);
  or _67065_ (_15501_, _15500_, _15499_);
  nand _67066_ (_15502_, _15497_, _15494_);
  and _67067_ (_15503_, _15502_, _15501_);
  nand _67068_ (_15504_, _15503_, _08035_);
  and _67069_ (_15505_, _15504_, _15487_);
  or _67070_ (_15506_, _15505_, _03614_);
  nor _67071_ (_15508_, _10373_, _08623_);
  or _67072_ (_15509_, _15508_, _08624_);
  and _67073_ (_15510_, _08621_, _15509_);
  nor _67074_ (_15511_, _08621_, _15509_);
  nor _67075_ (_15512_, _15511_, _15510_);
  and _67076_ (_15513_, _10376_, \oc8051_golden_model_1.PSW [7]);
  not _67077_ (_15514_, _15513_);
  nor _67078_ (_15515_, _15514_, _15512_);
  and _67079_ (_15516_, _15514_, _15512_);
  nor _67080_ (_15517_, _15516_, _15515_);
  nand _67081_ (_15519_, _15517_, _03614_);
  and _67082_ (_15520_, _15519_, _08109_);
  and _67083_ (_15521_, _15520_, _15506_);
  nor _67084_ (_15522_, _03471_, \oc8051_golden_model_1.ACC [0]);
  nor _67085_ (_15523_, _15522_, _08665_);
  nor _67086_ (_15524_, _15523_, _11491_);
  nor _67087_ (_15525_, _08661_, _15524_);
  and _67088_ (_15526_, _08661_, _15524_);
  nor _67089_ (_15527_, _15526_, _15525_);
  not _67090_ (_15528_, _10396_);
  or _67091_ (_15530_, _15528_, _15527_);
  and _67092_ (_15531_, _15530_, \oc8051_golden_model_1.PSW [7]);
  nor _67093_ (_15532_, _15527_, \oc8051_golden_model_1.PSW [7]);
  or _67094_ (_15533_, _15532_, _15531_);
  nand _67095_ (_15534_, _15528_, _15527_);
  and _67096_ (_15535_, _15534_, _15533_);
  nor _67097_ (_15536_, _15535_, _08109_);
  or _67098_ (_15537_, _15536_, _03311_);
  or _67099_ (_15538_, _15537_, _15521_);
  nand _67100_ (_15539_, _03877_, _03311_);
  and _67101_ (_15541_, _15539_, _03500_);
  and _67102_ (_15542_, _15541_, _15538_);
  nor _67103_ (_15543_, _12326_, _08358_);
  nor _67104_ (_15544_, _15543_, _15436_);
  nor _67105_ (_15545_, _15544_, _03500_);
  or _67106_ (_15546_, _15545_, _07314_);
  or _67107_ (_15547_, _15546_, _15542_);
  and _67108_ (_15548_, _15547_, _15408_);
  or _67109_ (_15549_, _15548_, _03479_);
  and _67110_ (_15550_, _06718_, _05227_);
  nor _67111_ (_15552_, _15550_, _15400_);
  nand _67112_ (_15553_, _15552_, _03479_);
  and _67113_ (_15554_, _15553_, _03474_);
  and _67114_ (_15555_, _15554_, _15549_);
  nor _67115_ (_15556_, _12384_, _07918_);
  nor _67116_ (_15557_, _15556_, _15400_);
  nor _67117_ (_15558_, _15557_, _03474_);
  or _67118_ (_15559_, _15558_, _07328_);
  or _67119_ (_15560_, _15559_, _15555_);
  or _67120_ (_15561_, _07520_, _07677_);
  and _67121_ (_15563_, _15561_, _15560_);
  or _67122_ (_15564_, _15563_, _03231_);
  and _67123_ (_15565_, _15564_, _15405_);
  or _67124_ (_15566_, _15565_, _03437_);
  and _67125_ (_15567_, _05227_, _06261_);
  nor _67126_ (_15568_, _15567_, _15400_);
  nand _67127_ (_15569_, _15568_, _03437_);
  and _67128_ (_15570_, _15569_, _08386_);
  and _67129_ (_15571_, _15570_, _15566_);
  nor _67130_ (_15572_, _08386_, _03877_);
  or _67131_ (_15574_, _15572_, _08392_);
  or _67132_ (_15575_, _15574_, _15571_);
  or _67133_ (_15576_, _07801_, _03936_);
  and _67134_ (_15577_, _15576_, _08396_);
  and _67135_ (_15578_, _15577_, _15575_);
  and _67136_ (_15579_, _08401_, _07801_);
  or _67137_ (_15580_, _15579_, _15578_);
  and _67138_ (_15581_, _15580_, _15269_);
  not _67139_ (_15582_, _04129_);
  nand _67140_ (_15583_, _07801_, _15268_);
  nand _67141_ (_15585_, _15583_, _15582_);
  or _67142_ (_15586_, _15585_, _15581_);
  and _67143_ (_15587_, _03650_, _03193_);
  not _67144_ (_15588_, _15587_);
  or _67145_ (_15589_, _07801_, _15588_);
  and _67146_ (_15590_, _15589_, _14991_);
  and _67147_ (_15591_, _15590_, _15586_);
  or _67148_ (_15592_, _07752_, _03043_);
  and _67149_ (_15593_, _15592_, _08405_);
  or _67150_ (_15594_, _15593_, _15591_);
  and _67151_ (_15596_, _15594_, _15404_);
  or _67152_ (_15597_, _15596_, _03767_);
  or _67153_ (_15598_, _12401_, _03768_);
  and _67154_ (_15599_, _15598_, _08416_);
  and _67155_ (_15600_, _15599_, _15597_);
  and _67156_ (_15601_, _08415_, _08661_);
  or _67157_ (_15602_, _15601_, _03636_);
  or _67158_ (_15603_, _15602_, _15600_);
  and _67159_ (_15604_, _15603_, _15403_);
  or _67160_ (_15605_, _15604_, _03769_);
  or _67161_ (_15607_, _15400_, _04501_);
  and _67162_ (_15608_, _15607_, _14870_);
  and _67163_ (_15609_, _15608_, _15605_);
  or _67164_ (_15610_, _15609_, _15399_);
  and _67165_ (_15611_, _15610_, _08446_);
  and _67166_ (_15612_, _08445_, _07750_);
  or _67167_ (_15613_, _15612_, _03755_);
  or _67168_ (_15614_, _15613_, _15611_);
  or _67169_ (_15615_, _12399_, _07911_);
  and _67170_ (_15616_, _15615_, _07910_);
  and _67171_ (_15618_, _15616_, _15614_);
  and _67172_ (_15619_, _08659_, _07909_);
  or _67173_ (_15620_, _15619_, _15618_);
  and _67174_ (_15621_, _15620_, _05769_);
  not _67175_ (_15622_, _09953_);
  or _67176_ (_15623_, _15568_, _12400_);
  nor _67177_ (_15624_, _15623_, _04505_);
  or _67178_ (_15625_, _15624_, _15622_);
  or _67179_ (_15626_, _15625_, _15621_);
  not _67180_ (_15627_, _09954_);
  nand _67181_ (_15629_, _15622_, _07800_);
  and _67182_ (_15630_, _15629_, _15627_);
  and _67183_ (_15631_, _15630_, _15626_);
  nor _67184_ (_15632_, _07800_, _15627_);
  or _67185_ (_15633_, _15632_, _08469_);
  or _67186_ (_15634_, _15633_, _15631_);
  nand _67187_ (_15635_, _08469_, _07751_);
  and _67188_ (_15636_, _15635_, _08473_);
  and _67189_ (_15637_, _15636_, _15634_);
  nand _67190_ (_15638_, _12400_, _08480_);
  and _67191_ (_15640_, _15638_, _08479_);
  or _67192_ (_15641_, _15640_, _15637_);
  and _67193_ (_15642_, _15641_, _15398_);
  or _67194_ (_15643_, _15642_, _03758_);
  nor _67195_ (_15644_, _12272_, _07918_);
  nor _67196_ (_15645_, _15644_, _15400_);
  nand _67197_ (_15646_, _15645_, _03758_);
  and _67198_ (_15647_, _15646_, _07830_);
  and _67199_ (_15648_, _15647_, _15643_);
  and _67200_ (_15649_, _07894_, _07879_);
  nor _67201_ (_15651_, _15649_, _07895_);
  and _67202_ (_15652_, _15651_, _08490_);
  or _67203_ (_15653_, _15652_, _07825_);
  or _67204_ (_15654_, _15653_, _15648_);
  and _67205_ (_15655_, _15654_, _15397_);
  or _67206_ (_15656_, _15655_, _03765_);
  and _67207_ (_15657_, _08538_, _08261_);
  nor _67208_ (_15658_, _15657_, _08539_);
  or _67209_ (_15659_, _15658_, _03766_);
  and _67210_ (_15660_, _15659_, _08557_);
  and _67211_ (_15662_, _15660_, _15656_);
  and _67212_ (_15663_, _08568_, _08326_);
  nor _67213_ (_15664_, _15663_, _08569_);
  and _67214_ (_15665_, _15664_, _08523_);
  or _67215_ (_15666_, _15665_, _08555_);
  or _67216_ (_15667_, _15666_, _15662_);
  nand _67217_ (_15668_, _08555_, _03233_);
  and _67218_ (_15669_, _15668_, _07780_);
  and _67219_ (_15670_, _15669_, _15667_);
  and _67220_ (_15671_, _07808_, _07802_);
  nor _67221_ (_15672_, _15671_, _07809_);
  and _67222_ (_15673_, _15672_, _15069_);
  or _67223_ (_15674_, _15673_, _15670_);
  and _67224_ (_15675_, _15674_, _07732_);
  and _67225_ (_15676_, _07759_, _07753_);
  nor _67226_ (_15677_, _15676_, _07760_);
  and _67227_ (_15678_, _15677_, _07731_);
  or _67228_ (_15679_, _15678_, _03524_);
  or _67229_ (_15680_, _15679_, _15675_);
  and _67230_ (_15681_, _15680_, _15394_);
  and _67231_ (_15683_, _08668_, _08662_);
  nor _67232_ (_15684_, _15683_, _08669_);
  and _67233_ (_15685_, _15684_, _08597_);
  or _67234_ (_15686_, _15685_, _07729_);
  or _67235_ (_15687_, _15686_, _15681_);
  and _67236_ (_15688_, _15687_, _15390_);
  or _67237_ (_15689_, _15688_, _03790_);
  nand _67238_ (_15690_, _15424_, _03790_);
  and _67239_ (_15691_, _15690_, _08688_);
  and _67240_ (_15692_, _15691_, _15689_);
  and _67241_ (_15694_, _07954_, _03321_);
  nor _67242_ (_15695_, _08693_, _07506_);
  or _67243_ (_15696_, _15695_, _15694_);
  nor _67244_ (_15697_, _15696_, _08692_);
  nor _67245_ (_15698_, _15697_, _10828_);
  or _67246_ (_15699_, _15698_, _15692_);
  nand _67247_ (_15700_, _08692_, _07500_);
  and _67248_ (_15701_, _15700_, _03152_);
  and _67249_ (_15702_, _15701_, _15699_);
  nor _67250_ (_15703_, _15456_, _03152_);
  or _67251_ (_15705_, _15703_, _03520_);
  or _67252_ (_15706_, _15705_, _15702_);
  and _67253_ (_15707_, _12456_, _05227_);
  nor _67254_ (_15708_, _15707_, _15400_);
  nand _67255_ (_15709_, _15708_, _03520_);
  and _67256_ (_15710_, _15709_, _08710_);
  and _67257_ (_15711_, _15710_, _15706_);
  and _67258_ (_15712_, _08717_, \oc8051_golden_model_1.ACC [2]);
  nor _67259_ (_15713_, _08717_, \oc8051_golden_model_1.ACC [2]);
  nor _67260_ (_15714_, _15713_, _15712_);
  nor _67261_ (_15716_, _15714_, _08716_);
  nor _67262_ (_15717_, _15716_, _10851_);
  or _67263_ (_15718_, _15717_, _15711_);
  nand _67264_ (_15719_, _08716_, _07500_);
  and _67265_ (_15720_, _15719_, _42963_);
  and _67266_ (_15721_, _15720_, _15718_);
  or _67267_ (_15722_, _15721_, _15389_);
  and _67268_ (_43205_, _15722_, _41755_);
  nor _67269_ (_15723_, _42963_, _07500_);
  nor _67270_ (_15724_, _07795_, _07797_);
  nor _67271_ (_15726_, _15724_, _07810_);
  and _67272_ (_15727_, _15724_, _07810_);
  nor _67273_ (_15728_, _15727_, _15726_);
  nand _67274_ (_15729_, _15728_, _15069_);
  nor _67275_ (_15730_, _05227_, _07500_);
  nor _67276_ (_15731_, _12597_, _07918_);
  nor _67277_ (_15732_, _15731_, _15730_);
  nor _67278_ (_15733_, _15732_, _03759_);
  or _67279_ (_15734_, _12602_, _07911_);
  and _67280_ (_15735_, _15734_, _07910_);
  and _67281_ (_15737_, _03650_, _03191_);
  not _67282_ (_15738_, _15737_);
  nor _67283_ (_15739_, _03665_, _10544_);
  not _67284_ (_15740_, _15739_);
  or _67285_ (_15741_, _07777_, _10544_);
  and _67286_ (_15742_, _15741_, _15740_);
  nor _67287_ (_15743_, _15742_, _07798_);
  and _67288_ (_15744_, _12598_, _05227_);
  nor _67289_ (_15745_, _15744_, _15730_);
  nand _67290_ (_15746_, _15745_, _03636_);
  nor _67291_ (_15748_, _07746_, _07748_);
  or _67292_ (_15749_, _15748_, _04126_);
  and _67293_ (_15750_, _08397_, _15269_);
  or _67294_ (_15751_, _15750_, _15724_);
  nand _67295_ (_15752_, _03432_, _03231_);
  nor _67296_ (_15753_, _07918_, _04843_);
  nor _67297_ (_15754_, _15753_, _15730_);
  nand _67298_ (_15755_, _15754_, _07314_);
  and _67299_ (_15756_, _03877_, \oc8051_golden_model_1.ACC [2]);
  nor _67300_ (_15757_, _15525_, _15756_);
  nor _67301_ (_15759_, _10392_, _15757_);
  and _67302_ (_15760_, _10392_, _15757_);
  nor _67303_ (_15761_, _15760_, _15759_);
  and _67304_ (_15762_, _15761_, \oc8051_golden_model_1.PSW [7]);
  nor _67305_ (_15763_, _15761_, \oc8051_golden_model_1.PSW [7]);
  nor _67306_ (_15764_, _15763_, _15762_);
  and _67307_ (_15765_, _15764_, _15531_);
  nor _67308_ (_15766_, _15764_, _15531_);
  nor _67309_ (_15767_, _15766_, _15765_);
  or _67310_ (_15768_, _15767_, _08109_);
  nor _67311_ (_15770_, _05792_, _07500_);
  and _67312_ (_15771_, _12490_, _05792_);
  and _67313_ (_15772_, _15771_, _12507_);
  nor _67314_ (_15773_, _15772_, _15770_);
  nor _67315_ (_15774_, _15773_, _03506_);
  nand _67316_ (_15775_, _07928_, _04843_);
  nand _67317_ (_15776_, _07933_, _04843_);
  nor _67318_ (_15777_, _04012_, _07500_);
  and _67319_ (_15778_, _04012_, _07500_);
  or _67320_ (_15779_, _15778_, _15777_);
  or _67321_ (_15781_, _15779_, _07933_);
  and _67322_ (_15782_, _15781_, _07936_);
  and _67323_ (_15783_, _15782_, _15776_);
  and _67324_ (_15784_, _15783_, _05847_);
  or _67325_ (_15785_, _15784_, _06717_);
  or _67326_ (_15786_, _15783_, _07935_);
  and _67327_ (_15787_, _15786_, _03208_);
  or _67328_ (_15788_, _15787_, _04438_);
  and _67329_ (_15789_, _15788_, _04444_);
  and _67330_ (_15790_, _15789_, _15785_);
  nor _67331_ (_15792_, _12486_, _07918_);
  nor _67332_ (_15793_, _15792_, _15730_);
  nor _67333_ (_15794_, _15793_, _04444_);
  or _67334_ (_15795_, _15794_, _07948_);
  or _67335_ (_15796_, _15795_, _15790_);
  not _67336_ (_15797_, \oc8051_golden_model_1.PSW [6]);
  nor _67337_ (_15798_, _07954_, _15797_);
  nor _67338_ (_15799_, _15798_, \oc8051_golden_model_1.ACC [3]);
  nor _67339_ (_15800_, _15799_, _07955_);
  or _67340_ (_15801_, _15800_, _11538_);
  and _67341_ (_15803_, _15801_, _15796_);
  or _67342_ (_15804_, _15803_, _03516_);
  nor _67343_ (_15805_, _15771_, _15770_);
  nand _67344_ (_15806_, _15805_, _03516_);
  and _67345_ (_15807_, _15806_, _03983_);
  and _67346_ (_15808_, _15807_, _15804_);
  nor _67347_ (_15809_, _15754_, _03983_);
  or _67348_ (_15810_, _15809_, _07928_);
  or _67349_ (_15811_, _15810_, _15808_);
  and _67350_ (_15812_, _15811_, _15775_);
  or _67351_ (_15814_, _15812_, _04458_);
  or _67352_ (_15815_, _06717_, _07987_);
  and _67353_ (_15816_, _15815_, _03583_);
  and _67354_ (_15817_, _15816_, _15814_);
  nor _67355_ (_15818_, _08143_, _03583_);
  or _67356_ (_15819_, _15818_, _07991_);
  or _67357_ (_15820_, _15819_, _15817_);
  nand _67358_ (_15821_, _07991_, _05834_);
  and _67359_ (_15822_, _15821_, _15820_);
  or _67360_ (_15823_, _15822_, _03512_);
  and _67361_ (_15825_, _12500_, _05792_);
  nor _67362_ (_15826_, _15825_, _15770_);
  nand _67363_ (_15827_, _15826_, _03512_);
  and _67364_ (_15828_, _15827_, _03506_);
  and _67365_ (_15829_, _15828_, _15823_);
  or _67366_ (_15830_, _15829_, _15774_);
  and _67367_ (_15831_, _15830_, _06800_);
  nor _67368_ (_15832_, _07272_, _07270_);
  nor _67369_ (_15833_, _15832_, _07273_);
  and _67370_ (_15834_, _15833_, _06794_);
  or _67371_ (_15836_, _15834_, _11700_);
  or _67372_ (_15837_, _15836_, _15831_);
  and _67373_ (_15838_, _05026_, \oc8051_golden_model_1.ACC [2]);
  nor _67374_ (_15839_, _15474_, _15838_);
  and _67375_ (_15840_, _15839_, _15724_);
  nor _67376_ (_15841_, _15839_, _15724_);
  or _67377_ (_15842_, _15841_, _15840_);
  nor _67378_ (_15843_, _15842_, _07888_);
  and _67379_ (_15844_, _15842_, _07888_);
  nor _67380_ (_15845_, _15844_, _15843_);
  and _67381_ (_15847_, _15845_, _15480_);
  nor _67382_ (_15848_, _15845_, _15480_);
  nor _67383_ (_15849_, _15848_, _15847_);
  and _67384_ (_15850_, _15849_, _11706_);
  or _67385_ (_15851_, _15850_, _07922_);
  and _67386_ (_15852_, _15851_, _15837_);
  and _67387_ (_15853_, _15849_, _11705_);
  or _67388_ (_15854_, _15853_, _08035_);
  or _67389_ (_15855_, _15854_, _15852_);
  and _67390_ (_15856_, _06569_, \oc8051_golden_model_1.ACC [2]);
  nor _67391_ (_15858_, _15492_, _15856_);
  nor _67392_ (_15859_, _15858_, _15748_);
  and _67393_ (_15860_, _15858_, _15748_);
  nor _67394_ (_15861_, _15860_, _15859_);
  and _67395_ (_15862_, _15861_, \oc8051_golden_model_1.PSW [7]);
  nor _67396_ (_15863_, _15861_, \oc8051_golden_model_1.PSW [7]);
  nor _67397_ (_15864_, _15863_, _15862_);
  and _67398_ (_15865_, _15864_, _15499_);
  nor _67399_ (_15866_, _15864_, _15499_);
  or _67400_ (_15867_, _15866_, _15865_);
  nand _67401_ (_15869_, _15867_, _08035_);
  and _67402_ (_15870_, _15869_, _03619_);
  and _67403_ (_15871_, _15870_, _15855_);
  and _67404_ (_15872_, _10377_, \oc8051_golden_model_1.PSW [7]);
  nor _67405_ (_15873_, _15510_, _08619_);
  nor _67406_ (_15874_, _10371_, _15873_);
  and _67407_ (_15875_, _10371_, _15873_);
  or _67408_ (_15876_, _15875_, _15874_);
  not _67409_ (_15877_, _15515_);
  and _67410_ (_15878_, _15877_, _15876_);
  nor _67411_ (_15880_, _15878_, _15872_);
  nor _67412_ (_15881_, _15880_, _03619_);
  or _67413_ (_15882_, _15881_, _08108_);
  or _67414_ (_15883_, _15882_, _15871_);
  and _67415_ (_15884_, _15883_, _15768_);
  or _67416_ (_15885_, _15884_, _03311_);
  nand _67417_ (_15886_, _03432_, _03311_);
  and _67418_ (_15887_, _15886_, _03500_);
  and _67419_ (_15888_, _15887_, _15885_);
  nor _67420_ (_15889_, _12525_, _08358_);
  nor _67421_ (_15891_, _15889_, _15770_);
  nor _67422_ (_15892_, _15891_, _03500_);
  or _67423_ (_15893_, _15892_, _07314_);
  or _67424_ (_15894_, _15893_, _15888_);
  and _67425_ (_15895_, _15894_, _15755_);
  or _67426_ (_15896_, _15895_, _03479_);
  and _67427_ (_15897_, _06717_, _05227_);
  nor _67428_ (_15898_, _15897_, _15730_);
  nand _67429_ (_15899_, _15898_, _03479_);
  and _67430_ (_15900_, _15899_, _03474_);
  and _67431_ (_15902_, _15900_, _15896_);
  nor _67432_ (_15903_, _12583_, _07918_);
  nor _67433_ (_15904_, _15903_, _15730_);
  nor _67434_ (_15905_, _15904_, _03474_);
  or _67435_ (_15906_, _15905_, _07328_);
  or _67436_ (_15907_, _15906_, _15902_);
  or _67437_ (_15908_, _07466_, _07677_);
  and _67438_ (_15909_, _15908_, _15907_);
  or _67439_ (_15910_, _15909_, _03231_);
  and _67440_ (_15911_, _15910_, _15752_);
  or _67441_ (_15913_, _15911_, _03437_);
  and _67442_ (_15914_, _05227_, _06217_);
  nor _67443_ (_15915_, _15914_, _15730_);
  nand _67444_ (_15916_, _15915_, _03437_);
  and _67445_ (_15917_, _15916_, _08386_);
  and _67446_ (_15918_, _15917_, _15913_);
  or _67447_ (_15919_, _08386_, _03432_);
  nand _67448_ (_15920_, _15919_, _15750_);
  or _67449_ (_15921_, _15920_, _15918_);
  nand _67450_ (_15922_, _15921_, _15751_);
  and _67451_ (_15924_, _15922_, _15588_);
  nor _67452_ (_15925_, _15724_, _15588_);
  or _67453_ (_15926_, _15925_, _14990_);
  nor _67454_ (_15927_, _15926_, _15924_);
  or _67455_ (_15928_, _15748_, _03043_);
  and _67456_ (_15929_, _15928_, _08405_);
  or _67457_ (_15930_, _15929_, _15927_);
  and _67458_ (_15931_, _15930_, _15749_);
  or _67459_ (_15932_, _15931_, _03767_);
  or _67460_ (_15933_, _12604_, _03768_);
  and _67461_ (_15935_, _15933_, _08416_);
  and _67462_ (_15936_, _15935_, _15932_);
  and _67463_ (_15937_, _08415_, _10392_);
  or _67464_ (_15938_, _15937_, _03636_);
  or _67465_ (_15939_, _15938_, _15936_);
  and _67466_ (_15940_, _15939_, _15746_);
  or _67467_ (_15941_, _15940_, _03769_);
  or _67468_ (_15942_, _15730_, _04501_);
  and _67469_ (_15943_, _15942_, _15742_);
  and _67470_ (_15944_, _15943_, _15941_);
  or _67471_ (_15946_, _15944_, _15743_);
  and _67472_ (_15947_, _15946_, _15738_);
  and _67473_ (_15948_, _07797_, _15737_);
  or _67474_ (_15949_, _15948_, _15947_);
  and _67475_ (_15950_, _15949_, _08446_);
  and _67476_ (_15951_, _08445_, _07748_);
  or _67477_ (_15952_, _15951_, _03755_);
  or _67478_ (_15953_, _15952_, _15950_);
  and _67479_ (_15954_, _15953_, _15735_);
  and _67480_ (_15955_, _08657_, _07909_);
  or _67481_ (_15957_, _15955_, _15954_);
  and _67482_ (_15958_, _15957_, _05769_);
  or _67483_ (_15959_, _15915_, _12603_);
  nor _67484_ (_15960_, _15959_, _04505_);
  or _67485_ (_15961_, _15960_, _15622_);
  or _67486_ (_15962_, _15961_, _15958_);
  nand _67487_ (_15963_, _15622_, _07795_);
  and _67488_ (_15964_, _15963_, _15627_);
  and _67489_ (_15965_, _15964_, _15962_);
  nor _67490_ (_15966_, _07795_, _15627_);
  or _67491_ (_15968_, _15966_, _08469_);
  or _67492_ (_15969_, _15968_, _15965_);
  nand _67493_ (_15970_, _08469_, _07746_);
  and _67494_ (_15971_, _15970_, _08473_);
  and _67495_ (_15972_, _15971_, _15969_);
  nand _67496_ (_15973_, _12603_, _08480_);
  and _67497_ (_15974_, _15973_, _08479_);
  or _67498_ (_15975_, _15974_, _15972_);
  nand _67499_ (_15976_, _08477_, _08658_);
  and _67500_ (_15977_, _15976_, _03759_);
  and _67501_ (_15979_, _15977_, _15975_);
  or _67502_ (_15980_, _15979_, _15733_);
  and _67503_ (_15981_, _15980_, _07830_);
  and _67504_ (_15982_, _07896_, _07873_);
  nor _67505_ (_15983_, _15982_, _07897_);
  and _67506_ (_15984_, _15983_, _08490_);
  or _67507_ (_15985_, _15984_, _07825_);
  or _67508_ (_15986_, _15985_, _15981_);
  and _67509_ (_15987_, _08508_, _08074_);
  nor _67510_ (_15988_, _15987_, _08509_);
  or _67511_ (_15990_, _15988_, _08495_);
  and _67512_ (_15991_, _15990_, _03766_);
  and _67513_ (_15992_, _15991_, _15986_);
  and _67514_ (_15993_, _08540_, _08256_);
  nor _67515_ (_15994_, _15993_, _08541_);
  and _67516_ (_15995_, _15994_, _03765_);
  or _67517_ (_15996_, _15995_, _08523_);
  or _67518_ (_15997_, _15996_, _15992_);
  and _67519_ (_15998_, _08570_, _08321_);
  nor _67520_ (_15999_, _15998_, _08571_);
  or _67521_ (_16001_, _15999_, _08557_);
  and _67522_ (_16002_, _16001_, _08556_);
  and _67523_ (_16003_, _16002_, _15997_);
  nand _67524_ (_16004_, _08555_, \oc8051_golden_model_1.ACC [2]);
  nand _67525_ (_16005_, _16004_, _07780_);
  or _67526_ (_16006_, _16005_, _16003_);
  and _67527_ (_16007_, _16006_, _15729_);
  or _67528_ (_16008_, _16007_, _07731_);
  nor _67529_ (_16009_, _15748_, _07761_);
  and _67530_ (_16010_, _15748_, _07761_);
  nor _67531_ (_16012_, _16010_, _16009_);
  nand _67532_ (_16013_, _16012_, _07731_);
  and _67533_ (_16014_, _16013_, _03526_);
  and _67534_ (_16015_, _16014_, _16008_);
  nor _67535_ (_16016_, _08631_, _10371_);
  and _67536_ (_16017_, _08631_, _10371_);
  nor _67537_ (_16018_, _16017_, _16016_);
  and _67538_ (_16019_, _16018_, _03524_);
  or _67539_ (_16020_, _16019_, _08597_);
  or _67540_ (_16021_, _16020_, _16015_);
  nor _67541_ (_16023_, _08670_, _10392_);
  and _67542_ (_16024_, _08670_, _10392_);
  nor _67543_ (_16025_, _16024_, _16023_);
  nand _67544_ (_16026_, _16025_, _08597_);
  and _67545_ (_16027_, _16026_, _10803_);
  and _67546_ (_16028_, _16027_, _16021_);
  and _67547_ (_16029_, _07729_, \oc8051_golden_model_1.ACC [2]);
  or _67548_ (_16030_, _16029_, _03790_);
  or _67549_ (_16031_, _16030_, _16028_);
  nand _67550_ (_16032_, _15793_, _03790_);
  and _67551_ (_16034_, _16032_, _08688_);
  and _67552_ (_16035_, _16034_, _16031_);
  nor _67553_ (_16036_, _15694_, _07500_);
  or _67554_ (_16037_, _16036_, _08694_);
  and _67555_ (_16038_, _16037_, _08687_);
  or _67556_ (_16039_, _16038_, _08692_);
  or _67557_ (_16040_, _16039_, _16035_);
  nand _67558_ (_16041_, _08692_, _07405_);
  and _67559_ (_16042_, _16041_, _03152_);
  and _67560_ (_16043_, _16042_, _16040_);
  nor _67561_ (_16045_, _15826_, _03152_);
  or _67562_ (_16046_, _16045_, _03520_);
  or _67563_ (_16047_, _16046_, _16043_);
  and _67564_ (_16048_, _12658_, _05227_);
  nor _67565_ (_16049_, _16048_, _15730_);
  nand _67566_ (_16050_, _16049_, _03520_);
  and _67567_ (_16051_, _16050_, _08710_);
  and _67568_ (_16052_, _16051_, _16047_);
  or _67569_ (_16053_, _15712_, \oc8051_golden_model_1.ACC [3]);
  and _67570_ (_16054_, _16053_, _08718_);
  and _67571_ (_16056_, _16054_, _08709_);
  or _67572_ (_16057_, _16056_, _08716_);
  or _67573_ (_16058_, _16057_, _16052_);
  nand _67574_ (_16059_, _08716_, _07405_);
  and _67575_ (_16060_, _16059_, _42963_);
  and _67576_ (_16061_, _16060_, _16058_);
  or _67577_ (_16062_, _16061_, _15723_);
  and _67578_ (_43206_, _16062_, _41755_);
  nor _67579_ (_16063_, _42963_, _07405_);
  nand _67580_ (_16064_, _07729_, _07500_);
  nand _67581_ (_16066_, _08555_, _07500_);
  nor _67582_ (_16067_, _08542_, _08530_);
  nor _67583_ (_16068_, _16067_, _08543_);
  or _67584_ (_16069_, _16068_, _03766_);
  and _67585_ (_16070_, _16069_, _08557_);
  nand _67586_ (_16071_, _08469_, _07744_);
  nand _67587_ (_16072_, _08458_, _07793_);
  or _67588_ (_16073_, _12842_, _07911_);
  and _67589_ (_16074_, _16073_, _07910_);
  and _67590_ (_16075_, _14871_, _07792_);
  nor _67591_ (_16077_, _05227_, _07405_);
  and _67592_ (_16078_, _12711_, _05227_);
  nor _67593_ (_16079_, _16078_, _16077_);
  nand _67594_ (_16080_, _16079_, _03636_);
  or _67595_ (_16081_, _08406_, _07745_);
  nand _67596_ (_16082_, _04249_, _03231_);
  nor _67597_ (_16083_, _05712_, _07918_);
  nor _67598_ (_16084_, _16083_, _16077_);
  nand _67599_ (_16085_, _16084_, _07314_);
  or _67600_ (_16086_, _15873_, _10369_);
  and _67601_ (_16088_, _16086_, _11474_);
  nor _67602_ (_16089_, _08615_, _16088_);
  and _67603_ (_16090_, _08615_, _16088_);
  nor _67604_ (_16091_, _16090_, _16089_);
  not _67605_ (_16092_, _15872_);
  nor _67606_ (_16093_, _16092_, _16091_);
  and _67607_ (_16094_, _16092_, _16091_);
  nor _67608_ (_16095_, _16094_, _16093_);
  nand _67609_ (_16096_, _16095_, _03614_);
  and _67610_ (_16097_, _16096_, _08109_);
  nand _67611_ (_16099_, _07928_, _05712_);
  nand _67612_ (_16100_, _07933_, _05712_);
  nor _67613_ (_16101_, _04012_, _07405_);
  and _67614_ (_16102_, _04012_, _07405_);
  or _67615_ (_16103_, _16102_, _16101_);
  or _67616_ (_16104_, _16103_, _07933_);
  and _67617_ (_16105_, _16104_, _07936_);
  and _67618_ (_16106_, _16105_, _16100_);
  and _67619_ (_16107_, _07935_, _06722_);
  or _67620_ (_16108_, _16107_, _16106_);
  and _67621_ (_16110_, _16108_, _07946_);
  nor _67622_ (_16111_, _12733_, _07918_);
  nor _67623_ (_16112_, _16111_, _16077_);
  nor _67624_ (_16113_, _16112_, _04444_);
  or _67625_ (_16114_, _16113_, _07948_);
  or _67626_ (_16115_, _16114_, _16110_);
  nor _67627_ (_16116_, _07955_, \oc8051_golden_model_1.ACC [4]);
  nor _67628_ (_16117_, _16116_, _07961_);
  not _67629_ (_16118_, _16117_);
  nand _67630_ (_16119_, _16118_, _07948_);
  and _67631_ (_16121_, _16119_, _03576_);
  and _67632_ (_16122_, _16121_, _16115_);
  nor _67633_ (_16123_, _05792_, _07405_);
  and _67634_ (_16124_, _12737_, _05792_);
  nor _67635_ (_16125_, _16124_, _16123_);
  nor _67636_ (_16126_, _16125_, _03517_);
  nor _67637_ (_16127_, _16084_, _03983_);
  or _67638_ (_16128_, _16127_, _07928_);
  or _67639_ (_16129_, _16128_, _16126_);
  or _67640_ (_16130_, _16129_, _16122_);
  and _67641_ (_16132_, _16130_, _16099_);
  or _67642_ (_16133_, _16132_, _04458_);
  or _67643_ (_16134_, _06722_, _07987_);
  and _67644_ (_16135_, _16134_, _03583_);
  and _67645_ (_16136_, _16135_, _16133_);
  nor _67646_ (_16137_, _08222_, _03583_);
  or _67647_ (_16138_, _16137_, _07991_);
  or _67648_ (_16139_, _16138_, _16136_);
  nand _67649_ (_16140_, _07991_, _03321_);
  and _67650_ (_16141_, _16140_, _16139_);
  or _67651_ (_16143_, _16141_, _03512_);
  and _67652_ (_16144_, _12718_, _05792_);
  nor _67653_ (_16145_, _16144_, _16123_);
  nand _67654_ (_16146_, _16145_, _03512_);
  and _67655_ (_16147_, _16146_, _03506_);
  and _67656_ (_16148_, _16147_, _16143_);
  and _67657_ (_16149_, _16124_, _12752_);
  nor _67658_ (_16150_, _16149_, _16123_);
  nor _67659_ (_16151_, _16150_, _03506_);
  or _67660_ (_16152_, _16151_, _06794_);
  or _67661_ (_16154_, _16152_, _16148_);
  nor _67662_ (_16155_, _07275_, _07273_);
  nor _67663_ (_16156_, _16155_, _07276_);
  or _67664_ (_16157_, _16156_, _06800_);
  and _67665_ (_16158_, _16157_, _16154_);
  or _67666_ (_16159_, _16158_, _07923_);
  or _67667_ (_16160_, _15847_, _15843_);
  nor _67668_ (_16161_, _04843_, \oc8051_golden_model_1.ACC [3]);
  nand _67669_ (_16162_, _04843_, \oc8051_golden_model_1.ACC [3]);
  and _67670_ (_16163_, _15839_, _16162_);
  or _67671_ (_16165_, _16163_, _16161_);
  nor _67672_ (_16166_, _16165_, _07794_);
  and _67673_ (_16167_, _16165_, _07794_);
  nor _67674_ (_16168_, _16167_, _16166_);
  and _67675_ (_16169_, _16168_, \oc8051_golden_model_1.PSW [7]);
  nor _67676_ (_16170_, _16168_, \oc8051_golden_model_1.PSW [7]);
  nor _67677_ (_16171_, _16170_, _16169_);
  and _67678_ (_16172_, _16171_, _16160_);
  nor _67679_ (_16173_, _16171_, _16160_);
  nor _67680_ (_16174_, _16173_, _16172_);
  or _67681_ (_16176_, _16174_, _07922_);
  and _67682_ (_16177_, _16176_, _16159_);
  or _67683_ (_16178_, _16177_, _08035_);
  or _67684_ (_16179_, _15865_, _15862_);
  and _67685_ (_16180_, _06717_, _07500_);
  or _67686_ (_16181_, _06717_, _07500_);
  and _67687_ (_16182_, _15858_, _16181_);
  or _67688_ (_16183_, _16182_, _16180_);
  nor _67689_ (_16184_, _16183_, _07745_);
  and _67690_ (_16185_, _16183_, _07745_);
  nor _67691_ (_16187_, _16185_, _16184_);
  and _67692_ (_16188_, _16187_, \oc8051_golden_model_1.PSW [7]);
  nor _67693_ (_16189_, _16187_, \oc8051_golden_model_1.PSW [7]);
  nor _67694_ (_16190_, _16189_, _16188_);
  and _67695_ (_16191_, _16190_, _16179_);
  nor _67696_ (_16192_, _16190_, _16179_);
  nor _67697_ (_16193_, _16192_, _16191_);
  or _67698_ (_16194_, _16193_, _08037_);
  and _67699_ (_16195_, _16194_, _16178_);
  or _67700_ (_16196_, _16195_, _03614_);
  and _67701_ (_16198_, _16196_, _16097_);
  or _67702_ (_16199_, _15765_, _15762_);
  or _67703_ (_16200_, _15757_, _11497_);
  and _67704_ (_16201_, _16200_, _11496_);
  nor _67705_ (_16202_, _08656_, _16201_);
  and _67706_ (_16203_, _08656_, _16201_);
  nor _67707_ (_16204_, _16203_, _16202_);
  and _67708_ (_16205_, _16204_, \oc8051_golden_model_1.PSW [7]);
  nor _67709_ (_16206_, _16204_, \oc8051_golden_model_1.PSW [7]);
  nor _67710_ (_16207_, _16206_, _16205_);
  and _67711_ (_16209_, _16207_, _16199_);
  nor _67712_ (_16210_, _16207_, _16199_);
  nor _67713_ (_16211_, _16210_, _16209_);
  and _67714_ (_16212_, _16211_, _08108_);
  or _67715_ (_16213_, _16212_, _03311_);
  or _67716_ (_16214_, _16213_, _16198_);
  nand _67717_ (_16215_, _04249_, _03311_);
  and _67718_ (_16216_, _16215_, _03500_);
  and _67719_ (_16217_, _16216_, _16214_);
  nor _67720_ (_16218_, _12716_, _08358_);
  nor _67721_ (_16220_, _16218_, _16123_);
  nor _67722_ (_16221_, _16220_, _03500_);
  or _67723_ (_16222_, _16221_, _07314_);
  or _67724_ (_16223_, _16222_, _16217_);
  and _67725_ (_16224_, _16223_, _16085_);
  or _67726_ (_16225_, _16224_, _03479_);
  and _67727_ (_16226_, _06722_, _05227_);
  nor _67728_ (_16227_, _16226_, _16077_);
  nand _67729_ (_16228_, _16227_, _03479_);
  and _67730_ (_16229_, _16228_, _03474_);
  and _67731_ (_16231_, _16229_, _16225_);
  nor _67732_ (_16232_, _12827_, _07918_);
  nor _67733_ (_16233_, _16232_, _16077_);
  nor _67734_ (_16234_, _16233_, _03474_);
  or _67735_ (_16235_, _16234_, _07328_);
  or _67736_ (_16236_, _16235_, _16231_);
  or _67737_ (_16237_, _07412_, _07677_);
  and _67738_ (_16238_, _16237_, _16236_);
  or _67739_ (_16239_, _16238_, _03231_);
  and _67740_ (_16240_, _16239_, _16082_);
  or _67741_ (_16242_, _16240_, _03437_);
  and _67742_ (_16243_, _06233_, _05227_);
  nor _67743_ (_16244_, _16243_, _16077_);
  nand _67744_ (_16245_, _16244_, _03437_);
  and _67745_ (_16246_, _16245_, _08386_);
  and _67746_ (_16247_, _16246_, _16242_);
  nor _67747_ (_16248_, _08386_, _04249_);
  or _67748_ (_16249_, _16248_, _16247_);
  nor _67749_ (_16250_, _04325_, _03932_);
  and _67750_ (_16251_, _16250_, _03936_);
  nor _67751_ (_16253_, _07827_, _04121_);
  not _67752_ (_16254_, _16253_);
  and _67753_ (_16255_, _16254_, _16251_);
  and _67754_ (_16256_, _16255_, _16249_);
  not _67755_ (_16257_, _16255_);
  and _67756_ (_16258_, _16257_, _07794_);
  or _67757_ (_16259_, _16258_, _08405_);
  or _67758_ (_16260_, _16259_, _16256_);
  and _67759_ (_16261_, _16260_, _16081_);
  or _67760_ (_16262_, _16261_, _03767_);
  or _67761_ (_16264_, _12844_, _03768_);
  and _67762_ (_16265_, _16264_, _08416_);
  and _67763_ (_16266_, _16265_, _16262_);
  and _67764_ (_16267_, _08415_, _08656_);
  or _67765_ (_16268_, _16267_, _03636_);
  or _67766_ (_16269_, _16268_, _16266_);
  and _67767_ (_16270_, _16269_, _16080_);
  or _67768_ (_16271_, _16270_, _03769_);
  or _67769_ (_16272_, _16077_, _04501_);
  and _67770_ (_16273_, _16272_, _14870_);
  and _67771_ (_16275_, _16273_, _16271_);
  or _67772_ (_16276_, _16275_, _16075_);
  and _67773_ (_16277_, _16276_, _08446_);
  and _67774_ (_16278_, _08445_, _07743_);
  or _67775_ (_16279_, _16278_, _03755_);
  or _67776_ (_16280_, _16279_, _16277_);
  and _67777_ (_16281_, _16280_, _16074_);
  and _67778_ (_16282_, _08654_, _07909_);
  or _67779_ (_16283_, _16282_, _16281_);
  and _67780_ (_16284_, _16283_, _05769_);
  or _67781_ (_16286_, _16244_, _12843_);
  nor _67782_ (_16287_, _16286_, _04505_);
  or _67783_ (_16288_, _16287_, _08458_);
  or _67784_ (_16289_, _16288_, _16284_);
  and _67785_ (_16290_, _16289_, _16072_);
  or _67786_ (_16291_, _16290_, _08465_);
  nand _67787_ (_16292_, _08465_, _07793_);
  and _67788_ (_16293_, _16292_, _15029_);
  and _67789_ (_16294_, _16293_, _16291_);
  nor _67790_ (_16295_, _07793_, _15029_);
  or _67791_ (_16297_, _16295_, _08469_);
  or _67792_ (_16298_, _16297_, _16294_);
  and _67793_ (_16299_, _16298_, _16071_);
  or _67794_ (_16300_, _16299_, _03761_);
  nand _67795_ (_16301_, _12843_, _03761_);
  and _67796_ (_16302_, _16301_, _08480_);
  and _67797_ (_16303_, _16302_, _16300_);
  nor _67798_ (_16304_, _08480_, _08655_);
  or _67799_ (_16305_, _16304_, _03758_);
  or _67800_ (_16306_, _16305_, _16303_);
  nor _67801_ (_16308_, _12710_, _07918_);
  nor _67802_ (_16309_, _16308_, _16077_);
  nand _67803_ (_16310_, _16309_, _03758_);
  and _67804_ (_16311_, _16310_, _07830_);
  and _67805_ (_16312_, _16311_, _16306_);
  nor _67806_ (_16313_, _07898_, _07863_);
  nor _67807_ (_16314_, _16313_, _07899_);
  and _67808_ (_16315_, _16314_, _08490_);
  or _67809_ (_16316_, _16315_, _07825_);
  or _67810_ (_16317_, _16316_, _16312_);
  nor _67811_ (_16319_, _08510_, _08066_);
  nor _67812_ (_16320_, _16319_, _08511_);
  or _67813_ (_16321_, _16320_, _08495_);
  and _67814_ (_16322_, _16321_, _16317_);
  or _67815_ (_16323_, _16322_, _03765_);
  and _67816_ (_16324_, _16323_, _16070_);
  nor _67817_ (_16325_, _08572_, _08315_);
  nor _67818_ (_16326_, _16325_, _08573_);
  and _67819_ (_16327_, _16326_, _08523_);
  or _67820_ (_16328_, _16327_, _08555_);
  or _67821_ (_16330_, _16328_, _16324_);
  and _67822_ (_16331_, _16330_, _16066_);
  or _67823_ (_16332_, _16331_, _15069_);
  nor _67824_ (_16333_, _07812_, _07794_);
  nor _67825_ (_16334_, _16333_, _07813_);
  or _67826_ (_16335_, _16334_, _07780_);
  and _67827_ (_16336_, _16335_, _07732_);
  and _67828_ (_16337_, _16336_, _16332_);
  nor _67829_ (_16338_, _07763_, _07745_);
  nor _67830_ (_16339_, _16338_, _07764_);
  and _67831_ (_16341_, _16339_, _07731_);
  or _67832_ (_16342_, _16341_, _03524_);
  or _67833_ (_16343_, _16342_, _16337_);
  nor _67834_ (_16344_, _08633_, _08615_);
  nor _67835_ (_16345_, _16344_, _08634_);
  or _67836_ (_16346_, _16345_, _03526_);
  and _67837_ (_16347_, _16346_, _08598_);
  and _67838_ (_16348_, _16347_, _16343_);
  nor _67839_ (_16349_, _08672_, _08656_);
  nor _67840_ (_16350_, _16349_, _08673_);
  and _67841_ (_16352_, _16350_, _08597_);
  or _67842_ (_16353_, _16352_, _07729_);
  or _67843_ (_16354_, _16353_, _16348_);
  and _67844_ (_16355_, _16354_, _16064_);
  or _67845_ (_16356_, _16355_, _03790_);
  nand _67846_ (_16357_, _16112_, _03790_);
  and _67847_ (_16358_, _16357_, _08688_);
  and _67848_ (_16359_, _16358_, _16356_);
  and _67849_ (_16360_, _08694_, _07405_);
  nor _67850_ (_16361_, _08694_, _07405_);
  nor _67851_ (_16363_, _16361_, _16360_);
  not _67852_ (_16364_, _16363_);
  and _67853_ (_16365_, _16364_, _08687_);
  or _67854_ (_16366_, _16365_, _08692_);
  or _67855_ (_16367_, _16366_, _16359_);
  nand _67856_ (_16368_, _08692_, _07399_);
  and _67857_ (_16369_, _16368_, _03152_);
  and _67858_ (_16370_, _16369_, _16367_);
  nor _67859_ (_16371_, _16145_, _03152_);
  or _67860_ (_16372_, _16371_, _03520_);
  or _67861_ (_16374_, _16372_, _16370_);
  and _67862_ (_16375_, _12893_, _05227_);
  nor _67863_ (_16376_, _16375_, _16077_);
  nand _67864_ (_16377_, _16376_, _03520_);
  and _67865_ (_16378_, _16377_, _08710_);
  and _67866_ (_16379_, _16378_, _16374_);
  and _67867_ (_16380_, _08718_, _07405_);
  nor _67868_ (_16381_, _16380_, _08719_);
  and _67869_ (_16382_, _16381_, _08709_);
  or _67870_ (_16383_, _16382_, _08716_);
  or _67871_ (_16385_, _16383_, _16379_);
  nand _67872_ (_16386_, _08716_, _07399_);
  and _67873_ (_16387_, _16386_, _42963_);
  and _67874_ (_16388_, _16387_, _16385_);
  or _67875_ (_16389_, _16388_, _16063_);
  and _67876_ (_43207_, _16389_, _41755_);
  nor _67877_ (_16390_, _42963_, _07399_);
  and _67878_ (_16391_, _07900_, _07857_);
  nor _67879_ (_16392_, _16391_, _07901_);
  or _67880_ (_16393_, _16392_, _07830_);
  nand _67881_ (_16395_, _08469_, _07740_);
  nand _67882_ (_16396_, _08458_, _07788_);
  nor _67883_ (_16397_, _05227_, _07399_);
  and _67884_ (_16398_, _13036_, _05227_);
  nor _67885_ (_16399_, _16398_, _16397_);
  nand _67886_ (_16400_, _16399_, _03636_);
  or _67887_ (_16401_, _07741_, _04126_);
  and _67888_ (_16402_, _03633_, _03193_);
  and _67889_ (_16403_, _03655_, _03193_);
  not _67890_ (_16404_, _16403_);
  nor _67891_ (_16406_, _07790_, _07788_);
  or _67892_ (_16407_, _16406_, _16404_);
  nand _67893_ (_16408_, _03834_, _03231_);
  nor _67894_ (_16409_, _05422_, _07918_);
  nor _67895_ (_16410_, _16409_, _16397_);
  nand _67896_ (_16411_, _16410_, _07314_);
  and _67897_ (_16412_, _04249_, \oc8051_golden_model_1.ACC [4]);
  nor _67898_ (_16413_, _16202_, _16412_);
  nor _67899_ (_16414_, _08652_, _16413_);
  and _67900_ (_16415_, _08652_, _16413_);
  nor _67901_ (_16417_, _16415_, _16414_);
  and _67902_ (_16418_, _16417_, \oc8051_golden_model_1.PSW [7]);
  nor _67903_ (_16419_, _16417_, \oc8051_golden_model_1.PSW [7]);
  nor _67904_ (_16420_, _16419_, _16418_);
  nor _67905_ (_16421_, _16209_, _16205_);
  not _67906_ (_16422_, _16421_);
  and _67907_ (_16423_, _16422_, _16420_);
  nor _67908_ (_16424_, _16422_, _16420_);
  nor _67909_ (_16425_, _16424_, _16423_);
  or _67910_ (_16426_, _16425_, _08109_);
  not _67911_ (_16428_, _16406_);
  and _67912_ (_16429_, _05712_, \oc8051_golden_model_1.ACC [4]);
  nor _67913_ (_16430_, _16166_, _16429_);
  and _67914_ (_16431_, _16430_, _16428_);
  nor _67915_ (_16432_, _16430_, _16428_);
  nor _67916_ (_16433_, _16432_, _16431_);
  nor _67917_ (_16434_, _16433_, _07888_);
  and _67918_ (_16435_, _16433_, _07888_);
  nor _67919_ (_16436_, _16435_, _16434_);
  nor _67920_ (_16437_, _16172_, _16169_);
  not _67921_ (_16439_, _16437_);
  and _67922_ (_16440_, _16439_, _16436_);
  nor _67923_ (_16441_, _16439_, _16436_);
  nor _67924_ (_16442_, _16441_, _16440_);
  or _67925_ (_16443_, _16442_, _07922_);
  nor _67926_ (_16444_, _05792_, _07399_);
  and _67927_ (_16445_, _12934_, _05792_);
  and _67928_ (_16446_, _16445_, _12949_);
  nor _67929_ (_16447_, _16446_, _16444_);
  nor _67930_ (_16448_, _16447_, _03506_);
  nand _67931_ (_16450_, _07928_, _05422_);
  nand _67932_ (_16451_, _07933_, _05422_);
  nor _67933_ (_16452_, _04012_, _07399_);
  and _67934_ (_16453_, _04012_, _07399_);
  or _67935_ (_16454_, _16453_, _16452_);
  or _67936_ (_16455_, _16454_, _07933_);
  and _67937_ (_16456_, _16455_, _07936_);
  and _67938_ (_16457_, _16456_, _16451_);
  and _67939_ (_16458_, _07935_, _06721_);
  or _67940_ (_16459_, _16458_, _16457_);
  and _67941_ (_16461_, _16459_, _07946_);
  not _67942_ (_16462_, _16397_);
  or _67943_ (_16463_, _12930_, _07918_);
  and _67944_ (_16464_, _16463_, _16462_);
  nor _67945_ (_16465_, _16464_, _04444_);
  or _67946_ (_16466_, _16465_, _07948_);
  or _67947_ (_16467_, _16466_, _16461_);
  and _67948_ (_16468_, _11549_, _07963_);
  nor _67949_ (_16469_, _11549_, _07963_);
  nor _67950_ (_16470_, _16469_, _16468_);
  nand _67951_ (_16472_, _16470_, _07948_);
  and _67952_ (_16473_, _16472_, _03576_);
  and _67953_ (_16474_, _16473_, _16467_);
  nor _67954_ (_16475_, _16445_, _16444_);
  nor _67955_ (_16476_, _16475_, _03517_);
  nor _67956_ (_16477_, _16410_, _03983_);
  or _67957_ (_16478_, _16477_, _07928_);
  or _67958_ (_16479_, _16478_, _16476_);
  or _67959_ (_16480_, _16479_, _16474_);
  and _67960_ (_16481_, _16480_, _16450_);
  or _67961_ (_16483_, _16481_, _04458_);
  or _67962_ (_16484_, _06721_, _07987_);
  and _67963_ (_16485_, _16484_, _03583_);
  and _67964_ (_16486_, _16485_, _16483_);
  nor _67965_ (_16487_, _08205_, _03583_);
  or _67966_ (_16488_, _16487_, _07991_);
  or _67967_ (_16489_, _16488_, _16486_);
  nand _67968_ (_16490_, _07991_, _03233_);
  and _67969_ (_16491_, _16490_, _16489_);
  or _67970_ (_16492_, _16491_, _03512_);
  and _67971_ (_16494_, _12914_, _05792_);
  nor _67972_ (_16495_, _16494_, _16444_);
  nand _67973_ (_16496_, _16495_, _03512_);
  and _67974_ (_16497_, _16496_, _03506_);
  and _67975_ (_16498_, _16497_, _16492_);
  or _67976_ (_16499_, _16498_, _16448_);
  and _67977_ (_16500_, _16499_, _06800_);
  nor _67978_ (_16501_, _07278_, _07276_);
  nor _67979_ (_16502_, _16501_, _07279_);
  and _67980_ (_16503_, _16502_, _06794_);
  or _67981_ (_16505_, _16503_, _07923_);
  or _67982_ (_16506_, _16505_, _16500_);
  and _67983_ (_16507_, _16506_, _16443_);
  or _67984_ (_16508_, _16507_, _08035_);
  and _67985_ (_16509_, _06661_, \oc8051_golden_model_1.ACC [4]);
  nor _67986_ (_16510_, _16184_, _16509_);
  nor _67987_ (_16511_, _16510_, _07741_);
  and _67988_ (_16512_, _16510_, _07741_);
  nor _67989_ (_16513_, _16512_, _16511_);
  and _67990_ (_16514_, _16513_, \oc8051_golden_model_1.PSW [7]);
  nor _67991_ (_16516_, _16513_, \oc8051_golden_model_1.PSW [7]);
  nor _67992_ (_16517_, _16516_, _16514_);
  nor _67993_ (_16518_, _16191_, _16188_);
  not _67994_ (_16519_, _16518_);
  and _67995_ (_16520_, _16519_, _16517_);
  nor _67996_ (_16521_, _16519_, _16517_);
  nor _67997_ (_16522_, _16521_, _16520_);
  or _67998_ (_16523_, _16522_, _08037_);
  and _67999_ (_16524_, _16523_, _03619_);
  and _68000_ (_16525_, _16524_, _16508_);
  nor _68001_ (_16527_, _16089_, _08612_);
  nor _68002_ (_16528_, _08610_, _16527_);
  and _68003_ (_16529_, _08610_, _16527_);
  or _68004_ (_16530_, _16529_, _16528_);
  not _68005_ (_16531_, _16093_);
  nor _68006_ (_16532_, _16531_, _16530_);
  and _68007_ (_16533_, _16531_, _16530_);
  nor _68008_ (_16534_, _16533_, _16532_);
  nand _68009_ (_16535_, _16534_, _08109_);
  and _68010_ (_16536_, _16535_, _10431_);
  or _68011_ (_16538_, _16536_, _16525_);
  and _68012_ (_16539_, _16538_, _16426_);
  or _68013_ (_16540_, _16539_, _03311_);
  nand _68014_ (_16541_, _03834_, _03311_);
  and _68015_ (_16542_, _16541_, _03500_);
  and _68016_ (_16543_, _16542_, _16540_);
  nor _68017_ (_16544_, _12912_, _08358_);
  nor _68018_ (_16545_, _16544_, _16444_);
  nor _68019_ (_16546_, _16545_, _03500_);
  or _68020_ (_16547_, _16546_, _07314_);
  or _68021_ (_16549_, _16547_, _16543_);
  and _68022_ (_16550_, _16549_, _16411_);
  or _68023_ (_16551_, _16550_, _03479_);
  and _68024_ (_16552_, _06721_, _05227_);
  nor _68025_ (_16553_, _16552_, _16397_);
  nand _68026_ (_16554_, _16553_, _03479_);
  and _68027_ (_16555_, _16554_, _03474_);
  and _68028_ (_16556_, _16555_, _16551_);
  nor _68029_ (_16557_, _13021_, _07918_);
  nor _68030_ (_16558_, _16557_, _16397_);
  nor _68031_ (_16560_, _16558_, _03474_);
  or _68032_ (_16561_, _16560_, _07328_);
  or _68033_ (_16562_, _16561_, _16556_);
  or _68034_ (_16563_, _07382_, _07677_);
  and _68035_ (_16564_, _16563_, _16562_);
  or _68036_ (_16565_, _16564_, _03231_);
  and _68037_ (_16566_, _16565_, _16408_);
  or _68038_ (_16567_, _16566_, _03437_);
  and _68039_ (_16568_, _06211_, _05227_);
  nor _68040_ (_16569_, _16568_, _16397_);
  nand _68041_ (_16572_, _16569_, _03437_);
  and _68042_ (_16573_, _16572_, _08386_);
  and _68043_ (_16574_, _16573_, _16567_);
  nor _68044_ (_16575_, _08386_, _03834_);
  or _68045_ (_16576_, _16575_, _16403_);
  or _68046_ (_16577_, _16576_, _16574_);
  and _68047_ (_16578_, _16577_, _16407_);
  nor _68048_ (_16579_, _16578_, _16402_);
  and _68049_ (_16580_, _16428_, _04127_);
  nand _68050_ (_16581_, _03925_, _03193_);
  or _68051_ (_16583_, _16581_, _03043_);
  nand _68052_ (_16584_, _15270_, _16583_);
  or _68053_ (_16585_, _16584_, _16580_);
  nor _68054_ (_16586_, _16585_, _16579_);
  and _68055_ (_16587_, _16584_, _16406_);
  or _68056_ (_16588_, _16587_, _04129_);
  or _68057_ (_16589_, _16588_, _16586_);
  or _68058_ (_16590_, _16406_, _15588_);
  and _68059_ (_16591_, _16590_, _14991_);
  and _68060_ (_16592_, _16591_, _16589_);
  and _68061_ (_16594_, _08405_, _07741_);
  or _68062_ (_16595_, _16594_, _16592_);
  and _68063_ (_16596_, _16595_, _16401_);
  or _68064_ (_16597_, _16596_, _03767_);
  or _68065_ (_16598_, _13042_, _03768_);
  and _68066_ (_16599_, _16598_, _08416_);
  and _68067_ (_16600_, _16599_, _16597_);
  and _68068_ (_16601_, _08415_, _08652_);
  or _68069_ (_16602_, _16601_, _03636_);
  or _68070_ (_16603_, _16602_, _16600_);
  and _68071_ (_16605_, _16603_, _16400_);
  or _68072_ (_16606_, _16605_, _03769_);
  or _68073_ (_16607_, _16397_, _04501_);
  and _68074_ (_16608_, _16607_, _15741_);
  and _68075_ (_16609_, _16608_, _16606_);
  nor _68076_ (_16610_, _15741_, _07791_);
  or _68077_ (_16611_, _16610_, _16609_);
  and _68078_ (_16612_, _16611_, _15740_);
  and _68079_ (_16613_, _15739_, _07790_);
  or _68080_ (_16614_, _16613_, _16612_);
  and _68081_ (_16616_, _16614_, _15738_);
  and _68082_ (_16617_, _07790_, _15737_);
  or _68083_ (_16618_, _16617_, _16616_);
  and _68084_ (_16619_, _16618_, _08446_);
  and _68085_ (_16620_, _08445_, _07739_);
  or _68086_ (_16621_, _16620_, _03755_);
  or _68087_ (_16622_, _16621_, _16619_);
  or _68088_ (_16623_, _13040_, _07911_);
  and _68089_ (_16624_, _16623_, _07910_);
  and _68090_ (_16625_, _16624_, _16622_);
  and _68091_ (_16627_, _08650_, _07909_);
  or _68092_ (_16628_, _16627_, _16625_);
  and _68093_ (_16629_, _16628_, _05769_);
  or _68094_ (_16630_, _16569_, _13041_);
  nor _68095_ (_16631_, _16630_, _04505_);
  or _68096_ (_16632_, _16631_, _08458_);
  or _68097_ (_16633_, _16632_, _16629_);
  and _68098_ (_16634_, _16633_, _16396_);
  or _68099_ (_16635_, _16634_, _08465_);
  nor _68100_ (_16636_, _07788_, _04161_);
  or _68101_ (_16638_, _16636_, _08466_);
  and _68102_ (_16639_, _16638_, _16635_);
  nor _68103_ (_16640_, _07788_, _15029_);
  or _68104_ (_16641_, _16640_, _08469_);
  or _68105_ (_16642_, _16641_, _16639_);
  and _68106_ (_16643_, _16642_, _16395_);
  or _68107_ (_16644_, _16643_, _03761_);
  nand _68108_ (_16645_, _13041_, _03761_);
  and _68109_ (_16646_, _16645_, _08480_);
  and _68110_ (_16647_, _16646_, _16644_);
  nor _68111_ (_16649_, _08480_, _08651_);
  or _68112_ (_16650_, _16649_, _16647_);
  and _68113_ (_16651_, _16650_, _03759_);
  nor _68114_ (_16652_, _13035_, _07918_);
  nor _68115_ (_16653_, _16652_, _16397_);
  nor _68116_ (_16654_, _16653_, _03759_);
  or _68117_ (_16655_, _16654_, _08490_);
  or _68118_ (_16656_, _16655_, _16651_);
  and _68119_ (_16657_, _16656_, _16393_);
  or _68120_ (_16658_, _16657_, _07825_);
  and _68121_ (_16660_, _08512_, _08063_);
  nor _68122_ (_16661_, _16660_, _08513_);
  or _68123_ (_16662_, _16661_, _08495_);
  and _68124_ (_16663_, _16662_, _03766_);
  and _68125_ (_16664_, _16663_, _16658_);
  and _68126_ (_16665_, _08544_, _08247_);
  nor _68127_ (_16666_, _16665_, _08545_);
  and _68128_ (_16667_, _16666_, _03765_);
  or _68129_ (_16668_, _16667_, _08523_);
  or _68130_ (_16669_, _16668_, _16664_);
  and _68131_ (_16671_, _08574_, _08312_);
  nor _68132_ (_16672_, _16671_, _08575_);
  or _68133_ (_16673_, _16672_, _08557_);
  and _68134_ (_16674_, _16673_, _08556_);
  and _68135_ (_16675_, _16674_, _16669_);
  nand _68136_ (_16676_, _08555_, \oc8051_golden_model_1.ACC [4]);
  nand _68137_ (_16677_, _16676_, _07779_);
  or _68138_ (_16678_, _16677_, _16675_);
  and _68139_ (_16679_, _16428_, _07814_);
  nor _68140_ (_16680_, _16428_, _07814_);
  nor _68141_ (_16682_, _16680_, _16679_);
  or _68142_ (_16683_, _16682_, _07779_);
  and _68143_ (_16684_, _16683_, _07775_);
  and _68144_ (_16685_, _16684_, _16678_);
  and _68145_ (_16686_, _16682_, _07774_);
  or _68146_ (_16687_, _16686_, _07731_);
  or _68147_ (_16688_, _16687_, _16685_);
  and _68148_ (_16689_, _07765_, _07742_);
  nor _68149_ (_16690_, _16689_, _07766_);
  or _68150_ (_16691_, _16690_, _07732_);
  and _68151_ (_16693_, _16691_, _03526_);
  and _68152_ (_16694_, _16693_, _16688_);
  and _68153_ (_16695_, _08635_, _08610_);
  nor _68154_ (_16696_, _16695_, _08636_);
  and _68155_ (_16697_, _16696_, _03524_);
  or _68156_ (_16698_, _16697_, _08597_);
  or _68157_ (_16699_, _16698_, _16694_);
  and _68158_ (_16700_, _08674_, _08653_);
  nor _68159_ (_16701_, _16700_, _08675_);
  or _68160_ (_16702_, _16701_, _08598_);
  and _68161_ (_16704_, _16702_, _10803_);
  and _68162_ (_16705_, _16704_, _16699_);
  and _68163_ (_16706_, _07729_, \oc8051_golden_model_1.ACC [4]);
  or _68164_ (_16707_, _16706_, _03790_);
  or _68165_ (_16708_, _16707_, _16705_);
  nand _68166_ (_16709_, _16464_, _03790_);
  and _68167_ (_16710_, _16709_, _08688_);
  and _68168_ (_16711_, _16710_, _16708_);
  nor _68169_ (_16712_, _16360_, _07399_);
  or _68170_ (_16713_, _16712_, _08695_);
  and _68171_ (_16715_, _16713_, _08687_);
  or _68172_ (_16716_, _16715_, _08692_);
  or _68173_ (_16717_, _16716_, _16711_);
  nand _68174_ (_16718_, _08692_, _07346_);
  and _68175_ (_16719_, _16718_, _03152_);
  and _68176_ (_16720_, _16719_, _16717_);
  nor _68177_ (_16721_, _16495_, _03152_);
  or _68178_ (_16722_, _16721_, _03520_);
  or _68179_ (_16723_, _16722_, _16720_);
  and _68180_ (_16724_, _13097_, _05227_);
  nor _68181_ (_16726_, _16724_, _16397_);
  nand _68182_ (_16727_, _16726_, _03520_);
  and _68183_ (_16728_, _16727_, _08710_);
  and _68184_ (_16729_, _16728_, _16723_);
  nor _68185_ (_16730_, _08719_, \oc8051_golden_model_1.ACC [5]);
  nor _68186_ (_16731_, _16730_, _08720_);
  and _68187_ (_16732_, _16731_, _08709_);
  or _68188_ (_16733_, _16732_, _08716_);
  or _68189_ (_16734_, _16733_, _16729_);
  nand _68190_ (_16735_, _08716_, _07346_);
  and _68191_ (_16737_, _16735_, _42963_);
  and _68192_ (_16738_, _16737_, _16734_);
  or _68193_ (_16739_, _16738_, _16390_);
  and _68194_ (_43208_, _16739_, _41755_);
  nor _68195_ (_16740_, _42963_, _07346_);
  nand _68196_ (_16741_, _07729_, _07399_);
  nor _68197_ (_16742_, _07767_, _07738_);
  nor _68198_ (_16743_, _16742_, _07768_);
  or _68199_ (_16744_, _16743_, _07732_);
  nand _68200_ (_16745_, _08477_, _08647_);
  nand _68201_ (_16747_, _08458_, _07786_);
  nor _68202_ (_16748_, _05227_, _07346_);
  and _68203_ (_16749_, _13253_, _05227_);
  nor _68204_ (_16750_, _16749_, _16748_);
  nand _68205_ (_16751_, _16750_, _03636_);
  or _68206_ (_16752_, _08406_, _07738_);
  or _68207_ (_16753_, _07787_, _16404_);
  nand _68208_ (_16754_, _03561_, _03231_);
  nor _68209_ (_16755_, _05327_, _07918_);
  nor _68210_ (_16756_, _16755_, _16748_);
  nand _68211_ (_16758_, _16756_, _07314_);
  or _68212_ (_16759_, _16527_, _08608_);
  and _68213_ (_16760_, _16759_, _11479_);
  nor _68214_ (_16761_, _16760_, _08606_);
  and _68215_ (_16762_, _16760_, _08606_);
  nor _68216_ (_16763_, _16762_, _16761_);
  not _68217_ (_16764_, _16532_);
  nor _68218_ (_16765_, _16764_, _16763_);
  and _68219_ (_16766_, _16764_, _16763_);
  nor _68220_ (_16767_, _16766_, _16765_);
  nand _68221_ (_16769_, _16767_, _03614_);
  and _68222_ (_16770_, _16769_, _08109_);
  or _68223_ (_16771_, _06721_, _07399_);
  and _68224_ (_16772_, _06721_, _07399_);
  or _68225_ (_16773_, _16510_, _16772_);
  and _68226_ (_16774_, _16773_, _16771_);
  nor _68227_ (_16775_, _16774_, _07738_);
  and _68228_ (_16776_, _16774_, _07738_);
  nor _68229_ (_16777_, _16776_, _16775_);
  nor _68230_ (_16778_, _16520_, _16514_);
  and _68231_ (_16780_, _16778_, \oc8051_golden_model_1.PSW [7]);
  or _68232_ (_16781_, _16780_, _16777_);
  nand _68233_ (_16782_, _16780_, _16777_);
  and _68234_ (_16783_, _16782_, _16781_);
  and _68235_ (_16784_, _16783_, _08035_);
  nand _68236_ (_16785_, _07928_, _05327_);
  nand _68237_ (_16786_, _07933_, _05327_);
  nor _68238_ (_16787_, _04012_, _07346_);
  and _68239_ (_16788_, _04012_, _07346_);
  or _68240_ (_16789_, _16788_, _16787_);
  or _68241_ (_16791_, _16789_, _07933_);
  and _68242_ (_16792_, _16791_, _07936_);
  and _68243_ (_16793_, _16792_, _16786_);
  and _68244_ (_16794_, _07935_, _06713_);
  or _68245_ (_16795_, _16794_, _16793_);
  and _68246_ (_16796_, _16795_, _07946_);
  nor _68247_ (_16797_, _13122_, _07918_);
  nor _68248_ (_16798_, _16797_, _16748_);
  nor _68249_ (_16799_, _16798_, _04444_);
  or _68250_ (_16800_, _16799_, _07948_);
  or _68251_ (_16802_, _16800_, _16796_);
  not _68252_ (_16803_, _07965_);
  nor _68253_ (_16804_, _16469_, _16803_);
  and _68254_ (_16805_, _11548_, _07966_);
  nor _68255_ (_16806_, _16805_, _16804_);
  nand _68256_ (_16807_, _16806_, _07948_);
  and _68257_ (_16808_, _16807_, _03576_);
  and _68258_ (_16809_, _16808_, _16802_);
  nor _68259_ (_16810_, _05792_, _07346_);
  and _68260_ (_16811_, _13145_, _05792_);
  nor _68261_ (_16813_, _16811_, _16810_);
  nor _68262_ (_16814_, _16813_, _03517_);
  nor _68263_ (_16815_, _16756_, _03983_);
  or _68264_ (_16816_, _16815_, _07928_);
  or _68265_ (_16817_, _16816_, _16814_);
  or _68266_ (_16818_, _16817_, _16809_);
  and _68267_ (_16819_, _16818_, _16785_);
  or _68268_ (_16820_, _16819_, _04458_);
  or _68269_ (_16821_, _06713_, _07987_);
  and _68270_ (_16822_, _16821_, _03583_);
  and _68271_ (_16824_, _16822_, _16820_);
  nor _68272_ (_16825_, _08125_, _03583_);
  or _68273_ (_16826_, _16825_, _07991_);
  or _68274_ (_16827_, _16826_, _16824_);
  nand _68275_ (_16828_, _07991_, _07506_);
  and _68276_ (_16829_, _16828_, _16827_);
  or _68277_ (_16830_, _16829_, _03512_);
  and _68278_ (_16831_, _13130_, _05792_);
  nor _68279_ (_16832_, _16831_, _16810_);
  nand _68280_ (_16833_, _16832_, _03512_);
  and _68281_ (_16835_, _16833_, _03506_);
  and _68282_ (_16836_, _16835_, _16830_);
  and _68283_ (_16837_, _16811_, _13160_);
  nor _68284_ (_16838_, _16837_, _16810_);
  nor _68285_ (_16839_, _16838_, _03506_);
  or _68286_ (_16840_, _16839_, _06794_);
  or _68287_ (_16841_, _16840_, _16836_);
  nor _68288_ (_16842_, _07281_, _07279_);
  nor _68289_ (_16843_, _16842_, _07282_);
  or _68290_ (_16844_, _16843_, _06800_);
  and _68291_ (_16846_, _16844_, _16841_);
  or _68292_ (_16847_, _16846_, _07923_);
  nand _68293_ (_16848_, _05422_, \oc8051_golden_model_1.ACC [5]);
  nor _68294_ (_16849_, _05422_, \oc8051_golden_model_1.ACC [5]);
  or _68295_ (_16850_, _16430_, _16849_);
  and _68296_ (_16851_, _16850_, _16848_);
  nor _68297_ (_16852_, _16851_, _07787_);
  and _68298_ (_16853_, _16851_, _07787_);
  nor _68299_ (_16854_, _16853_, _16852_);
  nor _68300_ (_16855_, _16440_, _16434_);
  and _68301_ (_16857_, _16855_, \oc8051_golden_model_1.PSW [7]);
  or _68302_ (_16858_, _16857_, _16854_);
  nand _68303_ (_16859_, _16857_, _16854_);
  and _68304_ (_16860_, _16859_, _16858_);
  or _68305_ (_16861_, _16860_, _07922_);
  and _68306_ (_16862_, _16861_, _08037_);
  and _68307_ (_16863_, _16862_, _16847_);
  or _68308_ (_16864_, _16863_, _03614_);
  or _68309_ (_16865_, _16864_, _16784_);
  and _68310_ (_16866_, _16865_, _16770_);
  or _68311_ (_16868_, _16413_, _11504_);
  and _68312_ (_16869_, _16868_, _11503_);
  nor _68313_ (_16870_, _16869_, _08649_);
  and _68314_ (_16871_, _16869_, _08649_);
  nor _68315_ (_16872_, _16871_, _16870_);
  nor _68316_ (_16873_, _16423_, _16418_);
  and _68317_ (_16874_, _16873_, \oc8051_golden_model_1.PSW [7]);
  nor _68318_ (_16875_, _16874_, _16872_);
  and _68319_ (_16876_, _16874_, _16872_);
  nor _68320_ (_16877_, _16876_, _16875_);
  and _68321_ (_16879_, _16877_, _08108_);
  or _68322_ (_16880_, _16879_, _03311_);
  or _68323_ (_16881_, _16880_, _16866_);
  nand _68324_ (_16882_, _03561_, _03311_);
  and _68325_ (_16883_, _16882_, _03500_);
  and _68326_ (_16884_, _16883_, _16881_);
  nor _68327_ (_16885_, _13178_, _08358_);
  nor _68328_ (_16886_, _16885_, _16810_);
  nor _68329_ (_16887_, _16886_, _03500_);
  or _68330_ (_16888_, _16887_, _07314_);
  or _68331_ (_16890_, _16888_, _16884_);
  and _68332_ (_16891_, _16890_, _16758_);
  or _68333_ (_16892_, _16891_, _03479_);
  and _68334_ (_16893_, _06713_, _05227_);
  nor _68335_ (_16894_, _16893_, _16748_);
  nand _68336_ (_16895_, _16894_, _03479_);
  and _68337_ (_16896_, _16895_, _03474_);
  and _68338_ (_16897_, _16896_, _16892_);
  nor _68339_ (_16898_, _13237_, _07918_);
  nor _68340_ (_16899_, _16898_, _16748_);
  nor _68341_ (_16901_, _16899_, _03474_);
  or _68342_ (_16902_, _16901_, _07328_);
  or _68343_ (_16903_, _16902_, _16897_);
  not _68344_ (_16904_, _07347_);
  and _68345_ (_16905_, _07352_, _16904_);
  or _68346_ (_16906_, _16905_, _07677_);
  and _68347_ (_16907_, _16906_, _16903_);
  or _68348_ (_16908_, _16907_, _03231_);
  and _68349_ (_16909_, _16908_, _16754_);
  or _68350_ (_16910_, _16909_, _03437_);
  and _68351_ (_16912_, _13244_, _05227_);
  nor _68352_ (_16913_, _16912_, _16748_);
  nand _68353_ (_16914_, _16913_, _03437_);
  and _68354_ (_16915_, _16914_, _08386_);
  and _68355_ (_16916_, _16915_, _16910_);
  nor _68356_ (_16917_, _08386_, _03561_);
  or _68357_ (_16918_, _16917_, _16403_);
  or _68358_ (_16919_, _16918_, _16916_);
  and _68359_ (_16920_, _16919_, _16753_);
  or _68360_ (_16921_, _16920_, _16402_);
  not _68361_ (_16923_, _07787_);
  and _68362_ (_16924_, _16923_, _16402_);
  nor _68363_ (_16925_, _16924_, _03935_);
  and _68364_ (_16926_, _16925_, _16921_);
  nor _68365_ (_16927_, _07787_, _03043_);
  nor _68366_ (_16928_, _16927_, _16581_);
  or _68367_ (_16929_, _16928_, _16926_);
  or _68368_ (_16930_, _07787_, _03933_);
  and _68369_ (_16931_, _16930_, _16929_);
  or _68370_ (_16932_, _16931_, _04325_);
  nand _68371_ (_16934_, _16923_, _04325_);
  and _68372_ (_16935_, _16934_, _16254_);
  and _68373_ (_16936_, _16935_, _16932_);
  and _68374_ (_16937_, _16253_, _07787_);
  or _68375_ (_16938_, _16937_, _08405_);
  or _68376_ (_16939_, _16938_, _16936_);
  and _68377_ (_16940_, _16939_, _16752_);
  or _68378_ (_16941_, _16940_, _03767_);
  or _68379_ (_16942_, _13259_, _03768_);
  and _68380_ (_16943_, _16942_, _08416_);
  and _68381_ (_16945_, _16943_, _16941_);
  nor _68382_ (_16946_, _08416_, _08648_);
  or _68383_ (_16947_, _16946_, _03636_);
  or _68384_ (_16948_, _16947_, _16945_);
  and _68385_ (_16949_, _16948_, _16751_);
  or _68386_ (_16950_, _16949_, _03769_);
  or _68387_ (_16951_, _16748_, _04501_);
  and _68388_ (_16952_, _16951_, _08435_);
  and _68389_ (_16953_, _16952_, _16950_);
  and _68390_ (_16954_, _08436_, _07785_);
  or _68391_ (_16956_, _16954_, _04135_);
  or _68392_ (_16957_, _16956_, _16953_);
  or _68393_ (_16958_, _07785_, _08440_);
  and _68394_ (_16959_, _16958_, _08446_);
  and _68395_ (_16960_, _16959_, _16957_);
  and _68396_ (_16961_, _08445_, _07736_);
  or _68397_ (_16962_, _16961_, _03755_);
  or _68398_ (_16963_, _16962_, _16960_);
  or _68399_ (_16964_, _13257_, _07911_);
  and _68400_ (_16965_, _16964_, _07910_);
  and _68401_ (_16967_, _16965_, _16963_);
  and _68402_ (_16968_, _08646_, _07909_);
  or _68403_ (_16969_, _16968_, _16967_);
  and _68404_ (_16970_, _16969_, _05769_);
  or _68405_ (_16971_, _16913_, _13258_);
  nor _68406_ (_16972_, _16971_, _04505_);
  or _68407_ (_16973_, _16972_, _08458_);
  or _68408_ (_16974_, _16973_, _16970_);
  and _68409_ (_16975_, _16974_, _16747_);
  or _68410_ (_16976_, _16975_, _08465_);
  nor _68411_ (_16978_, _07786_, _04161_);
  or _68412_ (_16979_, _16978_, _08466_);
  and _68413_ (_16980_, _16979_, _16976_);
  nor _68414_ (_16981_, _07786_, _15029_);
  or _68415_ (_16982_, _16981_, _08469_);
  or _68416_ (_16983_, _16982_, _16980_);
  nand _68417_ (_16984_, _08469_, _07737_);
  and _68418_ (_16985_, _16984_, _08473_);
  and _68419_ (_16986_, _16985_, _16983_);
  nand _68420_ (_16987_, _13258_, _08480_);
  and _68421_ (_16989_, _16987_, _08479_);
  or _68422_ (_16990_, _16989_, _16986_);
  and _68423_ (_16991_, _16990_, _16745_);
  or _68424_ (_16992_, _16991_, _03758_);
  nor _68425_ (_16993_, _13251_, _07918_);
  nor _68426_ (_16994_, _16993_, _16748_);
  nand _68427_ (_16995_, _16994_, _03758_);
  and _68428_ (_16996_, _16995_, _07830_);
  and _68429_ (_16997_, _16996_, _16992_);
  nor _68430_ (_16998_, _07902_, _07846_);
  nor _68431_ (_17000_, _16998_, _07903_);
  or _68432_ (_17001_, _17000_, _07825_);
  and _68433_ (_17002_, _17001_, _10581_);
  or _68434_ (_17003_, _17002_, _16997_);
  nor _68435_ (_17004_, _08514_, _08099_);
  nor _68436_ (_17005_, _17004_, _08515_);
  or _68437_ (_17006_, _17005_, _08495_);
  and _68438_ (_17007_, _17006_, _03766_);
  and _68439_ (_17008_, _17007_, _17003_);
  nor _68440_ (_17009_, _08546_, _08527_);
  nor _68441_ (_17011_, _17009_, _08547_);
  or _68442_ (_17012_, _17011_, _08523_);
  and _68443_ (_17013_, _17012_, _08525_);
  or _68444_ (_17014_, _17013_, _17008_);
  nor _68445_ (_17015_, _08576_, _08346_);
  nor _68446_ (_17016_, _17015_, _08577_);
  or _68447_ (_17017_, _17016_, _08557_);
  and _68448_ (_17018_, _17017_, _17014_);
  or _68449_ (_17019_, _17018_, _08555_);
  nand _68450_ (_17020_, _08555_, _07399_);
  and _68451_ (_17022_, _17020_, _07780_);
  and _68452_ (_17023_, _17022_, _17019_);
  nor _68453_ (_17024_, _07816_, _07787_);
  nor _68454_ (_17025_, _17024_, _07817_);
  or _68455_ (_17026_, _17025_, _07731_);
  and _68456_ (_17027_, _17026_, _10603_);
  or _68457_ (_17028_, _17027_, _17023_);
  and _68458_ (_17029_, _17028_, _16744_);
  or _68459_ (_17030_, _17029_, _03524_);
  nor _68460_ (_17031_, _08637_, _08606_);
  nor _68461_ (_17033_, _17031_, _08638_);
  or _68462_ (_17034_, _17033_, _03526_);
  and _68463_ (_17035_, _17034_, _08598_);
  and _68464_ (_17036_, _17035_, _17030_);
  nor _68465_ (_17037_, _08676_, _08649_);
  nor _68466_ (_17038_, _17037_, _08677_);
  and _68467_ (_17039_, _17038_, _08597_);
  or _68468_ (_17040_, _17039_, _07729_);
  or _68469_ (_17041_, _17040_, _17036_);
  and _68470_ (_17042_, _17041_, _16741_);
  or _68471_ (_17044_, _17042_, _03790_);
  nand _68472_ (_17045_, _16798_, _03790_);
  and _68473_ (_17046_, _17045_, _08688_);
  and _68474_ (_17047_, _17046_, _17044_);
  nor _68475_ (_17048_, _08695_, _07346_);
  or _68476_ (_17049_, _17048_, _08696_);
  nor _68477_ (_17050_, _17049_, _08692_);
  nor _68478_ (_17051_, _17050_, _10828_);
  or _68479_ (_17052_, _17051_, _17047_);
  nand _68480_ (_17053_, _08692_, _05834_);
  and _68481_ (_17055_, _17053_, _03152_);
  and _68482_ (_17056_, _17055_, _17052_);
  nor _68483_ (_17057_, _16832_, _03152_);
  or _68484_ (_17058_, _17057_, _03520_);
  or _68485_ (_17059_, _17058_, _17056_);
  and _68486_ (_17060_, _13312_, _05227_);
  nor _68487_ (_17061_, _17060_, _16748_);
  nand _68488_ (_17062_, _17061_, _03520_);
  and _68489_ (_17063_, _17062_, _08710_);
  and _68490_ (_17064_, _17063_, _17059_);
  nor _68491_ (_17066_, _08720_, \oc8051_golden_model_1.ACC [6]);
  nor _68492_ (_17067_, _17066_, _08721_);
  and _68493_ (_17068_, _17067_, _08709_);
  or _68494_ (_17069_, _17068_, _08716_);
  or _68495_ (_17070_, _17069_, _17064_);
  nand _68496_ (_17071_, _08716_, _05834_);
  and _68497_ (_17072_, _17071_, _42963_);
  and _68498_ (_17073_, _17072_, _17070_);
  or _68499_ (_17074_, _17073_, _16740_);
  and _68500_ (_43209_, _17074_, _41755_);
  not _68501_ (_17076_, _03882_);
  not _68502_ (_17077_, \oc8051_golden_model_1.SBUF [0]);
  nor _68503_ (_17078_, _05185_, _17077_);
  and _68504_ (_17079_, _05941_, _05185_);
  nor _68505_ (_17080_, _17079_, _17078_);
  and _68506_ (_17081_, _17080_, _17076_);
  and _68507_ (_17082_, _05185_, \oc8051_golden_model_1.ACC [0]);
  nor _68508_ (_17083_, _17082_, _17078_);
  nor _68509_ (_17084_, _17083_, _03583_);
  nor _68510_ (_17085_, _17083_, _04427_);
  nor _68511_ (_17087_, _04426_, _17077_);
  or _68512_ (_17088_, _17087_, _17085_);
  and _68513_ (_17089_, _17088_, _04444_);
  nor _68514_ (_17090_, _17080_, _04444_);
  or _68515_ (_17091_, _17090_, _17089_);
  and _68516_ (_17092_, _17091_, _03983_);
  and _68517_ (_17093_, _05185_, _04419_);
  nor _68518_ (_17094_, _17093_, _17078_);
  nor _68519_ (_17095_, _17094_, _03983_);
  nor _68520_ (_17096_, _17095_, _17092_);
  nor _68521_ (_17098_, _17096_, _03575_);
  or _68522_ (_17099_, _17098_, _07314_);
  nor _68523_ (_17100_, _17099_, _17084_);
  and _68524_ (_17101_, _17094_, _07314_);
  nor _68525_ (_17102_, _17101_, _17100_);
  nor _68526_ (_17103_, _17102_, _03479_);
  and _68527_ (_17104_, _06715_, _05185_);
  nor _68528_ (_17105_, _17078_, _06044_);
  not _68529_ (_17106_, _17105_);
  nor _68530_ (_17107_, _17106_, _17104_);
  nor _68531_ (_17109_, _17107_, _17103_);
  nor _68532_ (_17110_, _17109_, _03221_);
  nor _68533_ (_17111_, _11975_, _08737_);
  or _68534_ (_17112_, _17078_, _03474_);
  nor _68535_ (_17113_, _17112_, _17111_);
  or _68536_ (_17114_, _17113_, _03437_);
  nor _68537_ (_17115_, _17114_, _17110_);
  and _68538_ (_17116_, _05185_, _06202_);
  nor _68539_ (_17117_, _17116_, _17078_);
  nor _68540_ (_17118_, _17117_, _03438_);
  or _68541_ (_17120_, _17118_, _17115_);
  and _68542_ (_17121_, _17120_, _04499_);
  and _68543_ (_17122_, _11990_, _05185_);
  nor _68544_ (_17123_, _17122_, _17078_);
  nor _68545_ (_17124_, _17123_, _04499_);
  or _68546_ (_17125_, _17124_, _17121_);
  nor _68547_ (_17126_, _17125_, _03769_);
  and _68548_ (_17127_, _11995_, _05185_);
  or _68549_ (_17128_, _17078_, _04501_);
  nor _68550_ (_17129_, _17128_, _17127_);
  or _68551_ (_17131_, _17129_, _04504_);
  nor _68552_ (_17132_, _17131_, _17126_);
  or _68553_ (_17133_, _17117_, _04505_);
  nor _68554_ (_17134_, _17133_, _17079_);
  nor _68555_ (_17135_, _17134_, _17132_);
  nor _68556_ (_17136_, _17135_, _03752_);
  nor _68557_ (_17137_, _17078_, _05617_);
  or _68558_ (_17138_, _17137_, _03753_);
  nor _68559_ (_17139_, _17138_, _17083_);
  or _68560_ (_17140_, _17139_, _17136_);
  and _68561_ (_17142_, _17140_, _03759_);
  nor _68562_ (_17143_, _11988_, _08737_);
  nor _68563_ (_17144_, _17143_, _17078_);
  nor _68564_ (_17145_, _17144_, _03759_);
  or _68565_ (_17146_, _17145_, _17142_);
  and _68566_ (_17147_, _17146_, _04517_);
  nor _68567_ (_17148_, _11870_, _08737_);
  nor _68568_ (_17149_, _17148_, _17078_);
  nor _68569_ (_17150_, _17149_, _04517_);
  nor _68570_ (_17151_, _17150_, _17076_);
  not _68571_ (_17153_, _17151_);
  nor _68572_ (_17154_, _17153_, _17147_);
  nor _68573_ (_17155_, _17154_, _17081_);
  or _68574_ (_17156_, _17155_, _42967_);
  or _68575_ (_17157_, _42963_, \oc8051_golden_model_1.SBUF [0]);
  and _68576_ (_17158_, _17157_, _41755_);
  and _68577_ (_43210_, _17158_, _17156_);
  nor _68578_ (_17159_, _05185_, \oc8051_golden_model_1.SBUF [1]);
  and _68579_ (_17160_, _12252_, _05185_);
  nor _68580_ (_17161_, _17160_, _17159_);
  nor _68581_ (_17163_, _17161_, _04192_);
  and _68582_ (_17164_, _06714_, _05185_);
  not _68583_ (_17165_, \oc8051_golden_model_1.SBUF [1]);
  nor _68584_ (_17166_, _05185_, _17165_);
  nor _68585_ (_17167_, _17166_, _06044_);
  not _68586_ (_17168_, _17167_);
  nor _68587_ (_17169_, _17168_, _17164_);
  not _68588_ (_17170_, _17169_);
  and _68589_ (_17171_, _05185_, _03233_);
  nor _68590_ (_17172_, _17171_, _17159_);
  and _68591_ (_17174_, _17172_, _03575_);
  nor _68592_ (_17175_, _08737_, _04603_);
  nor _68593_ (_17176_, _17175_, _17166_);
  nor _68594_ (_17177_, _17176_, _03983_);
  and _68595_ (_17178_, _17172_, _04426_);
  nor _68596_ (_17179_, _04426_, _17165_);
  or _68597_ (_17180_, _17179_, _17178_);
  and _68598_ (_17181_, _17180_, _04444_);
  and _68599_ (_17182_, _17161_, _03570_);
  or _68600_ (_17183_, _17182_, _17181_);
  and _68601_ (_17185_, _17183_, _03983_);
  nor _68602_ (_17186_, _17185_, _17177_);
  nor _68603_ (_17187_, _17186_, _03575_);
  or _68604_ (_17188_, _17187_, _07314_);
  nor _68605_ (_17189_, _17188_, _17174_);
  and _68606_ (_17190_, _17176_, _07314_);
  nor _68607_ (_17191_, _17190_, _17189_);
  nor _68608_ (_17192_, _17191_, _03479_);
  nor _68609_ (_17193_, _17192_, _03221_);
  and _68610_ (_17194_, _17193_, _17170_);
  not _68611_ (_17196_, _17159_);
  and _68612_ (_17197_, _12176_, _05185_);
  nor _68613_ (_17198_, _17197_, _03474_);
  and _68614_ (_17199_, _17198_, _17196_);
  nor _68615_ (_17200_, _17199_, _17194_);
  nor _68616_ (_17201_, _17200_, _03437_);
  and _68617_ (_17202_, _05185_, _04317_);
  not _68618_ (_17203_, _17202_);
  nor _68619_ (_17204_, _17159_, _03438_);
  and _68620_ (_17205_, _17204_, _17203_);
  nor _68621_ (_17207_, _17205_, _17201_);
  nor _68622_ (_17208_, _17207_, _03636_);
  nor _68623_ (_17209_, _12191_, _08737_);
  nor _68624_ (_17210_, _17209_, _04499_);
  and _68625_ (_17211_, _17210_, _17196_);
  nor _68626_ (_17212_, _17211_, _17208_);
  nor _68627_ (_17213_, _17212_, _03769_);
  nor _68628_ (_17214_, _12197_, _08737_);
  nor _68629_ (_17215_, _17214_, _04501_);
  and _68630_ (_17216_, _17215_, _17196_);
  nor _68631_ (_17218_, _17216_, _17213_);
  nor _68632_ (_17219_, _17218_, _04504_);
  nor _68633_ (_17220_, _12190_, _08737_);
  nor _68634_ (_17221_, _17220_, _05769_);
  and _68635_ (_17222_, _17221_, _17196_);
  nor _68636_ (_17223_, _17222_, _17219_);
  nor _68637_ (_17224_, _17223_, _03752_);
  nor _68638_ (_17225_, _17166_, _05569_);
  nor _68639_ (_17226_, _17225_, _03753_);
  and _68640_ (_17227_, _17226_, _17172_);
  nor _68641_ (_17229_, _17227_, _17224_);
  nor _68642_ (_17230_, _17229_, _03758_);
  and _68643_ (_17231_, _17202_, _05940_);
  nor _68644_ (_17232_, _17231_, _03759_);
  and _68645_ (_17233_, _17232_, _17196_);
  nor _68646_ (_17234_, _17233_, _17230_);
  nor _68647_ (_17235_, _17234_, _03760_);
  nand _68648_ (_17236_, _17171_, _05940_);
  nor _68649_ (_17237_, _17159_, _04517_);
  and _68650_ (_17238_, _17237_, _17236_);
  or _68651_ (_17240_, _17238_, _03790_);
  nor _68652_ (_17241_, _17240_, _17235_);
  nor _68653_ (_17242_, _17241_, _17163_);
  and _68654_ (_17243_, _17242_, _03521_);
  nor _68655_ (_17244_, _17166_, _17160_);
  nor _68656_ (_17245_, _17244_, _03521_);
  or _68657_ (_17246_, _17245_, _17243_);
  or _68658_ (_17247_, _17246_, _42967_);
  or _68659_ (_17248_, _42963_, \oc8051_golden_model_1.SBUF [1]);
  and _68660_ (_17249_, _17248_, _41755_);
  and _68661_ (_43211_, _17249_, _17247_);
  not _68662_ (_17251_, \oc8051_golden_model_1.SBUF [2]);
  nor _68663_ (_17252_, _05185_, _17251_);
  nor _68664_ (_17253_, _12400_, _08737_);
  nor _68665_ (_17254_, _17253_, _17252_);
  nor _68666_ (_17255_, _17254_, _04517_);
  nor _68667_ (_17256_, _08737_, _05026_);
  nor _68668_ (_17257_, _17256_, _17252_);
  and _68669_ (_17258_, _17257_, _07314_);
  and _68670_ (_17259_, _05185_, \oc8051_golden_model_1.ACC [2]);
  nor _68671_ (_17261_, _17259_, _17252_);
  nor _68672_ (_17262_, _17261_, _04427_);
  nor _68673_ (_17263_, _04426_, _17251_);
  or _68674_ (_17264_, _17263_, _17262_);
  and _68675_ (_17265_, _17264_, _04444_);
  nor _68676_ (_17266_, _12282_, _08737_);
  nor _68677_ (_17267_, _17266_, _17252_);
  nor _68678_ (_17268_, _17267_, _04444_);
  or _68679_ (_17269_, _17268_, _17265_);
  and _68680_ (_17270_, _17269_, _03983_);
  nor _68681_ (_17272_, _17257_, _03983_);
  nor _68682_ (_17273_, _17272_, _17270_);
  nor _68683_ (_17274_, _17273_, _03575_);
  nor _68684_ (_17275_, _17261_, _03583_);
  nor _68685_ (_17276_, _17275_, _07314_);
  not _68686_ (_17277_, _17276_);
  nor _68687_ (_17278_, _17277_, _17274_);
  nor _68688_ (_17279_, _17278_, _17258_);
  nor _68689_ (_17280_, _17279_, _03479_);
  and _68690_ (_17281_, _06718_, _05185_);
  nor _68691_ (_17282_, _17252_, _06044_);
  not _68692_ (_17283_, _17282_);
  nor _68693_ (_17284_, _17283_, _17281_);
  nor _68694_ (_17285_, _17284_, _17280_);
  nor _68695_ (_17286_, _17285_, _03221_);
  nor _68696_ (_17287_, _12384_, _08737_);
  or _68697_ (_17288_, _17252_, _03474_);
  nor _68698_ (_17289_, _17288_, _17287_);
  or _68699_ (_17290_, _17289_, _03437_);
  nor _68700_ (_17291_, _17290_, _17286_);
  and _68701_ (_17294_, _05185_, _06261_);
  nor _68702_ (_17295_, _17294_, _17252_);
  nor _68703_ (_17296_, _17295_, _03438_);
  or _68704_ (_17297_, _17296_, _17291_);
  and _68705_ (_17298_, _17297_, _04499_);
  and _68706_ (_17299_, _12273_, _05185_);
  nor _68707_ (_17300_, _17299_, _17252_);
  nor _68708_ (_17301_, _17300_, _04499_);
  or _68709_ (_17302_, _17301_, _17298_);
  nor _68710_ (_17303_, _17302_, _03769_);
  and _68711_ (_17304_, _12401_, _05185_);
  or _68712_ (_17305_, _17252_, _04501_);
  nor _68713_ (_17306_, _17305_, _17304_);
  or _68714_ (_17307_, _17306_, _04504_);
  nor _68715_ (_17308_, _17307_, _17303_);
  nor _68716_ (_17309_, _17252_, _05665_);
  or _68717_ (_17310_, _17295_, _04505_);
  nor _68718_ (_17311_, _17310_, _17309_);
  nor _68719_ (_17312_, _17311_, _17308_);
  nor _68720_ (_17313_, _17312_, _03752_);
  or _68721_ (_17316_, _17309_, _03753_);
  or _68722_ (_17317_, _17316_, _17261_);
  and _68723_ (_17318_, _17317_, _03759_);
  not _68724_ (_17319_, _17318_);
  nor _68725_ (_17320_, _17319_, _17313_);
  nor _68726_ (_17321_, _12272_, _08737_);
  or _68727_ (_17322_, _17252_, _03759_);
  nor _68728_ (_17323_, _17322_, _17321_);
  or _68729_ (_17324_, _17323_, _03760_);
  nor _68730_ (_17325_, _17324_, _17320_);
  nor _68731_ (_17327_, _17325_, _17255_);
  nor _68732_ (_17328_, _17327_, _03790_);
  nor _68733_ (_17329_, _17267_, _04192_);
  or _68734_ (_17330_, _17329_, _03520_);
  nor _68735_ (_17331_, _17330_, _17328_);
  and _68736_ (_17332_, _12456_, _05185_);
  or _68737_ (_17333_, _17252_, _03521_);
  nor _68738_ (_17334_, _17333_, _17332_);
  nor _68739_ (_17335_, _17334_, _17331_);
  or _68740_ (_17336_, _17335_, _42967_);
  or _68741_ (_17338_, _42963_, \oc8051_golden_model_1.SBUF [2]);
  and _68742_ (_17339_, _17338_, _41755_);
  and _68743_ (_43212_, _17339_, _17336_);
  not _68744_ (_17340_, \oc8051_golden_model_1.SBUF [3]);
  nor _68745_ (_17341_, _05185_, _17340_);
  and _68746_ (_17342_, _06717_, _05185_);
  nor _68747_ (_17343_, _17342_, _17341_);
  or _68748_ (_17344_, _17343_, _06044_);
  and _68749_ (_17345_, _05185_, \oc8051_golden_model_1.ACC [3]);
  nor _68750_ (_17346_, _17345_, _17341_);
  nor _68751_ (_17348_, _17346_, _04427_);
  nor _68752_ (_17349_, _04426_, _17340_);
  or _68753_ (_17350_, _17349_, _17348_);
  and _68754_ (_17351_, _17350_, _04444_);
  nor _68755_ (_17352_, _12486_, _08737_);
  nor _68756_ (_17353_, _17352_, _17341_);
  nor _68757_ (_17354_, _17353_, _04444_);
  or _68758_ (_17355_, _17354_, _17351_);
  and _68759_ (_17356_, _17355_, _03983_);
  nor _68760_ (_17357_, _08737_, _04843_);
  nor _68761_ (_17359_, _17357_, _17341_);
  nor _68762_ (_17360_, _17359_, _03983_);
  nor _68763_ (_17361_, _17360_, _17356_);
  nor _68764_ (_17362_, _17361_, _03575_);
  nor _68765_ (_17363_, _17346_, _03583_);
  nor _68766_ (_17364_, _17363_, _07314_);
  not _68767_ (_17365_, _17364_);
  nor _68768_ (_17366_, _17365_, _17362_);
  and _68769_ (_17367_, _17359_, _07314_);
  or _68770_ (_17368_, _17367_, _03479_);
  or _68771_ (_17370_, _17368_, _17366_);
  and _68772_ (_17371_, _17370_, _03474_);
  and _68773_ (_17372_, _17371_, _17344_);
  nor _68774_ (_17373_, _12583_, _08737_);
  or _68775_ (_17374_, _17341_, _03474_);
  nor _68776_ (_17375_, _17374_, _17373_);
  or _68777_ (_17376_, _17375_, _03437_);
  nor _68778_ (_17377_, _17376_, _17372_);
  and _68779_ (_17378_, _05185_, _06217_);
  nor _68780_ (_17379_, _17378_, _17341_);
  nor _68781_ (_17381_, _17379_, _03438_);
  or _68782_ (_17382_, _17381_, _17377_);
  and _68783_ (_17383_, _17382_, _04499_);
  and _68784_ (_17384_, _12598_, _05185_);
  nor _68785_ (_17385_, _17384_, _17341_);
  nor _68786_ (_17386_, _17385_, _04499_);
  or _68787_ (_17387_, _17386_, _17383_);
  nor _68788_ (_17388_, _17387_, _03769_);
  and _68789_ (_17389_, _12604_, _05185_);
  or _68790_ (_17390_, _17341_, _04501_);
  nor _68791_ (_17392_, _17390_, _17389_);
  or _68792_ (_17393_, _17392_, _04504_);
  nor _68793_ (_17394_, _17393_, _17388_);
  nor _68794_ (_17395_, _17341_, _05521_);
  or _68795_ (_17396_, _17379_, _04505_);
  nor _68796_ (_17397_, _17396_, _17395_);
  nor _68797_ (_17398_, _17397_, _17394_);
  nor _68798_ (_17399_, _17398_, _03752_);
  or _68799_ (_17400_, _17395_, _03753_);
  or _68800_ (_17401_, _17400_, _17346_);
  and _68801_ (_17403_, _17401_, _03759_);
  not _68802_ (_17404_, _17403_);
  nor _68803_ (_17405_, _17404_, _17399_);
  nor _68804_ (_17406_, _12597_, _08737_);
  or _68805_ (_17407_, _17341_, _03759_);
  nor _68806_ (_17408_, _17407_, _17406_);
  or _68807_ (_17409_, _17408_, _03760_);
  nor _68808_ (_17410_, _17409_, _17405_);
  nor _68809_ (_17411_, _12603_, _08737_);
  nor _68810_ (_17412_, _17411_, _17341_);
  nor _68811_ (_17414_, _17412_, _04517_);
  or _68812_ (_17415_, _17414_, _03790_);
  nor _68813_ (_17416_, _17415_, _17410_);
  and _68814_ (_17417_, _17353_, _03790_);
  or _68815_ (_17418_, _17417_, _03520_);
  nor _68816_ (_17419_, _17418_, _17416_);
  and _68817_ (_17420_, _12658_, _05185_);
  nor _68818_ (_17421_, _17420_, _17341_);
  nor _68819_ (_17422_, _17421_, _03521_);
  or _68820_ (_17423_, _17422_, _17419_);
  or _68821_ (_17425_, _17423_, _42967_);
  or _68822_ (_17426_, _42963_, \oc8051_golden_model_1.SBUF [3]);
  and _68823_ (_17427_, _17426_, _41755_);
  and _68824_ (_43213_, _17427_, _17425_);
  not _68825_ (_17428_, \oc8051_golden_model_1.SBUF [4]);
  nor _68826_ (_17429_, _05185_, _17428_);
  and _68827_ (_17430_, _12844_, _05185_);
  nor _68828_ (_17431_, _17430_, _17429_);
  nor _68829_ (_17432_, _17431_, _04501_);
  and _68830_ (_17433_, _05185_, \oc8051_golden_model_1.ACC [4]);
  nor _68831_ (_17435_, _17433_, _17429_);
  nor _68832_ (_17436_, _17435_, _04427_);
  nor _68833_ (_17437_, _04426_, _17428_);
  or _68834_ (_17438_, _17437_, _17436_);
  and _68835_ (_17439_, _17438_, _04444_);
  nor _68836_ (_17440_, _12733_, _08737_);
  nor _68837_ (_17441_, _17440_, _17429_);
  nor _68838_ (_17442_, _17441_, _04444_);
  or _68839_ (_17443_, _17442_, _17439_);
  and _68840_ (_17444_, _17443_, _03983_);
  nor _68841_ (_17446_, _05712_, _08737_);
  nor _68842_ (_17447_, _17446_, _17429_);
  nor _68843_ (_17448_, _17447_, _03983_);
  nor _68844_ (_17449_, _17448_, _17444_);
  nor _68845_ (_17450_, _17449_, _03575_);
  nor _68846_ (_17451_, _17435_, _03583_);
  nor _68847_ (_17452_, _17451_, _07314_);
  not _68848_ (_17453_, _17452_);
  nor _68849_ (_17454_, _17453_, _17450_);
  and _68850_ (_17455_, _17447_, _07314_);
  or _68851_ (_17457_, _17455_, _03479_);
  nor _68852_ (_17458_, _17457_, _17454_);
  and _68853_ (_17459_, _06722_, _05185_);
  or _68854_ (_17460_, _17459_, _17429_);
  and _68855_ (_17461_, _17460_, _03479_);
  or _68856_ (_17462_, _17461_, _03221_);
  or _68857_ (_17463_, _17462_, _17458_);
  nor _68858_ (_17464_, _12827_, _08737_);
  or _68859_ (_17465_, _17429_, _03474_);
  or _68860_ (_17466_, _17465_, _17464_);
  and _68861_ (_17468_, _17466_, _03438_);
  and _68862_ (_17469_, _17468_, _17463_);
  and _68863_ (_17470_, _06233_, _05185_);
  nor _68864_ (_17471_, _17470_, _17429_);
  nor _68865_ (_17472_, _17471_, _03438_);
  or _68866_ (_17473_, _17472_, _03636_);
  nor _68867_ (_17474_, _17473_, _17469_);
  and _68868_ (_17475_, _12711_, _05185_);
  or _68869_ (_17476_, _17429_, _04499_);
  nor _68870_ (_17477_, _17476_, _17475_);
  or _68871_ (_17479_, _17477_, _03769_);
  nor _68872_ (_17480_, _17479_, _17474_);
  nor _68873_ (_17481_, _17480_, _17432_);
  nor _68874_ (_17482_, _17481_, _04504_);
  not _68875_ (_17483_, _17429_);
  and _68876_ (_17484_, _17483_, _05760_);
  or _68877_ (_17485_, _17471_, _04505_);
  nor _68878_ (_17486_, _17485_, _17484_);
  nor _68879_ (_17487_, _17486_, _17482_);
  nor _68880_ (_17488_, _17487_, _03752_);
  or _68881_ (_17490_, _17484_, _03753_);
  or _68882_ (_17491_, _17490_, _17435_);
  and _68883_ (_17492_, _17491_, _03759_);
  not _68884_ (_17493_, _17492_);
  nor _68885_ (_17494_, _17493_, _17488_);
  nor _68886_ (_17495_, _12710_, _08737_);
  or _68887_ (_17496_, _17429_, _03759_);
  nor _68888_ (_17497_, _17496_, _17495_);
  or _68889_ (_17498_, _17497_, _03760_);
  nor _68890_ (_17499_, _17498_, _17494_);
  nor _68891_ (_17501_, _12843_, _08737_);
  nor _68892_ (_17502_, _17501_, _17429_);
  nor _68893_ (_17503_, _17502_, _04517_);
  or _68894_ (_17504_, _17503_, _03790_);
  nor _68895_ (_17505_, _17504_, _17499_);
  and _68896_ (_17506_, _17441_, _03790_);
  or _68897_ (_17507_, _17506_, _03520_);
  nor _68898_ (_17508_, _17507_, _17505_);
  and _68899_ (_17509_, _12893_, _05185_);
  nor _68900_ (_17510_, _17509_, _17429_);
  nor _68901_ (_17512_, _17510_, _03521_);
  or _68902_ (_17513_, _17512_, _17508_);
  or _68903_ (_17514_, _17513_, _42967_);
  or _68904_ (_17515_, _42963_, \oc8051_golden_model_1.SBUF [4]);
  and _68905_ (_17516_, _17515_, _41755_);
  and _68906_ (_43214_, _17516_, _17514_);
  not _68907_ (_17517_, \oc8051_golden_model_1.SBUF [5]);
  nor _68908_ (_17518_, _05185_, _17517_);
  and _68909_ (_17519_, _13042_, _05185_);
  nor _68910_ (_17520_, _17519_, _17518_);
  nor _68911_ (_17522_, _17520_, _04501_);
  nor _68912_ (_17523_, _05422_, _08737_);
  nor _68913_ (_17524_, _17523_, _17518_);
  and _68914_ (_17525_, _17524_, _07314_);
  and _68915_ (_17526_, _05185_, \oc8051_golden_model_1.ACC [5]);
  nor _68916_ (_17527_, _17526_, _17518_);
  nor _68917_ (_17528_, _17527_, _04427_);
  nor _68918_ (_17529_, _04426_, _17517_);
  or _68919_ (_17530_, _17529_, _17528_);
  and _68920_ (_17531_, _17530_, _04444_);
  nor _68921_ (_17533_, _12930_, _08737_);
  nor _68922_ (_17534_, _17533_, _17518_);
  nor _68923_ (_17535_, _17534_, _04444_);
  or _68924_ (_17536_, _17535_, _17531_);
  and _68925_ (_17537_, _17536_, _03983_);
  nor _68926_ (_17538_, _17524_, _03983_);
  nor _68927_ (_17539_, _17538_, _17537_);
  nor _68928_ (_17540_, _17539_, _03575_);
  nor _68929_ (_17541_, _17527_, _03583_);
  nor _68930_ (_17542_, _17541_, _07314_);
  not _68931_ (_17544_, _17542_);
  nor _68932_ (_17545_, _17544_, _17540_);
  nor _68933_ (_17546_, _17545_, _17525_);
  nor _68934_ (_17547_, _17546_, _03479_);
  and _68935_ (_17548_, _06721_, _05185_);
  nor _68936_ (_17549_, _17518_, _06044_);
  not _68937_ (_17550_, _17549_);
  nor _68938_ (_17551_, _17550_, _17548_);
  or _68939_ (_17552_, _17551_, _03221_);
  nor _68940_ (_17553_, _17552_, _17547_);
  nor _68941_ (_17555_, _13021_, _08737_);
  nor _68942_ (_17556_, _17555_, _17518_);
  nor _68943_ (_17557_, _17556_, _03474_);
  or _68944_ (_17558_, _17557_, _03437_);
  or _68945_ (_17559_, _17558_, _17553_);
  and _68946_ (_17560_, _06211_, _05185_);
  nor _68947_ (_17561_, _17560_, _17518_);
  nand _68948_ (_17562_, _17561_, _03437_);
  and _68949_ (_17563_, _17562_, _17559_);
  nor _68950_ (_17564_, _17563_, _03636_);
  and _68951_ (_17566_, _13036_, _05185_);
  or _68952_ (_17567_, _17518_, _04499_);
  nor _68953_ (_17568_, _17567_, _17566_);
  or _68954_ (_17569_, _17568_, _03769_);
  nor _68955_ (_17570_, _17569_, _17564_);
  nor _68956_ (_17571_, _17570_, _17522_);
  nor _68957_ (_17572_, _17571_, _04504_);
  not _68958_ (_17573_, _17518_);
  and _68959_ (_17574_, _17573_, _05471_);
  or _68960_ (_17575_, _17561_, _04505_);
  nor _68961_ (_17577_, _17575_, _17574_);
  nor _68962_ (_17578_, _17577_, _17572_);
  nor _68963_ (_17579_, _17578_, _03752_);
  or _68964_ (_17580_, _17574_, _03753_);
  or _68965_ (_17581_, _17580_, _17527_);
  and _68966_ (_17582_, _17581_, _03759_);
  not _68967_ (_17583_, _17582_);
  nor _68968_ (_17584_, _17583_, _17579_);
  nor _68969_ (_17585_, _13035_, _08737_);
  or _68970_ (_17586_, _17518_, _03759_);
  nor _68971_ (_17588_, _17586_, _17585_);
  or _68972_ (_17589_, _17588_, _03760_);
  nor _68973_ (_17590_, _17589_, _17584_);
  nor _68974_ (_17591_, _13041_, _08737_);
  nor _68975_ (_17592_, _17591_, _17518_);
  nor _68976_ (_17593_, _17592_, _04517_);
  or _68977_ (_17594_, _17593_, _03790_);
  nor _68978_ (_17595_, _17594_, _17590_);
  and _68979_ (_17596_, _17534_, _03790_);
  or _68980_ (_17597_, _17596_, _03520_);
  nor _68981_ (_17599_, _17597_, _17595_);
  and _68982_ (_17600_, _13097_, _05185_);
  nor _68983_ (_17601_, _17600_, _17518_);
  nor _68984_ (_17602_, _17601_, _03521_);
  or _68985_ (_17603_, _17602_, _17599_);
  or _68986_ (_17604_, _17603_, _42967_);
  or _68987_ (_17605_, _42963_, \oc8051_golden_model_1.SBUF [5]);
  and _68988_ (_17606_, _17605_, _41755_);
  and _68989_ (_43217_, _17606_, _17604_);
  not _68990_ (_17607_, \oc8051_golden_model_1.SBUF [6]);
  nor _68991_ (_17609_, _05185_, _17607_);
  and _68992_ (_17610_, _13259_, _05185_);
  nor _68993_ (_17611_, _17610_, _17609_);
  nor _68994_ (_17612_, _17611_, _04501_);
  and _68995_ (_17613_, _05185_, \oc8051_golden_model_1.ACC [6]);
  nor _68996_ (_17614_, _17613_, _17609_);
  nor _68997_ (_17615_, _17614_, _03583_);
  nor _68998_ (_17616_, _17614_, _04427_);
  nor _68999_ (_17617_, _04426_, _17607_);
  or _69000_ (_17618_, _17617_, _17616_);
  and _69001_ (_17620_, _17618_, _04444_);
  nor _69002_ (_17621_, _13122_, _08737_);
  nor _69003_ (_17622_, _17621_, _17609_);
  nor _69004_ (_17623_, _17622_, _04444_);
  or _69005_ (_17624_, _17623_, _17620_);
  and _69006_ (_17625_, _17624_, _03983_);
  nor _69007_ (_17626_, _05327_, _08737_);
  nor _69008_ (_17627_, _17626_, _17609_);
  nor _69009_ (_17628_, _17627_, _03983_);
  nor _69010_ (_17629_, _17628_, _17625_);
  nor _69011_ (_17631_, _17629_, _03575_);
  or _69012_ (_17632_, _17631_, _07314_);
  nor _69013_ (_17633_, _17632_, _17615_);
  and _69014_ (_17634_, _17627_, _07314_);
  nor _69015_ (_17635_, _17634_, _17633_);
  nor _69016_ (_17636_, _17635_, _03479_);
  and _69017_ (_17637_, _06713_, _05185_);
  nor _69018_ (_17638_, _17609_, _06044_);
  not _69019_ (_17639_, _17638_);
  nor _69020_ (_17640_, _17639_, _17637_);
  or _69021_ (_17642_, _17640_, _03221_);
  nor _69022_ (_17643_, _17642_, _17636_);
  nor _69023_ (_17644_, _13237_, _08737_);
  nor _69024_ (_17645_, _17644_, _17609_);
  nor _69025_ (_17646_, _17645_, _03474_);
  or _69026_ (_17647_, _17646_, _03437_);
  or _69027_ (_17648_, _17647_, _17643_);
  and _69028_ (_17649_, _13244_, _05185_);
  nor _69029_ (_17650_, _17649_, _17609_);
  nand _69030_ (_17651_, _17650_, _03437_);
  and _69031_ (_17653_, _17651_, _17648_);
  nor _69032_ (_17654_, _17653_, _03636_);
  and _69033_ (_17655_, _13253_, _05185_);
  or _69034_ (_17656_, _17609_, _04499_);
  nor _69035_ (_17657_, _17656_, _17655_);
  or _69036_ (_17658_, _17657_, _03769_);
  nor _69037_ (_17659_, _17658_, _17654_);
  nor _69038_ (_17660_, _17659_, _17612_);
  nor _69039_ (_17661_, _17660_, _04504_);
  not _69040_ (_17662_, _17609_);
  and _69041_ (_17664_, _17662_, _05376_);
  or _69042_ (_17665_, _17650_, _04505_);
  nor _69043_ (_17666_, _17665_, _17664_);
  nor _69044_ (_17667_, _17666_, _17661_);
  nor _69045_ (_17668_, _17667_, _03752_);
  or _69046_ (_17669_, _17664_, _03753_);
  or _69047_ (_17670_, _17669_, _17614_);
  and _69048_ (_17671_, _17670_, _03759_);
  not _69049_ (_17672_, _17671_);
  nor _69050_ (_17673_, _17672_, _17668_);
  nor _69051_ (_17675_, _13251_, _08737_);
  or _69052_ (_17676_, _17609_, _03759_);
  nor _69053_ (_17677_, _17676_, _17675_);
  or _69054_ (_17678_, _17677_, _03760_);
  nor _69055_ (_17679_, _17678_, _17673_);
  nor _69056_ (_17680_, _13258_, _08737_);
  nor _69057_ (_17681_, _17680_, _17609_);
  nor _69058_ (_17682_, _17681_, _04517_);
  or _69059_ (_17683_, _17682_, _03790_);
  nor _69060_ (_17684_, _17683_, _17679_);
  and _69061_ (_17686_, _17622_, _03790_);
  or _69062_ (_17687_, _17686_, _03520_);
  nor _69063_ (_17688_, _17687_, _17684_);
  and _69064_ (_17689_, _13312_, _05185_);
  nor _69065_ (_17690_, _17689_, _17609_);
  nor _69066_ (_17691_, _17690_, _03521_);
  or _69067_ (_17692_, _17691_, _17688_);
  or _69068_ (_17693_, _17692_, _42967_);
  or _69069_ (_17694_, _42963_, \oc8051_golden_model_1.SBUF [6]);
  and _69070_ (_17695_, _17694_, _41755_);
  and _69071_ (_43218_, _17695_, _17693_);
  not _69072_ (_17697_, \oc8051_golden_model_1.SCON [0]);
  nor _69073_ (_17698_, _05248_, _17697_);
  and _69074_ (_17699_, _11995_, _05248_);
  nor _69075_ (_17700_, _17699_, _17698_);
  nor _69076_ (_17701_, _17700_, _04501_);
  and _69077_ (_17702_, _05248_, _04419_);
  nor _69078_ (_17703_, _17702_, _17698_);
  and _69079_ (_17704_, _17703_, _07314_);
  and _69080_ (_17705_, _05248_, \oc8051_golden_model_1.ACC [0]);
  nor _69081_ (_17707_, _17705_, _17698_);
  nor _69082_ (_17708_, _17707_, _04427_);
  nor _69083_ (_17709_, _04426_, _17697_);
  or _69084_ (_17710_, _17709_, _17708_);
  and _69085_ (_17711_, _17710_, _04444_);
  and _69086_ (_17712_, _05941_, _05248_);
  nor _69087_ (_17713_, _17712_, _17698_);
  nor _69088_ (_17714_, _17713_, _04444_);
  or _69089_ (_17715_, _17714_, _17711_);
  and _69090_ (_17716_, _17715_, _03517_);
  nor _69091_ (_17718_, _05805_, _17697_);
  and _69092_ (_17719_, _11887_, _05805_);
  nor _69093_ (_17720_, _17719_, _17718_);
  nor _69094_ (_17721_, _17720_, _03517_);
  nor _69095_ (_17722_, _17721_, _17716_);
  nor _69096_ (_17723_, _17722_, _03568_);
  nor _69097_ (_17724_, _17703_, _03983_);
  or _69098_ (_17725_, _17724_, _17723_);
  and _69099_ (_17726_, _17725_, _03583_);
  nor _69100_ (_17727_, _17707_, _03583_);
  or _69101_ (_17729_, _17727_, _17726_);
  and _69102_ (_17730_, _17729_, _03513_);
  and _69103_ (_17731_, _17698_, _03512_);
  or _69104_ (_17732_, _17731_, _17730_);
  and _69105_ (_17733_, _17732_, _03506_);
  nor _69106_ (_17734_, _17713_, _03506_);
  or _69107_ (_17735_, _17734_, _17733_);
  and _69108_ (_17736_, _17735_, _03500_);
  nor _69109_ (_17737_, _11916_, _08855_);
  nor _69110_ (_17738_, _17737_, _17718_);
  nor _69111_ (_17740_, _17738_, _03500_);
  or _69112_ (_17741_, _17740_, _07314_);
  nor _69113_ (_17742_, _17741_, _17736_);
  nor _69114_ (_17743_, _17742_, _17704_);
  nor _69115_ (_17744_, _17743_, _03479_);
  and _69116_ (_17745_, _06715_, _05248_);
  nor _69117_ (_17746_, _17698_, _06044_);
  not _69118_ (_17747_, _17746_);
  nor _69119_ (_17748_, _17747_, _17745_);
  or _69120_ (_17749_, _17748_, _03221_);
  nor _69121_ (_17751_, _17749_, _17744_);
  nor _69122_ (_17752_, _11975_, _08818_);
  nor _69123_ (_17753_, _17752_, _17698_);
  nor _69124_ (_17754_, _17753_, _03474_);
  or _69125_ (_17755_, _17754_, _03437_);
  or _69126_ (_17756_, _17755_, _17751_);
  and _69127_ (_17757_, _05248_, _06202_);
  nor _69128_ (_17758_, _17757_, _17698_);
  nand _69129_ (_17759_, _17758_, _03437_);
  and _69130_ (_17760_, _17759_, _17756_);
  nor _69131_ (_17762_, _17760_, _03636_);
  and _69132_ (_17763_, _11990_, _05248_);
  or _69133_ (_17764_, _17698_, _04499_);
  nor _69134_ (_17765_, _17764_, _17763_);
  or _69135_ (_17766_, _17765_, _03769_);
  nor _69136_ (_17767_, _17766_, _17762_);
  nor _69137_ (_17768_, _17767_, _17701_);
  nor _69138_ (_17769_, _17768_, _04504_);
  or _69139_ (_17770_, _17758_, _04505_);
  nor _69140_ (_17771_, _17770_, _17712_);
  nor _69141_ (_17773_, _17771_, _17769_);
  nor _69142_ (_17774_, _17773_, _03752_);
  and _69143_ (_17775_, _11994_, _05248_);
  or _69144_ (_17776_, _17775_, _17698_);
  and _69145_ (_17777_, _17776_, _03752_);
  or _69146_ (_17778_, _17777_, _17774_);
  and _69147_ (_17779_, _17778_, _03759_);
  nor _69148_ (_17780_, _11988_, _08818_);
  nor _69149_ (_17781_, _17780_, _17698_);
  nor _69150_ (_17782_, _17781_, _03759_);
  or _69151_ (_17784_, _17782_, _17779_);
  and _69152_ (_17785_, _17784_, _04517_);
  nor _69153_ (_17786_, _11870_, _08818_);
  nor _69154_ (_17787_, _17786_, _17698_);
  nor _69155_ (_17788_, _17787_, _04517_);
  or _69156_ (_17789_, _17788_, _17785_);
  and _69157_ (_17790_, _17789_, _04192_);
  nor _69158_ (_17791_, _17713_, _04192_);
  or _69159_ (_17792_, _17791_, _17790_);
  and _69160_ (_17793_, _17792_, _03152_);
  and _69161_ (_17795_, _17698_, _03151_);
  nor _69162_ (_17796_, _17795_, _17793_);
  or _69163_ (_17797_, _17796_, _03520_);
  or _69164_ (_17798_, _17713_, _03521_);
  and _69165_ (_17799_, _17798_, _17797_);
  nand _69166_ (_17800_, _17799_, _42963_);
  or _69167_ (_17801_, _42963_, \oc8051_golden_model_1.SCON [0]);
  and _69168_ (_17802_, _17801_, _41755_);
  and _69169_ (_43219_, _17802_, _17800_);
  not _69170_ (_17803_, \oc8051_golden_model_1.SCON [1]);
  nor _69171_ (_17805_, _05248_, _17803_);
  and _69172_ (_17806_, _06714_, _05248_);
  or _69173_ (_17807_, _17806_, _17805_);
  and _69174_ (_17808_, _17807_, _03479_);
  nor _69175_ (_17809_, _05248_, \oc8051_golden_model_1.SCON [1]);
  and _69176_ (_17810_, _05248_, _03233_);
  nor _69177_ (_17811_, _17810_, _17809_);
  and _69178_ (_17812_, _17811_, _04426_);
  nor _69179_ (_17813_, _04426_, _17803_);
  or _69180_ (_17814_, _17813_, _17812_);
  and _69181_ (_17816_, _17814_, _04444_);
  and _69182_ (_17817_, _12252_, _05248_);
  nor _69183_ (_17818_, _17817_, _17809_);
  and _69184_ (_17819_, _17818_, _03570_);
  or _69185_ (_17820_, _17819_, _17816_);
  and _69186_ (_17821_, _17820_, _03517_);
  and _69187_ (_17822_, _12083_, _05805_);
  nor _69188_ (_17823_, _05805_, _17803_);
  or _69189_ (_17824_, _17823_, _03568_);
  or _69190_ (_17825_, _17824_, _17822_);
  and _69191_ (_17827_, _17825_, _14165_);
  nor _69192_ (_17828_, _17827_, _17821_);
  nor _69193_ (_17829_, _08818_, _04603_);
  nor _69194_ (_17830_, _17829_, _17805_);
  and _69195_ (_17831_, _17830_, _03568_);
  nor _69196_ (_17832_, _17831_, _17828_);
  and _69197_ (_17833_, _17832_, _03583_);
  and _69198_ (_17834_, _17811_, _03575_);
  or _69199_ (_17835_, _17834_, _17833_);
  and _69200_ (_17836_, _17835_, _03513_);
  and _69201_ (_17838_, _12069_, _05805_);
  nor _69202_ (_17839_, _17838_, _17823_);
  nor _69203_ (_17840_, _17839_, _03513_);
  or _69204_ (_17841_, _17840_, _17836_);
  and _69205_ (_17842_, _17841_, _03506_);
  and _69206_ (_17843_, _17822_, _12098_);
  or _69207_ (_17844_, _17843_, _17823_);
  and _69208_ (_17845_, _17844_, _03505_);
  or _69209_ (_17846_, _17845_, _17842_);
  and _69210_ (_17847_, _17846_, _03500_);
  nor _69211_ (_17849_, _12116_, _08855_);
  nor _69212_ (_17850_, _17823_, _17849_);
  nor _69213_ (_17851_, _17850_, _03500_);
  or _69214_ (_17852_, _17851_, _07314_);
  nor _69215_ (_17853_, _17852_, _17847_);
  and _69216_ (_17854_, _17830_, _07314_);
  or _69217_ (_17855_, _17854_, _03479_);
  nor _69218_ (_17856_, _17855_, _17853_);
  or _69219_ (_17857_, _17856_, _17808_);
  and _69220_ (_17858_, _17857_, _03474_);
  nor _69221_ (_17860_, _12176_, _08818_);
  nor _69222_ (_17861_, _17860_, _17805_);
  nor _69223_ (_17862_, _17861_, _03474_);
  nor _69224_ (_17863_, _17862_, _17858_);
  nor _69225_ (_17864_, _17863_, _03437_);
  and _69226_ (_17865_, _05248_, _04317_);
  not _69227_ (_17866_, _17865_);
  nor _69228_ (_17867_, _17809_, _03438_);
  and _69229_ (_17868_, _17867_, _17866_);
  nor _69230_ (_17869_, _17868_, _17864_);
  nor _69231_ (_17871_, _17869_, _03636_);
  not _69232_ (_17872_, _17809_);
  nor _69233_ (_17873_, _12191_, _08818_);
  nor _69234_ (_17874_, _17873_, _04499_);
  and _69235_ (_17875_, _17874_, _17872_);
  nor _69236_ (_17876_, _17875_, _17871_);
  nor _69237_ (_17877_, _17876_, _03769_);
  nor _69238_ (_17878_, _12197_, _08818_);
  nor _69239_ (_17879_, _17878_, _04501_);
  and _69240_ (_17880_, _17879_, _17872_);
  nor _69241_ (_17882_, _17880_, _17877_);
  nor _69242_ (_17883_, _17882_, _04504_);
  nor _69243_ (_17884_, _12190_, _08818_);
  nor _69244_ (_17885_, _17884_, _05769_);
  and _69245_ (_17886_, _17885_, _17872_);
  nor _69246_ (_17887_, _17886_, _17883_);
  nor _69247_ (_17888_, _17887_, _03752_);
  nor _69248_ (_17889_, _17805_, _05569_);
  nor _69249_ (_17890_, _17889_, _03753_);
  and _69250_ (_17891_, _17890_, _17811_);
  nor _69251_ (_17893_, _17891_, _17888_);
  nor _69252_ (_17894_, _17893_, _03758_);
  and _69253_ (_17895_, _17865_, _05940_);
  nor _69254_ (_17896_, _17895_, _03759_);
  and _69255_ (_17897_, _17896_, _17872_);
  nor _69256_ (_17898_, _17897_, _17894_);
  nor _69257_ (_17899_, _17898_, _03760_);
  and _69258_ (_17900_, _17810_, _05940_);
  nor _69259_ (_17901_, _17900_, _04517_);
  and _69260_ (_17902_, _17901_, _17872_);
  or _69261_ (_17904_, _17902_, _17899_);
  and _69262_ (_17905_, _17904_, _04192_);
  and _69263_ (_17906_, _17818_, _03790_);
  or _69264_ (_17907_, _17906_, _17905_);
  and _69265_ (_17908_, _17907_, _03152_);
  nor _69266_ (_17909_, _17839_, _03152_);
  or _69267_ (_17910_, _17909_, _03520_);
  nor _69268_ (_17911_, _17910_, _17908_);
  nor _69269_ (_17912_, _17817_, _17805_);
  and _69270_ (_17913_, _17912_, _03520_);
  nor _69271_ (_17915_, _17913_, _17911_);
  or _69272_ (_17916_, _17915_, _42967_);
  or _69273_ (_17917_, _42963_, \oc8051_golden_model_1.SCON [1]);
  and _69274_ (_17918_, _17917_, _41755_);
  and _69275_ (_43222_, _17918_, _17916_);
  not _69276_ (_17919_, \oc8051_golden_model_1.SCON [2]);
  nor _69277_ (_17920_, _05248_, _17919_);
  and _69278_ (_17921_, _12401_, _05248_);
  nor _69279_ (_17922_, _17921_, _17920_);
  nor _69280_ (_17923_, _17922_, _04501_);
  nor _69281_ (_17925_, _08818_, _05026_);
  nor _69282_ (_17926_, _17925_, _17920_);
  and _69283_ (_17927_, _17926_, _07314_);
  nor _69284_ (_17928_, _17926_, _03983_);
  nor _69285_ (_17929_, _05805_, _17919_);
  and _69286_ (_17930_, _12278_, _05805_);
  nor _69287_ (_17931_, _17930_, _17929_);
  and _69288_ (_17932_, _17931_, _03516_);
  nor _69289_ (_17933_, _12282_, _08818_);
  nor _69290_ (_17934_, _17933_, _17920_);
  nor _69291_ (_17936_, _17934_, _04444_);
  nor _69292_ (_17937_, _04426_, _17919_);
  and _69293_ (_17938_, _05248_, \oc8051_golden_model_1.ACC [2]);
  nor _69294_ (_17939_, _17938_, _17920_);
  nor _69295_ (_17940_, _17939_, _04427_);
  nor _69296_ (_17941_, _17940_, _17937_);
  nor _69297_ (_17942_, _17941_, _03570_);
  or _69298_ (_17943_, _17942_, _03516_);
  nor _69299_ (_17944_, _17943_, _17936_);
  nor _69300_ (_17945_, _17944_, _17932_);
  and _69301_ (_17947_, _17945_, _03983_);
  or _69302_ (_17948_, _17947_, _17928_);
  and _69303_ (_17949_, _17948_, _03583_);
  nor _69304_ (_17950_, _17939_, _03583_);
  or _69305_ (_17951_, _17950_, _17949_);
  and _69306_ (_17952_, _17951_, _03513_);
  and _69307_ (_17953_, _12276_, _05805_);
  nor _69308_ (_17954_, _17953_, _17929_);
  nor _69309_ (_17955_, _17954_, _03513_);
  or _69310_ (_17956_, _17955_, _17952_);
  and _69311_ (_17958_, _17956_, _03506_);
  nor _69312_ (_17959_, _17929_, _12309_);
  nor _69313_ (_17960_, _17959_, _17931_);
  and _69314_ (_17961_, _17960_, _03505_);
  or _69315_ (_17962_, _17961_, _17958_);
  and _69316_ (_17963_, _17962_, _03500_);
  nor _69317_ (_17964_, _12326_, _08855_);
  nor _69318_ (_17965_, _17964_, _17929_);
  nor _69319_ (_17966_, _17965_, _03500_);
  nor _69320_ (_17967_, _17966_, _07314_);
  not _69321_ (_17969_, _17967_);
  nor _69322_ (_17970_, _17969_, _17963_);
  nor _69323_ (_17971_, _17970_, _17927_);
  nor _69324_ (_17972_, _17971_, _03479_);
  and _69325_ (_17973_, _06718_, _05248_);
  nor _69326_ (_17974_, _17920_, _06044_);
  not _69327_ (_17975_, _17974_);
  nor _69328_ (_17976_, _17975_, _17973_);
  or _69329_ (_17977_, _17976_, _03221_);
  nor _69330_ (_17978_, _17977_, _17972_);
  nor _69331_ (_17980_, _12384_, _08818_);
  nor _69332_ (_17981_, _17980_, _17920_);
  nor _69333_ (_17982_, _17981_, _03474_);
  or _69334_ (_17983_, _17982_, _03437_);
  or _69335_ (_17984_, _17983_, _17978_);
  and _69336_ (_17985_, _05248_, _06261_);
  nor _69337_ (_17986_, _17985_, _17920_);
  nand _69338_ (_17987_, _17986_, _03437_);
  and _69339_ (_17988_, _17987_, _17984_);
  nor _69340_ (_17989_, _17988_, _03636_);
  and _69341_ (_17991_, _12273_, _05248_);
  or _69342_ (_17992_, _17920_, _04499_);
  nor _69343_ (_17993_, _17992_, _17991_);
  or _69344_ (_17994_, _17993_, _03769_);
  nor _69345_ (_17995_, _17994_, _17989_);
  nor _69346_ (_17996_, _17995_, _17923_);
  nor _69347_ (_17997_, _17996_, _04504_);
  not _69348_ (_17998_, _17920_);
  and _69349_ (_17999_, _17998_, _05664_);
  or _69350_ (_18000_, _17986_, _04505_);
  nor _69351_ (_18002_, _18000_, _17999_);
  nor _69352_ (_18003_, _18002_, _17997_);
  nor _69353_ (_18004_, _18003_, _03752_);
  or _69354_ (_18005_, _17999_, _03753_);
  nor _69355_ (_18006_, _18005_, _17939_);
  or _69356_ (_18007_, _18006_, _18004_);
  and _69357_ (_18008_, _18007_, _03759_);
  nor _69358_ (_18009_, _12272_, _08818_);
  nor _69359_ (_18010_, _18009_, _17920_);
  nor _69360_ (_18011_, _18010_, _03759_);
  or _69361_ (_18013_, _18011_, _18008_);
  and _69362_ (_18014_, _18013_, _04517_);
  nor _69363_ (_18015_, _12400_, _08818_);
  nor _69364_ (_18016_, _18015_, _17920_);
  nor _69365_ (_18017_, _18016_, _04517_);
  or _69366_ (_18018_, _18017_, _18014_);
  and _69367_ (_18019_, _18018_, _04192_);
  nor _69368_ (_18020_, _17934_, _04192_);
  or _69369_ (_18021_, _18020_, _18019_);
  and _69370_ (_18022_, _18021_, _03152_);
  nor _69371_ (_18024_, _17954_, _03152_);
  or _69372_ (_18025_, _18024_, _18022_);
  and _69373_ (_18026_, _18025_, _03521_);
  and _69374_ (_18027_, _12456_, _05248_);
  nor _69375_ (_18028_, _18027_, _17920_);
  nor _69376_ (_18029_, _18028_, _03521_);
  or _69377_ (_18030_, _18029_, _18026_);
  or _69378_ (_18031_, _18030_, _42967_);
  or _69379_ (_18032_, _42963_, \oc8051_golden_model_1.SCON [2]);
  and _69380_ (_18033_, _18032_, _41755_);
  and _69381_ (_43223_, _18033_, _18031_);
  not _69382_ (_18035_, \oc8051_golden_model_1.SCON [3]);
  nor _69383_ (_18036_, _05248_, _18035_);
  and _69384_ (_18037_, _12604_, _05248_);
  nor _69385_ (_18038_, _18037_, _18036_);
  nor _69386_ (_18039_, _18038_, _04501_);
  nor _69387_ (_18040_, _08818_, _04843_);
  nor _69388_ (_18041_, _18040_, _18036_);
  and _69389_ (_18042_, _18041_, _07314_);
  and _69390_ (_18043_, _05248_, \oc8051_golden_model_1.ACC [3]);
  nor _69391_ (_18045_, _18043_, _18036_);
  nor _69392_ (_18046_, _18045_, _04427_);
  nor _69393_ (_18047_, _04426_, _18035_);
  or _69394_ (_18048_, _18047_, _18046_);
  and _69395_ (_18049_, _18048_, _04444_);
  nor _69396_ (_18050_, _12486_, _08818_);
  nor _69397_ (_18051_, _18050_, _18036_);
  nor _69398_ (_18052_, _18051_, _04444_);
  or _69399_ (_18053_, _18052_, _18049_);
  and _69400_ (_18054_, _18053_, _03517_);
  nor _69401_ (_18056_, _05805_, _18035_);
  and _69402_ (_18057_, _12490_, _05805_);
  nor _69403_ (_18058_, _18057_, _18056_);
  nor _69404_ (_18059_, _18058_, _03517_);
  or _69405_ (_18060_, _18059_, _03568_);
  or _69406_ (_18061_, _18060_, _18054_);
  nand _69407_ (_18062_, _18041_, _03568_);
  and _69408_ (_18063_, _18062_, _18061_);
  and _69409_ (_18064_, _18063_, _03583_);
  nor _69410_ (_18065_, _18045_, _03583_);
  or _69411_ (_18067_, _18065_, _18064_);
  and _69412_ (_18068_, _18067_, _03513_);
  and _69413_ (_18069_, _12500_, _05805_);
  nor _69414_ (_18070_, _18069_, _18056_);
  nor _69415_ (_18071_, _18070_, _03513_);
  or _69416_ (_18072_, _18071_, _03505_);
  or _69417_ (_18073_, _18072_, _18068_);
  nor _69418_ (_18074_, _18056_, _12507_);
  nor _69419_ (_18075_, _18074_, _18058_);
  or _69420_ (_18076_, _18075_, _03506_);
  and _69421_ (_18078_, _18076_, _03500_);
  and _69422_ (_18079_, _18078_, _18073_);
  nor _69423_ (_18080_, _12525_, _08855_);
  nor _69424_ (_18081_, _18080_, _18056_);
  nor _69425_ (_18082_, _18081_, _03500_);
  nor _69426_ (_18083_, _18082_, _07314_);
  not _69427_ (_18084_, _18083_);
  nor _69428_ (_18085_, _18084_, _18079_);
  nor _69429_ (_18086_, _18085_, _18042_);
  nor _69430_ (_18087_, _18086_, _03479_);
  and _69431_ (_18089_, _06717_, _05248_);
  nor _69432_ (_18090_, _18036_, _06044_);
  not _69433_ (_18091_, _18090_);
  nor _69434_ (_18092_, _18091_, _18089_);
  or _69435_ (_18093_, _18092_, _03221_);
  nor _69436_ (_18094_, _18093_, _18087_);
  nor _69437_ (_18095_, _12583_, _08818_);
  nor _69438_ (_18096_, _18095_, _18036_);
  nor _69439_ (_18097_, _18096_, _03474_);
  or _69440_ (_18098_, _18097_, _03437_);
  or _69441_ (_18100_, _18098_, _18094_);
  and _69442_ (_18101_, _05248_, _06217_);
  nor _69443_ (_18102_, _18101_, _18036_);
  nand _69444_ (_18103_, _18102_, _03437_);
  and _69445_ (_18104_, _18103_, _18100_);
  nor _69446_ (_18105_, _18104_, _03636_);
  and _69447_ (_18106_, _12598_, _05248_);
  or _69448_ (_18107_, _18036_, _04499_);
  nor _69449_ (_18108_, _18107_, _18106_);
  or _69450_ (_18109_, _18108_, _03769_);
  nor _69451_ (_18111_, _18109_, _18105_);
  nor _69452_ (_18112_, _18111_, _18039_);
  nor _69453_ (_18113_, _18112_, _04504_);
  not _69454_ (_18114_, _18036_);
  and _69455_ (_18115_, _18114_, _05520_);
  or _69456_ (_18116_, _18102_, _04505_);
  nor _69457_ (_18117_, _18116_, _18115_);
  nor _69458_ (_18118_, _18117_, _18113_);
  nor _69459_ (_18119_, _18118_, _03752_);
  or _69460_ (_18120_, _18115_, _03753_);
  or _69461_ (_18122_, _18120_, _18045_);
  and _69462_ (_18123_, _18122_, _03759_);
  not _69463_ (_18124_, _18123_);
  nor _69464_ (_18125_, _18124_, _18119_);
  nor _69465_ (_18126_, _12597_, _08818_);
  or _69466_ (_18127_, _18036_, _03759_);
  nor _69467_ (_18128_, _18127_, _18126_);
  or _69468_ (_18129_, _18128_, _03760_);
  nor _69469_ (_18130_, _18129_, _18125_);
  nor _69470_ (_18131_, _12603_, _08818_);
  nor _69471_ (_18133_, _18131_, _18036_);
  nor _69472_ (_18134_, _18133_, _04517_);
  or _69473_ (_18135_, _18134_, _18130_);
  and _69474_ (_18136_, _18135_, _04192_);
  nor _69475_ (_18137_, _18051_, _04192_);
  or _69476_ (_18138_, _18137_, _18136_);
  and _69477_ (_18139_, _18138_, _03152_);
  nor _69478_ (_18140_, _18070_, _03152_);
  or _69479_ (_18141_, _18140_, _18139_);
  and _69480_ (_18142_, _18141_, _03521_);
  and _69481_ (_18144_, _12658_, _05248_);
  nor _69482_ (_18145_, _18144_, _18036_);
  nor _69483_ (_18146_, _18145_, _03521_);
  or _69484_ (_18147_, _18146_, _18142_);
  or _69485_ (_18148_, _18147_, _42967_);
  or _69486_ (_18149_, _42963_, \oc8051_golden_model_1.SCON [3]);
  and _69487_ (_18150_, _18149_, _41755_);
  and _69488_ (_43224_, _18150_, _18148_);
  not _69489_ (_18151_, \oc8051_golden_model_1.SCON [4]);
  nor _69490_ (_18152_, _05248_, _18151_);
  and _69491_ (_18154_, _12844_, _05248_);
  nor _69492_ (_18155_, _18154_, _18152_);
  nor _69493_ (_18156_, _18155_, _04501_);
  nor _69494_ (_18157_, _05712_, _08818_);
  nor _69495_ (_18158_, _18157_, _18152_);
  and _69496_ (_18159_, _18158_, _07314_);
  and _69497_ (_18160_, _05248_, \oc8051_golden_model_1.ACC [4]);
  nor _69498_ (_18161_, _18160_, _18152_);
  nor _69499_ (_18162_, _18161_, _04427_);
  nor _69500_ (_18163_, _04426_, _18151_);
  or _69501_ (_18165_, _18163_, _18162_);
  and _69502_ (_18166_, _18165_, _04444_);
  nor _69503_ (_18167_, _12733_, _08818_);
  nor _69504_ (_18168_, _18167_, _18152_);
  nor _69505_ (_18169_, _18168_, _04444_);
  or _69506_ (_18170_, _18169_, _18166_);
  and _69507_ (_18171_, _18170_, _03517_);
  nor _69508_ (_18172_, _05805_, _18151_);
  and _69509_ (_18173_, _12737_, _05805_);
  nor _69510_ (_18174_, _18173_, _18172_);
  nor _69511_ (_18176_, _18174_, _03517_);
  or _69512_ (_18177_, _18176_, _03568_);
  or _69513_ (_18178_, _18177_, _18171_);
  nand _69514_ (_18179_, _18158_, _03568_);
  and _69515_ (_18180_, _18179_, _18178_);
  and _69516_ (_18181_, _18180_, _03583_);
  nor _69517_ (_18182_, _18161_, _03583_);
  or _69518_ (_18183_, _18182_, _18181_);
  and _69519_ (_18184_, _18183_, _03513_);
  and _69520_ (_18185_, _12718_, _05805_);
  nor _69521_ (_18187_, _18185_, _18172_);
  nor _69522_ (_18188_, _18187_, _03513_);
  or _69523_ (_18189_, _18188_, _18184_);
  and _69524_ (_18190_, _18189_, _03506_);
  nor _69525_ (_18191_, _18172_, _12752_);
  nor _69526_ (_18192_, _18191_, _18174_);
  and _69527_ (_18193_, _18192_, _03505_);
  or _69528_ (_18194_, _18193_, _18190_);
  and _69529_ (_18195_, _18194_, _03500_);
  nor _69530_ (_18196_, _12716_, _08855_);
  nor _69531_ (_18198_, _18196_, _18172_);
  nor _69532_ (_18199_, _18198_, _03500_);
  nor _69533_ (_18200_, _18199_, _07314_);
  not _69534_ (_18201_, _18200_);
  nor _69535_ (_18202_, _18201_, _18195_);
  nor _69536_ (_18203_, _18202_, _18159_);
  nor _69537_ (_18204_, _18203_, _03479_);
  and _69538_ (_18205_, _06722_, _05248_);
  nor _69539_ (_18206_, _18152_, _06044_);
  not _69540_ (_18207_, _18206_);
  nor _69541_ (_18209_, _18207_, _18205_);
  or _69542_ (_18210_, _18209_, _03221_);
  nor _69543_ (_18211_, _18210_, _18204_);
  nor _69544_ (_18212_, _12827_, _08818_);
  nor _69545_ (_18213_, _18212_, _18152_);
  nor _69546_ (_18214_, _18213_, _03474_);
  or _69547_ (_18215_, _18214_, _03437_);
  or _69548_ (_18216_, _18215_, _18211_);
  and _69549_ (_18217_, _06233_, _05248_);
  nor _69550_ (_18218_, _18217_, _18152_);
  nand _69551_ (_18220_, _18218_, _03437_);
  and _69552_ (_18221_, _18220_, _18216_);
  nor _69553_ (_18222_, _18221_, _03636_);
  and _69554_ (_18223_, _12711_, _05248_);
  or _69555_ (_18224_, _18152_, _04499_);
  nor _69556_ (_18225_, _18224_, _18223_);
  or _69557_ (_18226_, _18225_, _03769_);
  nor _69558_ (_18227_, _18226_, _18222_);
  nor _69559_ (_18228_, _18227_, _18156_);
  nor _69560_ (_18229_, _18228_, _04504_);
  not _69561_ (_18231_, _18152_);
  and _69562_ (_18232_, _18231_, _05760_);
  or _69563_ (_18233_, _18218_, _04505_);
  nor _69564_ (_18234_, _18233_, _18232_);
  nor _69565_ (_18235_, _18234_, _18229_);
  nor _69566_ (_18236_, _18235_, _03752_);
  or _69567_ (_18237_, _18232_, _03753_);
  or _69568_ (_18238_, _18237_, _18161_);
  and _69569_ (_18239_, _18238_, _03759_);
  not _69570_ (_18240_, _18239_);
  nor _69571_ (_18242_, _18240_, _18236_);
  nor _69572_ (_18243_, _12710_, _08818_);
  or _69573_ (_18244_, _18152_, _03759_);
  nor _69574_ (_18245_, _18244_, _18243_);
  or _69575_ (_18246_, _18245_, _03760_);
  nor _69576_ (_18247_, _18246_, _18242_);
  nor _69577_ (_18248_, _12843_, _08818_);
  nor _69578_ (_18249_, _18248_, _18152_);
  nor _69579_ (_18250_, _18249_, _04517_);
  or _69580_ (_18251_, _18250_, _18247_);
  and _69581_ (_18253_, _18251_, _04192_);
  nor _69582_ (_18254_, _18168_, _04192_);
  or _69583_ (_18255_, _18254_, _18253_);
  and _69584_ (_18256_, _18255_, _03152_);
  nor _69585_ (_18257_, _18187_, _03152_);
  or _69586_ (_18258_, _18257_, _18256_);
  and _69587_ (_18259_, _18258_, _03521_);
  and _69588_ (_18260_, _12893_, _05248_);
  nor _69589_ (_18261_, _18260_, _18152_);
  nor _69590_ (_18262_, _18261_, _03521_);
  or _69591_ (_18264_, _18262_, _18259_);
  or _69592_ (_18265_, _18264_, _42967_);
  or _69593_ (_18266_, _42963_, \oc8051_golden_model_1.SCON [4]);
  and _69594_ (_18267_, _18266_, _41755_);
  and _69595_ (_43225_, _18267_, _18265_);
  not _69596_ (_18268_, \oc8051_golden_model_1.SCON [5]);
  nor _69597_ (_18269_, _05248_, _18268_);
  and _69598_ (_18270_, _13042_, _05248_);
  nor _69599_ (_18271_, _18270_, _18269_);
  nor _69600_ (_18272_, _18271_, _04501_);
  nor _69601_ (_18274_, _05422_, _08818_);
  nor _69602_ (_18275_, _18274_, _18269_);
  and _69603_ (_18276_, _18275_, _07314_);
  and _69604_ (_18277_, _05248_, \oc8051_golden_model_1.ACC [5]);
  nor _69605_ (_18278_, _18277_, _18269_);
  nor _69606_ (_18279_, _18278_, _04427_);
  nor _69607_ (_18280_, _04426_, _18268_);
  or _69608_ (_18281_, _18280_, _18279_);
  and _69609_ (_18282_, _18281_, _04444_);
  nor _69610_ (_18283_, _12930_, _08818_);
  nor _69611_ (_18285_, _18283_, _18269_);
  nor _69612_ (_18286_, _18285_, _04444_);
  or _69613_ (_18287_, _18286_, _18282_);
  and _69614_ (_18288_, _18287_, _03517_);
  nor _69615_ (_18289_, _05805_, _18268_);
  and _69616_ (_18290_, _12934_, _05805_);
  nor _69617_ (_18291_, _18290_, _18289_);
  nor _69618_ (_18292_, _18291_, _03517_);
  or _69619_ (_18293_, _18292_, _03568_);
  or _69620_ (_18294_, _18293_, _18288_);
  nand _69621_ (_18296_, _18275_, _03568_);
  and _69622_ (_18297_, _18296_, _18294_);
  and _69623_ (_18298_, _18297_, _03583_);
  nor _69624_ (_18299_, _18278_, _03583_);
  or _69625_ (_18300_, _18299_, _18298_);
  and _69626_ (_18301_, _18300_, _03513_);
  and _69627_ (_18302_, _12914_, _05805_);
  nor _69628_ (_18303_, _18302_, _18289_);
  nor _69629_ (_18304_, _18303_, _03513_);
  or _69630_ (_18305_, _18304_, _18301_);
  and _69631_ (_18307_, _18305_, _03506_);
  nor _69632_ (_18308_, _18289_, _12949_);
  nor _69633_ (_18309_, _18308_, _18291_);
  and _69634_ (_18310_, _18309_, _03505_);
  or _69635_ (_18311_, _18310_, _18307_);
  and _69636_ (_18312_, _18311_, _03500_);
  nor _69637_ (_18313_, _12912_, _08855_);
  nor _69638_ (_18314_, _18313_, _18289_);
  nor _69639_ (_18315_, _18314_, _03500_);
  nor _69640_ (_18316_, _18315_, _07314_);
  not _69641_ (_18318_, _18316_);
  nor _69642_ (_18319_, _18318_, _18312_);
  nor _69643_ (_18320_, _18319_, _18276_);
  nor _69644_ (_18321_, _18320_, _03479_);
  and _69645_ (_18322_, _06721_, _05248_);
  nor _69646_ (_18323_, _18269_, _06044_);
  not _69647_ (_18324_, _18323_);
  nor _69648_ (_18325_, _18324_, _18322_);
  or _69649_ (_18326_, _18325_, _03221_);
  nor _69650_ (_18327_, _18326_, _18321_);
  nor _69651_ (_18329_, _13021_, _08818_);
  nor _69652_ (_18330_, _18329_, _18269_);
  nor _69653_ (_18331_, _18330_, _03474_);
  or _69654_ (_18332_, _18331_, _03437_);
  or _69655_ (_18333_, _18332_, _18327_);
  and _69656_ (_18334_, _06211_, _05248_);
  nor _69657_ (_18335_, _18334_, _18269_);
  nand _69658_ (_18336_, _18335_, _03437_);
  and _69659_ (_18337_, _18336_, _18333_);
  nor _69660_ (_18338_, _18337_, _03636_);
  and _69661_ (_18340_, _13036_, _05248_);
  or _69662_ (_18341_, _18269_, _04499_);
  nor _69663_ (_18342_, _18341_, _18340_);
  or _69664_ (_18343_, _18342_, _03769_);
  nor _69665_ (_18344_, _18343_, _18338_);
  nor _69666_ (_18345_, _18344_, _18272_);
  nor _69667_ (_18346_, _18345_, _04504_);
  not _69668_ (_18347_, _18269_);
  and _69669_ (_18348_, _18347_, _05471_);
  or _69670_ (_18349_, _18335_, _04505_);
  nor _69671_ (_18351_, _18349_, _18348_);
  nor _69672_ (_18352_, _18351_, _18346_);
  nor _69673_ (_18353_, _18352_, _03752_);
  or _69674_ (_18354_, _18348_, _03753_);
  or _69675_ (_18355_, _18354_, _18278_);
  and _69676_ (_18356_, _18355_, _03759_);
  not _69677_ (_18357_, _18356_);
  nor _69678_ (_18358_, _18357_, _18353_);
  nor _69679_ (_18359_, _13035_, _08818_);
  or _69680_ (_18360_, _18269_, _03759_);
  nor _69681_ (_18362_, _18360_, _18359_);
  or _69682_ (_18363_, _18362_, _03760_);
  nor _69683_ (_18364_, _18363_, _18358_);
  nor _69684_ (_18365_, _13041_, _08818_);
  nor _69685_ (_18366_, _18365_, _18269_);
  nor _69686_ (_18367_, _18366_, _04517_);
  or _69687_ (_18368_, _18367_, _18364_);
  and _69688_ (_18369_, _18368_, _04192_);
  nor _69689_ (_18370_, _18285_, _04192_);
  or _69690_ (_18371_, _18370_, _18369_);
  and _69691_ (_18373_, _18371_, _03152_);
  nor _69692_ (_18374_, _18303_, _03152_);
  or _69693_ (_18375_, _18374_, _18373_);
  and _69694_ (_18376_, _18375_, _03521_);
  and _69695_ (_18377_, _13097_, _05248_);
  nor _69696_ (_18378_, _18377_, _18269_);
  nor _69697_ (_18379_, _18378_, _03521_);
  or _69698_ (_18380_, _18379_, _18376_);
  or _69699_ (_18381_, _18380_, _42967_);
  or _69700_ (_18382_, _42963_, \oc8051_golden_model_1.SCON [5]);
  and _69701_ (_18384_, _18382_, _41755_);
  and _69702_ (_43226_, _18384_, _18381_);
  not _69703_ (_18385_, \oc8051_golden_model_1.SCON [6]);
  nor _69704_ (_18386_, _05248_, _18385_);
  and _69705_ (_18387_, _13259_, _05248_);
  nor _69706_ (_18388_, _18387_, _18386_);
  nor _69707_ (_18389_, _18388_, _04501_);
  nor _69708_ (_18390_, _05327_, _08818_);
  nor _69709_ (_18391_, _18390_, _18386_);
  and _69710_ (_18392_, _18391_, _07314_);
  and _69711_ (_18394_, _05248_, \oc8051_golden_model_1.ACC [6]);
  nor _69712_ (_18395_, _18394_, _18386_);
  nor _69713_ (_18396_, _18395_, _04427_);
  nor _69714_ (_18397_, _04426_, _18385_);
  or _69715_ (_18398_, _18397_, _18396_);
  and _69716_ (_18399_, _18398_, _04444_);
  nor _69717_ (_18400_, _13122_, _08818_);
  nor _69718_ (_18401_, _18400_, _18386_);
  nor _69719_ (_18402_, _18401_, _04444_);
  or _69720_ (_18403_, _18402_, _18399_);
  and _69721_ (_18405_, _18403_, _03517_);
  nor _69722_ (_18406_, _05805_, _18385_);
  and _69723_ (_18407_, _13145_, _05805_);
  nor _69724_ (_18408_, _18407_, _18406_);
  nor _69725_ (_18409_, _18408_, _03517_);
  or _69726_ (_18410_, _18409_, _03568_);
  or _69727_ (_18411_, _18410_, _18405_);
  nand _69728_ (_18412_, _18391_, _03568_);
  and _69729_ (_18413_, _18412_, _18411_);
  and _69730_ (_18414_, _18413_, _03583_);
  nor _69731_ (_18416_, _18395_, _03583_);
  or _69732_ (_18417_, _18416_, _18414_);
  and _69733_ (_18418_, _18417_, _03513_);
  and _69734_ (_18419_, _13130_, _05805_);
  nor _69735_ (_18420_, _18419_, _18406_);
  nor _69736_ (_18421_, _18420_, _03513_);
  or _69737_ (_18422_, _18421_, _03505_);
  or _69738_ (_18423_, _18422_, _18418_);
  nor _69739_ (_18424_, _18406_, _13160_);
  nor _69740_ (_18425_, _18424_, _18408_);
  or _69741_ (_18427_, _18425_, _03506_);
  and _69742_ (_18428_, _18427_, _03500_);
  and _69743_ (_18429_, _18428_, _18423_);
  nor _69744_ (_18430_, _13178_, _08855_);
  nor _69745_ (_18431_, _18430_, _18406_);
  nor _69746_ (_18432_, _18431_, _03500_);
  nor _69747_ (_18433_, _18432_, _07314_);
  not _69748_ (_18434_, _18433_);
  nor _69749_ (_18435_, _18434_, _18429_);
  nor _69750_ (_18436_, _18435_, _18392_);
  nor _69751_ (_18438_, _18436_, _03479_);
  and _69752_ (_18439_, _06713_, _05248_);
  nor _69753_ (_18440_, _18386_, _06044_);
  not _69754_ (_18441_, _18440_);
  nor _69755_ (_18442_, _18441_, _18439_);
  or _69756_ (_18443_, _18442_, _03221_);
  nor _69757_ (_18444_, _18443_, _18438_);
  nor _69758_ (_18445_, _13237_, _08818_);
  nor _69759_ (_18446_, _18445_, _18386_);
  nor _69760_ (_18447_, _18446_, _03474_);
  or _69761_ (_18449_, _18447_, _03437_);
  or _69762_ (_18450_, _18449_, _18444_);
  and _69763_ (_18451_, _13244_, _05248_);
  nor _69764_ (_18452_, _18451_, _18386_);
  nand _69765_ (_18453_, _18452_, _03437_);
  and _69766_ (_18454_, _18453_, _18450_);
  nor _69767_ (_18455_, _18454_, _03636_);
  and _69768_ (_18456_, _13253_, _05248_);
  or _69769_ (_18457_, _18386_, _04499_);
  nor _69770_ (_18458_, _18457_, _18456_);
  or _69771_ (_18460_, _18458_, _03769_);
  nor _69772_ (_18461_, _18460_, _18455_);
  nor _69773_ (_18462_, _18461_, _18389_);
  nor _69774_ (_18463_, _18462_, _04504_);
  not _69775_ (_18464_, _18386_);
  and _69776_ (_18465_, _18464_, _05376_);
  or _69777_ (_18466_, _18452_, _04505_);
  nor _69778_ (_18467_, _18466_, _18465_);
  nor _69779_ (_18468_, _18467_, _18463_);
  nor _69780_ (_18469_, _18468_, _03752_);
  or _69781_ (_18471_, _18465_, _03753_);
  or _69782_ (_18472_, _18471_, _18395_);
  and _69783_ (_18473_, _18472_, _03759_);
  not _69784_ (_18474_, _18473_);
  nor _69785_ (_18475_, _18474_, _18469_);
  nor _69786_ (_18476_, _13251_, _08818_);
  or _69787_ (_18477_, _18386_, _03759_);
  nor _69788_ (_18478_, _18477_, _18476_);
  or _69789_ (_18479_, _18478_, _03760_);
  nor _69790_ (_18480_, _18479_, _18475_);
  nor _69791_ (_18482_, _13258_, _08818_);
  nor _69792_ (_18483_, _18482_, _18386_);
  nor _69793_ (_18484_, _18483_, _04517_);
  or _69794_ (_18485_, _18484_, _18480_);
  and _69795_ (_18486_, _18485_, _04192_);
  nor _69796_ (_18487_, _18401_, _04192_);
  or _69797_ (_18488_, _18487_, _18486_);
  and _69798_ (_18489_, _18488_, _03152_);
  nor _69799_ (_18490_, _18420_, _03152_);
  or _69800_ (_18491_, _18490_, _18489_);
  and _69801_ (_18493_, _18491_, _03521_);
  and _69802_ (_18494_, _13312_, _05248_);
  nor _69803_ (_18495_, _18494_, _18386_);
  nor _69804_ (_18496_, _18495_, _03521_);
  or _69805_ (_18497_, _18496_, _18493_);
  or _69806_ (_18498_, _18497_, _42967_);
  or _69807_ (_18499_, _42963_, \oc8051_golden_model_1.SCON [6]);
  and _69808_ (_18500_, _18499_, _41755_);
  and _69809_ (_43227_, _18500_, _18498_);
  not _69810_ (_18501_, \oc8051_golden_model_1.PCON [0]);
  nor _69811_ (_18503_, _05208_, _18501_);
  nor _69812_ (_18504_, _05617_, _08940_);
  nor _69813_ (_18505_, _18504_, _18503_);
  and _69814_ (_18506_, _18505_, _17076_);
  and _69815_ (_18507_, _05208_, \oc8051_golden_model_1.ACC [0]);
  nor _69816_ (_18508_, _18507_, _18503_);
  nor _69817_ (_18509_, _18508_, _03583_);
  nor _69818_ (_18510_, _18509_, _07314_);
  nor _69819_ (_18511_, _18505_, _04444_);
  nor _69820_ (_18512_, _04426_, _18501_);
  nor _69821_ (_18514_, _18508_, _04427_);
  nor _69822_ (_18515_, _18514_, _18512_);
  nor _69823_ (_18516_, _18515_, _03570_);
  or _69824_ (_18517_, _18516_, _03568_);
  nor _69825_ (_18518_, _18517_, _18511_);
  or _69826_ (_18519_, _18518_, _03575_);
  and _69827_ (_18520_, _18519_, _18510_);
  and _69828_ (_18521_, _05208_, _04419_);
  and _69829_ (_18522_, _06039_, _03983_);
  or _69830_ (_18523_, _18522_, _18503_);
  nor _69831_ (_18525_, _18523_, _18521_);
  nor _69832_ (_18526_, _18525_, _18520_);
  nor _69833_ (_18527_, _18526_, _03479_);
  and _69834_ (_18528_, _06715_, _05208_);
  nor _69835_ (_18529_, _18503_, _06044_);
  not _69836_ (_18530_, _18529_);
  nor _69837_ (_18531_, _18530_, _18528_);
  nor _69838_ (_18532_, _18531_, _18527_);
  nor _69839_ (_18533_, _18532_, _03221_);
  nor _69840_ (_18534_, _11975_, _08940_);
  or _69841_ (_18536_, _18503_, _03474_);
  nor _69842_ (_18537_, _18536_, _18534_);
  or _69843_ (_18538_, _18537_, _03437_);
  nor _69844_ (_18539_, _18538_, _18533_);
  and _69845_ (_18540_, _05208_, _06202_);
  nor _69846_ (_18541_, _18540_, _18503_);
  nor _69847_ (_18542_, _18541_, _03438_);
  or _69848_ (_18543_, _18542_, _18539_);
  and _69849_ (_18544_, _18543_, _04499_);
  and _69850_ (_18545_, _11990_, _05208_);
  nor _69851_ (_18547_, _18545_, _18503_);
  nor _69852_ (_18548_, _18547_, _04499_);
  or _69853_ (_18549_, _18548_, _18544_);
  nor _69854_ (_18550_, _18549_, _03769_);
  and _69855_ (_18551_, _11995_, _05208_);
  or _69856_ (_18552_, _18503_, _04501_);
  nor _69857_ (_18553_, _18552_, _18551_);
  or _69858_ (_18554_, _18553_, _04504_);
  nor _69859_ (_18555_, _18554_, _18550_);
  or _69860_ (_18556_, _18541_, _04505_);
  nor _69861_ (_18558_, _18556_, _18504_);
  nor _69862_ (_18559_, _18558_, _18555_);
  nor _69863_ (_18560_, _18559_, _03752_);
  and _69864_ (_18561_, _11994_, _05208_);
  or _69865_ (_18562_, _18561_, _18503_);
  and _69866_ (_18563_, _18562_, _03752_);
  or _69867_ (_18564_, _18563_, _18560_);
  and _69868_ (_18565_, _18564_, _03759_);
  nor _69869_ (_18566_, _11988_, _08940_);
  nor _69870_ (_18567_, _18566_, _18503_);
  nor _69871_ (_18569_, _18567_, _03759_);
  or _69872_ (_18570_, _18569_, _18565_);
  and _69873_ (_18571_, _18570_, _04517_);
  nor _69874_ (_18572_, _11870_, _08940_);
  nor _69875_ (_18573_, _18572_, _18503_);
  nor _69876_ (_18574_, _18573_, _04517_);
  nor _69877_ (_18575_, _18574_, _17076_);
  not _69878_ (_18576_, _18575_);
  nor _69879_ (_18577_, _18576_, _18571_);
  nor _69880_ (_18578_, _18577_, _18506_);
  or _69881_ (_18580_, _18578_, _42967_);
  or _69882_ (_18581_, _42963_, \oc8051_golden_model_1.PCON [0]);
  and _69883_ (_18582_, _18581_, _41755_);
  and _69884_ (_43228_, _18582_, _18580_);
  nor _69885_ (_18583_, _05208_, \oc8051_golden_model_1.PCON [1]);
  and _69886_ (_18584_, _12252_, _05208_);
  nor _69887_ (_18585_, _18584_, _18583_);
  nor _69888_ (_18586_, _18585_, _04192_);
  and _69889_ (_18587_, _06714_, _05208_);
  not _69890_ (_18588_, \oc8051_golden_model_1.PCON [1]);
  nor _69891_ (_18590_, _05208_, _18588_);
  nor _69892_ (_18591_, _18590_, _06044_);
  not _69893_ (_18592_, _18591_);
  nor _69894_ (_18593_, _18592_, _18587_);
  not _69895_ (_18594_, _18593_);
  nor _69896_ (_18595_, _08940_, _04603_);
  nor _69897_ (_18596_, _18595_, _18590_);
  and _69898_ (_18597_, _18596_, _07314_);
  and _69899_ (_18598_, _05208_, _03233_);
  nor _69900_ (_18599_, _18598_, _18583_);
  and _69901_ (_18601_, _18599_, _03575_);
  nor _69902_ (_18602_, _18596_, _03983_);
  and _69903_ (_18603_, _18599_, _04426_);
  nor _69904_ (_18604_, _04426_, _18588_);
  or _69905_ (_18605_, _18604_, _18603_);
  and _69906_ (_18606_, _18605_, _04444_);
  and _69907_ (_18607_, _18585_, _03570_);
  or _69908_ (_18608_, _18607_, _18606_);
  and _69909_ (_18609_, _18608_, _03983_);
  nor _69910_ (_18610_, _18609_, _18602_);
  nor _69911_ (_18612_, _18610_, _03575_);
  or _69912_ (_18613_, _18612_, _07314_);
  nor _69913_ (_18614_, _18613_, _18601_);
  nor _69914_ (_18615_, _18614_, _18597_);
  nor _69915_ (_18616_, _18615_, _03479_);
  nor _69916_ (_18617_, _18616_, _03221_);
  and _69917_ (_18618_, _18617_, _18594_);
  not _69918_ (_18619_, _18583_);
  and _69919_ (_18620_, _12176_, _05208_);
  nor _69920_ (_18621_, _18620_, _03474_);
  and _69921_ (_18623_, _18621_, _18619_);
  nor _69922_ (_18624_, _18623_, _18618_);
  nor _69923_ (_18625_, _18624_, _03437_);
  and _69924_ (_18626_, _05208_, _04317_);
  not _69925_ (_18627_, _18626_);
  nor _69926_ (_18628_, _18583_, _03438_);
  and _69927_ (_18629_, _18628_, _18627_);
  nor _69928_ (_18630_, _18629_, _18625_);
  nor _69929_ (_18631_, _18630_, _03636_);
  nor _69930_ (_18632_, _12191_, _08940_);
  nor _69931_ (_18634_, _18632_, _04499_);
  and _69932_ (_18635_, _18634_, _18619_);
  nor _69933_ (_18636_, _18635_, _18631_);
  nor _69934_ (_18637_, _18636_, _03769_);
  nor _69935_ (_18638_, _12197_, _08940_);
  nor _69936_ (_18639_, _18638_, _04501_);
  and _69937_ (_18640_, _18639_, _18619_);
  nor _69938_ (_18641_, _18640_, _18637_);
  nor _69939_ (_18642_, _18641_, _04504_);
  nor _69940_ (_18643_, _12190_, _08940_);
  nor _69941_ (_18645_, _18643_, _05769_);
  and _69942_ (_18646_, _18645_, _18619_);
  nor _69943_ (_18647_, _18646_, _18642_);
  nor _69944_ (_18648_, _18647_, _03752_);
  nor _69945_ (_18649_, _18590_, _05569_);
  nor _69946_ (_18650_, _18649_, _03753_);
  and _69947_ (_18651_, _18650_, _18599_);
  nor _69948_ (_18652_, _18651_, _18648_);
  nor _69949_ (_18653_, _18652_, _03758_);
  and _69950_ (_18654_, _18626_, _05940_);
  nor _69951_ (_18656_, _18654_, _03759_);
  and _69952_ (_18657_, _18656_, _18619_);
  nor _69953_ (_18658_, _18657_, _18653_);
  nor _69954_ (_18659_, _18658_, _03760_);
  nand _69955_ (_18660_, _18598_, _05940_);
  nor _69956_ (_18661_, _18583_, _04517_);
  and _69957_ (_18662_, _18661_, _18660_);
  or _69958_ (_18663_, _18662_, _03790_);
  nor _69959_ (_18664_, _18663_, _18659_);
  nor _69960_ (_18665_, _18664_, _18586_);
  and _69961_ (_18667_, _18665_, _03521_);
  nor _69962_ (_18668_, _18590_, _18584_);
  nor _69963_ (_18669_, _18668_, _03521_);
  or _69964_ (_18670_, _18669_, _18667_);
  or _69965_ (_18671_, _18670_, _42967_);
  or _69966_ (_18672_, _42963_, \oc8051_golden_model_1.PCON [1]);
  and _69967_ (_18673_, _18672_, _41755_);
  and _69968_ (_43229_, _18673_, _18671_);
  not _69969_ (_18674_, \oc8051_golden_model_1.PCON [2]);
  nor _69970_ (_18675_, _05208_, _18674_);
  nor _69971_ (_18677_, _12400_, _08940_);
  nor _69972_ (_18678_, _18677_, _18675_);
  nor _69973_ (_18679_, _18678_, _04517_);
  nor _69974_ (_18680_, _08940_, _05026_);
  nor _69975_ (_18681_, _18680_, _18675_);
  and _69976_ (_18682_, _18681_, _07314_);
  and _69977_ (_18683_, _05208_, \oc8051_golden_model_1.ACC [2]);
  nor _69978_ (_18684_, _18683_, _18675_);
  nor _69979_ (_18685_, _18684_, _04427_);
  nor _69980_ (_18686_, _04426_, _18674_);
  or _69981_ (_18688_, _18686_, _18685_);
  and _69982_ (_18689_, _18688_, _04444_);
  nor _69983_ (_18690_, _12282_, _08940_);
  nor _69984_ (_18691_, _18690_, _18675_);
  nor _69985_ (_18692_, _18691_, _04444_);
  or _69986_ (_18693_, _18692_, _18689_);
  and _69987_ (_18694_, _18693_, _03983_);
  nor _69988_ (_18695_, _18681_, _03983_);
  nor _69989_ (_18696_, _18695_, _18694_);
  nor _69990_ (_18697_, _18696_, _03575_);
  nor _69991_ (_18699_, _18684_, _03583_);
  nor _69992_ (_18700_, _18699_, _07314_);
  not _69993_ (_18701_, _18700_);
  nor _69994_ (_18702_, _18701_, _18697_);
  nor _69995_ (_18703_, _18702_, _18682_);
  nor _69996_ (_18704_, _18703_, _03479_);
  and _69997_ (_18705_, _06718_, _05208_);
  nor _69998_ (_18706_, _18675_, _06044_);
  not _69999_ (_18707_, _18706_);
  nor _70000_ (_18708_, _18707_, _18705_);
  nor _70001_ (_18710_, _18708_, _18704_);
  nor _70002_ (_18711_, _18710_, _03221_);
  nor _70003_ (_18712_, _12384_, _08940_);
  or _70004_ (_18713_, _18675_, _03474_);
  nor _70005_ (_18714_, _18713_, _18712_);
  or _70006_ (_18715_, _18714_, _03437_);
  nor _70007_ (_18716_, _18715_, _18711_);
  and _70008_ (_18717_, _05208_, _06261_);
  nor _70009_ (_18718_, _18717_, _18675_);
  nor _70010_ (_18719_, _18718_, _03438_);
  or _70011_ (_18721_, _18719_, _18716_);
  and _70012_ (_18722_, _18721_, _04499_);
  and _70013_ (_18723_, _12273_, _05208_);
  nor _70014_ (_18724_, _18723_, _18675_);
  nor _70015_ (_18725_, _18724_, _04499_);
  or _70016_ (_18726_, _18725_, _18722_);
  nor _70017_ (_18727_, _18726_, _03769_);
  and _70018_ (_18728_, _12401_, _05208_);
  or _70019_ (_18729_, _18675_, _04501_);
  nor _70020_ (_18730_, _18729_, _18728_);
  or _70021_ (_18732_, _18730_, _04504_);
  nor _70022_ (_18733_, _18732_, _18727_);
  nor _70023_ (_18734_, _18675_, _05665_);
  or _70024_ (_18735_, _18718_, _04505_);
  nor _70025_ (_18736_, _18735_, _18734_);
  nor _70026_ (_18737_, _18736_, _18733_);
  nor _70027_ (_18738_, _18737_, _03752_);
  or _70028_ (_18739_, _18734_, _03753_);
  or _70029_ (_18740_, _18739_, _18684_);
  and _70030_ (_18741_, _18740_, _03759_);
  not _70031_ (_18743_, _18741_);
  nor _70032_ (_18744_, _18743_, _18738_);
  nor _70033_ (_18745_, _12272_, _08940_);
  or _70034_ (_18746_, _18675_, _03759_);
  nor _70035_ (_18747_, _18746_, _18745_);
  or _70036_ (_18748_, _18747_, _03760_);
  nor _70037_ (_18749_, _18748_, _18744_);
  nor _70038_ (_18750_, _18749_, _18679_);
  nor _70039_ (_18751_, _18750_, _03790_);
  nor _70040_ (_18752_, _18691_, _04192_);
  or _70041_ (_18754_, _18752_, _03520_);
  nor _70042_ (_18755_, _18754_, _18751_);
  and _70043_ (_18756_, _12456_, _05208_);
  or _70044_ (_18757_, _18675_, _03521_);
  nor _70045_ (_18758_, _18757_, _18756_);
  nor _70046_ (_18759_, _18758_, _18755_);
  or _70047_ (_18760_, _18759_, _42967_);
  or _70048_ (_18761_, _42963_, \oc8051_golden_model_1.PCON [2]);
  and _70049_ (_18762_, _18761_, _41755_);
  and _70050_ (_43230_, _18762_, _18760_);
  not _70051_ (_18764_, \oc8051_golden_model_1.PCON [3]);
  nor _70052_ (_18765_, _05208_, _18764_);
  and _70053_ (_18766_, _12604_, _05208_);
  nor _70054_ (_18767_, _18766_, _18765_);
  nor _70055_ (_18768_, _18767_, _04501_);
  nor _70056_ (_18769_, _08940_, _04843_);
  nor _70057_ (_18770_, _18769_, _18765_);
  and _70058_ (_18771_, _18770_, _07314_);
  and _70059_ (_18772_, _05208_, \oc8051_golden_model_1.ACC [3]);
  nor _70060_ (_18773_, _18772_, _18765_);
  nor _70061_ (_18775_, _18773_, _03583_);
  nor _70062_ (_18776_, _18773_, _04427_);
  nor _70063_ (_18777_, _04426_, _18764_);
  or _70064_ (_18778_, _18777_, _18776_);
  and _70065_ (_18779_, _18778_, _04444_);
  nor _70066_ (_18780_, _12486_, _08940_);
  nor _70067_ (_18781_, _18780_, _18765_);
  nor _70068_ (_18782_, _18781_, _04444_);
  or _70069_ (_18783_, _18782_, _18779_);
  and _70070_ (_18784_, _18783_, _03983_);
  nor _70071_ (_18786_, _18770_, _03983_);
  nor _70072_ (_18787_, _18786_, _18784_);
  nor _70073_ (_18788_, _18787_, _03575_);
  or _70074_ (_18789_, _18788_, _07314_);
  nor _70075_ (_18790_, _18789_, _18775_);
  nor _70076_ (_18791_, _18790_, _18771_);
  nor _70077_ (_18792_, _18791_, _03479_);
  and _70078_ (_18793_, _06717_, _05208_);
  nor _70079_ (_18794_, _18765_, _06044_);
  not _70080_ (_18795_, _18794_);
  nor _70081_ (_18797_, _18795_, _18793_);
  or _70082_ (_18798_, _18797_, _03221_);
  nor _70083_ (_18799_, _18798_, _18792_);
  nor _70084_ (_18800_, _12583_, _08940_);
  nor _70085_ (_18801_, _18800_, _18765_);
  nor _70086_ (_18802_, _18801_, _03474_);
  or _70087_ (_18803_, _18802_, _03437_);
  or _70088_ (_18804_, _18803_, _18799_);
  and _70089_ (_18805_, _05208_, _06217_);
  nor _70090_ (_18806_, _18805_, _18765_);
  nand _70091_ (_18808_, _18806_, _03437_);
  and _70092_ (_18809_, _18808_, _18804_);
  nor _70093_ (_18810_, _18809_, _03636_);
  and _70094_ (_18811_, _12598_, _05208_);
  or _70095_ (_18812_, _18765_, _04499_);
  nor _70096_ (_18813_, _18812_, _18811_);
  or _70097_ (_18814_, _18813_, _03769_);
  nor _70098_ (_18815_, _18814_, _18810_);
  nor _70099_ (_18816_, _18815_, _18768_);
  nor _70100_ (_18817_, _18816_, _04504_);
  not _70101_ (_18819_, _18765_);
  and _70102_ (_18820_, _18819_, _05520_);
  or _70103_ (_18821_, _18806_, _04505_);
  nor _70104_ (_18822_, _18821_, _18820_);
  nor _70105_ (_18823_, _18822_, _18817_);
  nor _70106_ (_18824_, _18823_, _03752_);
  or _70107_ (_18825_, _18820_, _03753_);
  nor _70108_ (_18826_, _18825_, _18773_);
  or _70109_ (_18827_, _18826_, _18824_);
  and _70110_ (_18828_, _18827_, _03759_);
  nor _70111_ (_18830_, _12597_, _08940_);
  nor _70112_ (_18831_, _18830_, _18765_);
  nor _70113_ (_18832_, _18831_, _03759_);
  or _70114_ (_18833_, _18832_, _18828_);
  and _70115_ (_18834_, _18833_, _04517_);
  nor _70116_ (_18835_, _12603_, _08940_);
  nor _70117_ (_18836_, _18835_, _18765_);
  nor _70118_ (_18837_, _18836_, _04517_);
  or _70119_ (_18838_, _18837_, _03790_);
  nor _70120_ (_18839_, _18838_, _18834_);
  and _70121_ (_18841_, _18781_, _03790_);
  or _70122_ (_18842_, _18841_, _03520_);
  nor _70123_ (_18843_, _18842_, _18839_);
  and _70124_ (_18844_, _12658_, _05208_);
  nor _70125_ (_18845_, _18844_, _18765_);
  nor _70126_ (_18846_, _18845_, _03521_);
  or _70127_ (_18847_, _18846_, _18843_);
  or _70128_ (_18848_, _18847_, _42967_);
  or _70129_ (_18849_, _42963_, \oc8051_golden_model_1.PCON [3]);
  and _70130_ (_18850_, _18849_, _41755_);
  and _70131_ (_43231_, _18850_, _18848_);
  not _70132_ (_18852_, \oc8051_golden_model_1.PCON [4]);
  nor _70133_ (_18853_, _05208_, _18852_);
  and _70134_ (_18854_, _12844_, _05208_);
  nor _70135_ (_18855_, _18854_, _18853_);
  nor _70136_ (_18856_, _18855_, _04501_);
  and _70137_ (_18857_, _05208_, \oc8051_golden_model_1.ACC [4]);
  nor _70138_ (_18858_, _18857_, _18853_);
  nor _70139_ (_18859_, _18858_, _03583_);
  nor _70140_ (_18860_, _18858_, _04427_);
  nor _70141_ (_18862_, _04426_, _18852_);
  or _70142_ (_18863_, _18862_, _18860_);
  and _70143_ (_18864_, _18863_, _04444_);
  nor _70144_ (_18865_, _12733_, _08940_);
  nor _70145_ (_18866_, _18865_, _18853_);
  nor _70146_ (_18867_, _18866_, _04444_);
  or _70147_ (_18868_, _18867_, _18864_);
  and _70148_ (_18869_, _18868_, _03983_);
  nor _70149_ (_18870_, _05712_, _08940_);
  nor _70150_ (_18871_, _18870_, _18853_);
  nor _70151_ (_18873_, _18871_, _03983_);
  nor _70152_ (_18874_, _18873_, _18869_);
  nor _70153_ (_18875_, _18874_, _03575_);
  or _70154_ (_18876_, _18875_, _07314_);
  nor _70155_ (_18877_, _18876_, _18859_);
  and _70156_ (_18878_, _18871_, _07314_);
  or _70157_ (_18879_, _18878_, _03479_);
  nor _70158_ (_18880_, _18879_, _18877_);
  and _70159_ (_18881_, _06722_, _05208_);
  or _70160_ (_18882_, _18881_, _18853_);
  and _70161_ (_18884_, _18882_, _03479_);
  or _70162_ (_18885_, _18884_, _03221_);
  or _70163_ (_18886_, _18885_, _18880_);
  nor _70164_ (_18887_, _12827_, _08940_);
  or _70165_ (_18888_, _18853_, _03474_);
  or _70166_ (_18889_, _18888_, _18887_);
  and _70167_ (_18890_, _18889_, _03438_);
  and _70168_ (_18891_, _18890_, _18886_);
  and _70169_ (_18892_, _06233_, _05208_);
  nor _70170_ (_18893_, _18892_, _18853_);
  nor _70171_ (_18895_, _18893_, _03438_);
  or _70172_ (_18896_, _18895_, _03636_);
  nor _70173_ (_18897_, _18896_, _18891_);
  and _70174_ (_18898_, _12711_, _05208_);
  or _70175_ (_18899_, _18853_, _04499_);
  nor _70176_ (_18900_, _18899_, _18898_);
  or _70177_ (_18901_, _18900_, _03769_);
  nor _70178_ (_18902_, _18901_, _18897_);
  nor _70179_ (_18903_, _18902_, _18856_);
  nor _70180_ (_18904_, _18903_, _04504_);
  not _70181_ (_18906_, _18853_);
  and _70182_ (_18907_, _18906_, _05760_);
  or _70183_ (_18908_, _18893_, _04505_);
  nor _70184_ (_18909_, _18908_, _18907_);
  nor _70185_ (_18910_, _18909_, _18904_);
  nor _70186_ (_18911_, _18910_, _03752_);
  or _70187_ (_18912_, _18907_, _03753_);
  nor _70188_ (_18913_, _18912_, _18858_);
  or _70189_ (_18914_, _18913_, _18911_);
  and _70190_ (_18915_, _18914_, _03759_);
  nor _70191_ (_18917_, _12710_, _08940_);
  nor _70192_ (_18918_, _18917_, _18853_);
  nor _70193_ (_18919_, _18918_, _03759_);
  or _70194_ (_18920_, _18919_, _18915_);
  and _70195_ (_18921_, _18920_, _04517_);
  nor _70196_ (_18922_, _12843_, _08940_);
  nor _70197_ (_18923_, _18922_, _18853_);
  nor _70198_ (_18924_, _18923_, _04517_);
  or _70199_ (_18925_, _18924_, _03790_);
  nor _70200_ (_18926_, _18925_, _18921_);
  and _70201_ (_18928_, _18866_, _03790_);
  or _70202_ (_18929_, _18928_, _03520_);
  nor _70203_ (_18930_, _18929_, _18926_);
  and _70204_ (_18931_, _12893_, _05208_);
  nor _70205_ (_18932_, _18931_, _18853_);
  nor _70206_ (_18933_, _18932_, _03521_);
  or _70207_ (_18934_, _18933_, _18930_);
  or _70208_ (_18935_, _18934_, _42967_);
  or _70209_ (_18936_, _42963_, \oc8051_golden_model_1.PCON [4]);
  and _70210_ (_18937_, _18936_, _41755_);
  and _70211_ (_43232_, _18937_, _18935_);
  not _70212_ (_18939_, \oc8051_golden_model_1.PCON [5]);
  nor _70213_ (_18940_, _05208_, _18939_);
  and _70214_ (_18941_, _13042_, _05208_);
  nor _70215_ (_18942_, _18941_, _18940_);
  nor _70216_ (_18943_, _18942_, _04501_);
  and _70217_ (_18944_, _05208_, \oc8051_golden_model_1.ACC [5]);
  nor _70218_ (_18945_, _18944_, _18940_);
  nor _70219_ (_18946_, _18945_, _03583_);
  nor _70220_ (_18947_, _18945_, _04427_);
  nor _70221_ (_18949_, _04426_, _18939_);
  or _70222_ (_18950_, _18949_, _18947_);
  and _70223_ (_18951_, _18950_, _04444_);
  nor _70224_ (_18952_, _12930_, _08940_);
  nor _70225_ (_18953_, _18952_, _18940_);
  nor _70226_ (_18954_, _18953_, _04444_);
  or _70227_ (_18955_, _18954_, _18951_);
  and _70228_ (_18956_, _18955_, _03983_);
  nor _70229_ (_18957_, _05422_, _08940_);
  nor _70230_ (_18958_, _18957_, _18940_);
  nor _70231_ (_18960_, _18958_, _03983_);
  nor _70232_ (_18961_, _18960_, _18956_);
  nor _70233_ (_18962_, _18961_, _03575_);
  or _70234_ (_18963_, _18962_, _07314_);
  nor _70235_ (_18964_, _18963_, _18946_);
  and _70236_ (_18965_, _18958_, _07314_);
  nor _70237_ (_18966_, _18965_, _18964_);
  nor _70238_ (_18967_, _18966_, _03479_);
  and _70239_ (_18968_, _06721_, _05208_);
  nor _70240_ (_18969_, _18940_, _06044_);
  not _70241_ (_18971_, _18969_);
  nor _70242_ (_18972_, _18971_, _18968_);
  or _70243_ (_18973_, _18972_, _03221_);
  nor _70244_ (_18974_, _18973_, _18967_);
  nor _70245_ (_18975_, _13021_, _08940_);
  nor _70246_ (_18976_, _18975_, _18940_);
  nor _70247_ (_18977_, _18976_, _03474_);
  or _70248_ (_18978_, _18977_, _03437_);
  or _70249_ (_18979_, _18978_, _18974_);
  and _70250_ (_18980_, _06211_, _05208_);
  nor _70251_ (_18982_, _18980_, _18940_);
  nand _70252_ (_18983_, _18982_, _03437_);
  and _70253_ (_18984_, _18983_, _18979_);
  nor _70254_ (_18985_, _18984_, _03636_);
  and _70255_ (_18986_, _13036_, _05208_);
  or _70256_ (_18987_, _18940_, _04499_);
  nor _70257_ (_18988_, _18987_, _18986_);
  or _70258_ (_18989_, _18988_, _03769_);
  nor _70259_ (_18990_, _18989_, _18985_);
  nor _70260_ (_18991_, _18990_, _18943_);
  nor _70261_ (_18993_, _18991_, _04504_);
  not _70262_ (_18994_, _18940_);
  and _70263_ (_18995_, _18994_, _05471_);
  or _70264_ (_18996_, _18982_, _04505_);
  nor _70265_ (_18997_, _18996_, _18995_);
  nor _70266_ (_18998_, _18997_, _18993_);
  nor _70267_ (_18999_, _18998_, _03752_);
  or _70268_ (_19000_, _18995_, _03753_);
  or _70269_ (_19001_, _19000_, _18945_);
  and _70270_ (_19002_, _19001_, _03759_);
  not _70271_ (_19004_, _19002_);
  nor _70272_ (_19005_, _19004_, _18999_);
  nor _70273_ (_19006_, _13035_, _08940_);
  or _70274_ (_19007_, _18940_, _03759_);
  nor _70275_ (_19008_, _19007_, _19006_);
  or _70276_ (_19009_, _19008_, _03760_);
  nor _70277_ (_19010_, _19009_, _19005_);
  nor _70278_ (_19011_, _13041_, _08940_);
  nor _70279_ (_19012_, _19011_, _18940_);
  nor _70280_ (_19013_, _19012_, _04517_);
  or _70281_ (_19015_, _19013_, _03790_);
  nor _70282_ (_19016_, _19015_, _19010_);
  and _70283_ (_19017_, _18953_, _03790_);
  or _70284_ (_19018_, _19017_, _03520_);
  nor _70285_ (_19019_, _19018_, _19016_);
  and _70286_ (_19020_, _13097_, _05208_);
  nor _70287_ (_19021_, _19020_, _18940_);
  nor _70288_ (_19022_, _19021_, _03521_);
  or _70289_ (_19023_, _19022_, _19019_);
  or _70290_ (_19024_, _19023_, _42967_);
  or _70291_ (_19026_, _42963_, \oc8051_golden_model_1.PCON [5]);
  and _70292_ (_19027_, _19026_, _41755_);
  and _70293_ (_43233_, _19027_, _19024_);
  not _70294_ (_19028_, \oc8051_golden_model_1.PCON [6]);
  nor _70295_ (_19029_, _05208_, _19028_);
  and _70296_ (_19030_, _13259_, _05208_);
  nor _70297_ (_19031_, _19030_, _19029_);
  nor _70298_ (_19032_, _19031_, _04501_);
  nor _70299_ (_19033_, _05327_, _08940_);
  nor _70300_ (_19034_, _19033_, _19029_);
  and _70301_ (_19036_, _19034_, _07314_);
  and _70302_ (_19037_, _05208_, \oc8051_golden_model_1.ACC [6]);
  nor _70303_ (_19038_, _19037_, _19029_);
  nor _70304_ (_19039_, _19038_, _04427_);
  nor _70305_ (_19040_, _04426_, _19028_);
  or _70306_ (_19041_, _19040_, _19039_);
  and _70307_ (_19042_, _19041_, _04444_);
  nor _70308_ (_19043_, _13122_, _08940_);
  nor _70309_ (_19044_, _19043_, _19029_);
  nor _70310_ (_19045_, _19044_, _04444_);
  or _70311_ (_19047_, _19045_, _19042_);
  and _70312_ (_19048_, _19047_, _03983_);
  nor _70313_ (_19049_, _19034_, _03983_);
  nor _70314_ (_19050_, _19049_, _19048_);
  nor _70315_ (_19051_, _19050_, _03575_);
  nor _70316_ (_19052_, _19038_, _03583_);
  nor _70317_ (_19053_, _19052_, _07314_);
  not _70318_ (_19054_, _19053_);
  nor _70319_ (_19055_, _19054_, _19051_);
  nor _70320_ (_19056_, _19055_, _19036_);
  nor _70321_ (_19058_, _19056_, _03479_);
  and _70322_ (_19059_, _06713_, _05208_);
  nor _70323_ (_19060_, _19029_, _06044_);
  not _70324_ (_19061_, _19060_);
  nor _70325_ (_19062_, _19061_, _19059_);
  or _70326_ (_19063_, _19062_, _03221_);
  nor _70327_ (_19064_, _19063_, _19058_);
  nor _70328_ (_19065_, _13237_, _08940_);
  nor _70329_ (_19066_, _19065_, _19029_);
  nor _70330_ (_19067_, _19066_, _03474_);
  or _70331_ (_19069_, _19067_, _03437_);
  or _70332_ (_19070_, _19069_, _19064_);
  and _70333_ (_19071_, _13244_, _05208_);
  nor _70334_ (_19072_, _19071_, _19029_);
  nand _70335_ (_19073_, _19072_, _03437_);
  and _70336_ (_19074_, _19073_, _19070_);
  nor _70337_ (_19075_, _19074_, _03636_);
  and _70338_ (_19076_, _13253_, _05208_);
  or _70339_ (_19077_, _19029_, _04499_);
  nor _70340_ (_19078_, _19077_, _19076_);
  or _70341_ (_19080_, _19078_, _03769_);
  nor _70342_ (_19081_, _19080_, _19075_);
  nor _70343_ (_19082_, _19081_, _19032_);
  nor _70344_ (_19083_, _19082_, _04504_);
  not _70345_ (_19084_, _19029_);
  and _70346_ (_19085_, _19084_, _05376_);
  or _70347_ (_19086_, _19072_, _04505_);
  nor _70348_ (_19087_, _19086_, _19085_);
  nor _70349_ (_19088_, _19087_, _19083_);
  nor _70350_ (_19089_, _19088_, _03752_);
  or _70351_ (_19091_, _19085_, _03753_);
  nor _70352_ (_19092_, _19091_, _19038_);
  or _70353_ (_19093_, _19092_, _19089_);
  and _70354_ (_19094_, _19093_, _03759_);
  nor _70355_ (_19095_, _13251_, _08940_);
  nor _70356_ (_19096_, _19095_, _19029_);
  nor _70357_ (_19097_, _19096_, _03759_);
  or _70358_ (_19098_, _19097_, _19094_);
  and _70359_ (_19099_, _19098_, _04517_);
  nor _70360_ (_19100_, _13258_, _08940_);
  nor _70361_ (_19102_, _19100_, _19029_);
  nor _70362_ (_19103_, _19102_, _04517_);
  or _70363_ (_19104_, _19103_, _03790_);
  nor _70364_ (_19105_, _19104_, _19099_);
  and _70365_ (_19106_, _19044_, _03790_);
  or _70366_ (_19107_, _19106_, _03520_);
  nor _70367_ (_19108_, _19107_, _19105_);
  and _70368_ (_19109_, _13312_, _05208_);
  nor _70369_ (_19110_, _19109_, _19029_);
  nor _70370_ (_19111_, _19110_, _03521_);
  or _70371_ (_19113_, _19111_, _19108_);
  or _70372_ (_19114_, _19113_, _42967_);
  or _70373_ (_19115_, _42963_, \oc8051_golden_model_1.PCON [6]);
  and _70374_ (_19116_, _19115_, _41755_);
  and _70375_ (_43234_, _19116_, _19114_);
  not _70376_ (_19117_, \oc8051_golden_model_1.TCON [0]);
  nor _70377_ (_19118_, _05236_, _19117_);
  and _70378_ (_19119_, _11995_, _05236_);
  nor _70379_ (_19120_, _19119_, _19118_);
  nor _70380_ (_19121_, _19120_, _04501_);
  and _70381_ (_19123_, _05236_, _04419_);
  nor _70382_ (_19124_, _19123_, _19118_);
  and _70383_ (_19125_, _19124_, _07314_);
  and _70384_ (_19126_, _05236_, \oc8051_golden_model_1.ACC [0]);
  nor _70385_ (_19127_, _19126_, _19118_);
  nor _70386_ (_19128_, _19127_, _04427_);
  nor _70387_ (_19129_, _04426_, _19117_);
  or _70388_ (_19130_, _19129_, _19128_);
  and _70389_ (_19131_, _19130_, _04444_);
  and _70390_ (_19132_, _05941_, _05236_);
  nor _70391_ (_19134_, _19132_, _19118_);
  nor _70392_ (_19135_, _19134_, _04444_);
  or _70393_ (_19136_, _19135_, _19131_);
  and _70394_ (_19137_, _19136_, _03517_);
  nor _70395_ (_19138_, _05799_, _19117_);
  and _70396_ (_19139_, _11887_, _05799_);
  nor _70397_ (_19140_, _19139_, _19138_);
  nor _70398_ (_19141_, _19140_, _03517_);
  nor _70399_ (_19142_, _19141_, _19137_);
  nor _70400_ (_19143_, _19142_, _03568_);
  nor _70401_ (_19145_, _19124_, _03983_);
  or _70402_ (_19146_, _19145_, _19143_);
  and _70403_ (_19147_, _19146_, _03583_);
  nor _70404_ (_19148_, _19127_, _03583_);
  or _70405_ (_19149_, _19148_, _19147_);
  and _70406_ (_19150_, _19149_, _03513_);
  and _70407_ (_19151_, _19118_, _03512_);
  or _70408_ (_19152_, _19151_, _19150_);
  and _70409_ (_19153_, _19152_, _03506_);
  nor _70410_ (_19154_, _19134_, _03506_);
  or _70411_ (_19156_, _19154_, _19153_);
  and _70412_ (_19157_, _19156_, _03500_);
  nor _70413_ (_19158_, _11916_, _09052_);
  nor _70414_ (_19159_, _19158_, _19138_);
  nor _70415_ (_19160_, _19159_, _03500_);
  or _70416_ (_19161_, _19160_, _07314_);
  nor _70417_ (_19162_, _19161_, _19157_);
  nor _70418_ (_19163_, _19162_, _19125_);
  nor _70419_ (_19164_, _19163_, _03479_);
  and _70420_ (_19165_, _06715_, _05236_);
  nor _70421_ (_19167_, _19118_, _06044_);
  not _70422_ (_19168_, _19167_);
  nor _70423_ (_19169_, _19168_, _19165_);
  or _70424_ (_19170_, _19169_, _03221_);
  nor _70425_ (_19171_, _19170_, _19164_);
  nor _70426_ (_19172_, _11975_, _09015_);
  nor _70427_ (_19173_, _19172_, _19118_);
  nor _70428_ (_19174_, _19173_, _03474_);
  or _70429_ (_19175_, _19174_, _03437_);
  or _70430_ (_19176_, _19175_, _19171_);
  and _70431_ (_19178_, _05236_, _06202_);
  nor _70432_ (_19179_, _19178_, _19118_);
  nand _70433_ (_19180_, _19179_, _03437_);
  and _70434_ (_19181_, _19180_, _19176_);
  nor _70435_ (_19182_, _19181_, _03636_);
  and _70436_ (_19183_, _11990_, _05236_);
  or _70437_ (_19184_, _19118_, _04499_);
  nor _70438_ (_19185_, _19184_, _19183_);
  or _70439_ (_19186_, _19185_, _03769_);
  nor _70440_ (_19187_, _19186_, _19182_);
  nor _70441_ (_19189_, _19187_, _19121_);
  nor _70442_ (_19190_, _19189_, _04504_);
  or _70443_ (_19191_, _19179_, _04505_);
  nor _70444_ (_19192_, _19191_, _19132_);
  nor _70445_ (_19193_, _19192_, _19190_);
  nor _70446_ (_19194_, _19193_, _03752_);
  and _70447_ (_19195_, _11994_, _05236_);
  or _70448_ (_19196_, _19195_, _19118_);
  and _70449_ (_19197_, _19196_, _03752_);
  or _70450_ (_19198_, _19197_, _19194_);
  and _70451_ (_19200_, _19198_, _03759_);
  nor _70452_ (_19201_, _11988_, _09015_);
  nor _70453_ (_19202_, _19201_, _19118_);
  nor _70454_ (_19203_, _19202_, _03759_);
  or _70455_ (_19204_, _19203_, _19200_);
  and _70456_ (_19205_, _19204_, _04517_);
  nor _70457_ (_19206_, _11870_, _09015_);
  nor _70458_ (_19207_, _19206_, _19118_);
  nor _70459_ (_19208_, _19207_, _04517_);
  or _70460_ (_19209_, _19208_, _19205_);
  and _70461_ (_19211_, _19209_, _04192_);
  nor _70462_ (_19212_, _19134_, _04192_);
  or _70463_ (_19213_, _19212_, _19211_);
  and _70464_ (_19214_, _19213_, _03152_);
  and _70465_ (_19215_, _19118_, _03151_);
  or _70466_ (_19216_, _19215_, _19214_);
  and _70467_ (_19217_, _19216_, _03521_);
  nor _70468_ (_19218_, _19134_, _03521_);
  or _70469_ (_19219_, _19218_, _19217_);
  or _70470_ (_19220_, _19219_, _42967_);
  or _70471_ (_19222_, _42963_, \oc8051_golden_model_1.TCON [0]);
  and _70472_ (_19223_, _19222_, _41755_);
  and _70473_ (_43237_, _19223_, _19220_);
  or _70474_ (_19224_, _05236_, \oc8051_golden_model_1.TCON [1]);
  and _70475_ (_19225_, _12252_, _05236_);
  not _70476_ (_19226_, _19225_);
  and _70477_ (_19227_, _19226_, _19224_);
  or _70478_ (_19228_, _19227_, _04444_);
  nand _70479_ (_19229_, _05236_, _03233_);
  and _70480_ (_19230_, _19229_, _19224_);
  and _70481_ (_19232_, _19230_, _04426_);
  not _70482_ (_19233_, \oc8051_golden_model_1.TCON [1]);
  nor _70483_ (_19234_, _04426_, _19233_);
  or _70484_ (_19235_, _19234_, _03570_);
  or _70485_ (_19236_, _19235_, _19232_);
  and _70486_ (_19237_, _19236_, _03517_);
  and _70487_ (_19238_, _19237_, _19228_);
  and _70488_ (_19239_, _12083_, _05799_);
  nor _70489_ (_19240_, _05799_, _19233_);
  or _70490_ (_19241_, _19240_, _03568_);
  or _70491_ (_19243_, _19241_, _19239_);
  and _70492_ (_19244_, _19243_, _14165_);
  or _70493_ (_19245_, _19244_, _19238_);
  nor _70494_ (_19246_, _05236_, _19233_);
  nor _70495_ (_19247_, _09015_, _04603_);
  or _70496_ (_19248_, _19247_, _19246_);
  or _70497_ (_19249_, _19248_, _03983_);
  and _70498_ (_19250_, _19249_, _19245_);
  or _70499_ (_19251_, _19250_, _03575_);
  or _70500_ (_19252_, _19230_, _03583_);
  and _70501_ (_19254_, _19252_, _03513_);
  and _70502_ (_19255_, _19254_, _19251_);
  and _70503_ (_19256_, _12069_, _05799_);
  or _70504_ (_19257_, _19256_, _19240_);
  and _70505_ (_19258_, _19257_, _03512_);
  or _70506_ (_19259_, _19258_, _03505_);
  or _70507_ (_19260_, _19259_, _19255_);
  and _70508_ (_19261_, _19239_, _12098_);
  or _70509_ (_19262_, _19240_, _03506_);
  or _70510_ (_19263_, _19262_, _19261_);
  and _70511_ (_19265_, _19263_, _19260_);
  and _70512_ (_19266_, _19265_, _03500_);
  nor _70513_ (_19267_, _12116_, _09052_);
  or _70514_ (_19268_, _19240_, _19267_);
  and _70515_ (_19269_, _19268_, _03499_);
  or _70516_ (_19270_, _19269_, _07314_);
  or _70517_ (_19271_, _19270_, _19266_);
  or _70518_ (_19272_, _19248_, _06039_);
  and _70519_ (_19273_, _19272_, _19271_);
  or _70520_ (_19274_, _19273_, _03479_);
  and _70521_ (_19276_, _06714_, _05236_);
  or _70522_ (_19277_, _19246_, _06044_);
  or _70523_ (_19278_, _19277_, _19276_);
  and _70524_ (_19279_, _19278_, _03474_);
  and _70525_ (_19280_, _19279_, _19274_);
  nor _70526_ (_19281_, _12176_, _09015_);
  or _70527_ (_19282_, _19281_, _19246_);
  and _70528_ (_19283_, _19282_, _03221_);
  or _70529_ (_19284_, _19283_, _19280_);
  and _70530_ (_19285_, _19284_, _03438_);
  nand _70531_ (_19287_, _05236_, _04317_);
  and _70532_ (_19288_, _19224_, _03437_);
  and _70533_ (_19289_, _19288_, _19287_);
  or _70534_ (_19290_, _19289_, _19285_);
  and _70535_ (_19291_, _19290_, _04499_);
  or _70536_ (_19292_, _12191_, _09015_);
  and _70537_ (_19293_, _19224_, _03636_);
  and _70538_ (_19294_, _19293_, _19292_);
  or _70539_ (_19295_, _19294_, _19291_);
  and _70540_ (_19296_, _19295_, _04501_);
  or _70541_ (_19298_, _12197_, _09015_);
  and _70542_ (_19299_, _19224_, _03769_);
  and _70543_ (_19300_, _19299_, _19298_);
  or _70544_ (_19301_, _19300_, _19296_);
  and _70545_ (_19302_, _19301_, _05769_);
  or _70546_ (_19303_, _12190_, _09015_);
  and _70547_ (_19304_, _19303_, _03754_);
  and _70548_ (_19305_, _19304_, _19224_);
  or _70549_ (_19306_, _19305_, _19302_);
  and _70550_ (_19307_, _19306_, _03753_);
  or _70551_ (_19309_, _19246_, _05569_);
  and _70552_ (_19310_, _19230_, _03752_);
  and _70553_ (_19311_, _19310_, _19309_);
  or _70554_ (_19312_, _19311_, _19307_);
  and _70555_ (_19313_, _19312_, _03759_);
  or _70556_ (_19314_, _19287_, _05569_);
  and _70557_ (_19315_, _19224_, _03758_);
  and _70558_ (_19316_, _19315_, _19314_);
  or _70559_ (_19317_, _19316_, _19313_);
  and _70560_ (_19318_, _19317_, _04517_);
  or _70561_ (_19320_, _19229_, _05569_);
  and _70562_ (_19321_, _19224_, _03760_);
  and _70563_ (_19322_, _19321_, _19320_);
  or _70564_ (_19323_, _19322_, _03790_);
  or _70565_ (_19324_, _19323_, _19318_);
  or _70566_ (_19325_, _19227_, _04192_);
  and _70567_ (_19326_, _19325_, _03152_);
  and _70568_ (_19327_, _19326_, _19324_);
  and _70569_ (_19328_, _19257_, _03151_);
  or _70570_ (_19329_, _19328_, _03520_);
  or _70571_ (_19331_, _19329_, _19327_);
  or _70572_ (_19332_, _19246_, _03521_);
  or _70573_ (_19333_, _19332_, _19225_);
  and _70574_ (_19334_, _19333_, _19331_);
  and _70575_ (_19335_, _19334_, _42963_);
  nor _70576_ (_19336_, \oc8051_golden_model_1.TCON [1], rst);
  nor _70577_ (_19337_, _19336_, _00000_);
  or _70578_ (_43238_, _19337_, _19335_);
  not _70579_ (_19338_, \oc8051_golden_model_1.TCON [2]);
  nor _70580_ (_19339_, _05236_, _19338_);
  and _70581_ (_19341_, _12401_, _05236_);
  nor _70582_ (_19342_, _19341_, _19339_);
  nor _70583_ (_19343_, _19342_, _04501_);
  nor _70584_ (_19344_, _09015_, _05026_);
  nor _70585_ (_19345_, _19344_, _19339_);
  and _70586_ (_19346_, _19345_, _07314_);
  nor _70587_ (_19347_, _19345_, _03983_);
  nor _70588_ (_19348_, _05799_, _19338_);
  and _70589_ (_19349_, _12278_, _05799_);
  nor _70590_ (_19350_, _19349_, _19348_);
  and _70591_ (_19352_, _19350_, _03516_);
  nor _70592_ (_19353_, _12282_, _09015_);
  nor _70593_ (_19354_, _19353_, _19339_);
  nor _70594_ (_19355_, _19354_, _04444_);
  nor _70595_ (_19356_, _04426_, _19338_);
  and _70596_ (_19357_, _05236_, \oc8051_golden_model_1.ACC [2]);
  nor _70597_ (_19358_, _19357_, _19339_);
  nor _70598_ (_19359_, _19358_, _04427_);
  nor _70599_ (_19360_, _19359_, _19356_);
  nor _70600_ (_19361_, _19360_, _03570_);
  or _70601_ (_19363_, _19361_, _03516_);
  nor _70602_ (_19364_, _19363_, _19355_);
  nor _70603_ (_19365_, _19364_, _19352_);
  and _70604_ (_19366_, _19365_, _03983_);
  or _70605_ (_19367_, _19366_, _19347_);
  and _70606_ (_19368_, _19367_, _03583_);
  nor _70607_ (_19369_, _19358_, _03583_);
  or _70608_ (_19370_, _19369_, _19368_);
  and _70609_ (_19371_, _19370_, _03513_);
  and _70610_ (_19372_, _12276_, _05799_);
  nor _70611_ (_19374_, _19372_, _19348_);
  nor _70612_ (_19375_, _19374_, _03513_);
  or _70613_ (_19376_, _19375_, _03505_);
  or _70614_ (_19377_, _19376_, _19371_);
  nor _70615_ (_19378_, _19348_, _12309_);
  nor _70616_ (_19379_, _19378_, _19350_);
  or _70617_ (_19380_, _19379_, _03506_);
  and _70618_ (_19381_, _19380_, _03500_);
  and _70619_ (_19382_, _19381_, _19377_);
  nor _70620_ (_19383_, _12326_, _09052_);
  nor _70621_ (_19385_, _19383_, _19348_);
  nor _70622_ (_19386_, _19385_, _03500_);
  nor _70623_ (_19387_, _19386_, _07314_);
  not _70624_ (_19388_, _19387_);
  nor _70625_ (_19389_, _19388_, _19382_);
  nor _70626_ (_19390_, _19389_, _19346_);
  nor _70627_ (_19391_, _19390_, _03479_);
  and _70628_ (_19392_, _06718_, _05236_);
  nor _70629_ (_19393_, _19339_, _06044_);
  not _70630_ (_19394_, _19393_);
  nor _70631_ (_19396_, _19394_, _19392_);
  or _70632_ (_19397_, _19396_, _03221_);
  nor _70633_ (_19398_, _19397_, _19391_);
  nor _70634_ (_19399_, _12384_, _09015_);
  nor _70635_ (_19400_, _19399_, _19339_);
  nor _70636_ (_19401_, _19400_, _03474_);
  or _70637_ (_19402_, _19401_, _03437_);
  or _70638_ (_19403_, _19402_, _19398_);
  and _70639_ (_19404_, _05236_, _06261_);
  nor _70640_ (_19405_, _19404_, _19339_);
  nand _70641_ (_19407_, _19405_, _03437_);
  and _70642_ (_19408_, _19407_, _19403_);
  nor _70643_ (_19409_, _19408_, _03636_);
  and _70644_ (_19410_, _12273_, _05236_);
  or _70645_ (_19411_, _19339_, _04499_);
  nor _70646_ (_19412_, _19411_, _19410_);
  or _70647_ (_19413_, _19412_, _03769_);
  nor _70648_ (_19414_, _19413_, _19409_);
  nor _70649_ (_19415_, _19414_, _19343_);
  nor _70650_ (_19416_, _19415_, _04504_);
  not _70651_ (_19418_, _19339_);
  and _70652_ (_19419_, _19418_, _05664_);
  or _70653_ (_19420_, _19405_, _04505_);
  nor _70654_ (_19421_, _19420_, _19419_);
  nor _70655_ (_19422_, _19421_, _19416_);
  nor _70656_ (_19423_, _19422_, _03752_);
  or _70657_ (_19424_, _19419_, _03753_);
  nor _70658_ (_19425_, _19424_, _19358_);
  or _70659_ (_19426_, _19425_, _19423_);
  and _70660_ (_19427_, _19426_, _03759_);
  nor _70661_ (_19429_, _12272_, _09015_);
  nor _70662_ (_19430_, _19429_, _19339_);
  nor _70663_ (_19431_, _19430_, _03759_);
  or _70664_ (_19432_, _19431_, _19427_);
  and _70665_ (_19433_, _19432_, _04517_);
  nor _70666_ (_19434_, _12400_, _09015_);
  nor _70667_ (_19435_, _19434_, _19339_);
  nor _70668_ (_19436_, _19435_, _04517_);
  or _70669_ (_19437_, _19436_, _19433_);
  and _70670_ (_19438_, _19437_, _04192_);
  nor _70671_ (_19440_, _19354_, _04192_);
  or _70672_ (_19441_, _19440_, _19438_);
  and _70673_ (_19442_, _19441_, _03152_);
  nor _70674_ (_19443_, _19374_, _03152_);
  or _70675_ (_19444_, _19443_, _19442_);
  and _70676_ (_19445_, _19444_, _03521_);
  and _70677_ (_19446_, _12456_, _05236_);
  nor _70678_ (_19447_, _19446_, _19339_);
  nor _70679_ (_19448_, _19447_, _03521_);
  or _70680_ (_19449_, _19448_, _19445_);
  or _70681_ (_19451_, _19449_, _42967_);
  or _70682_ (_19452_, _42963_, \oc8051_golden_model_1.TCON [2]);
  and _70683_ (_19453_, _19452_, _41755_);
  and _70684_ (_43239_, _19453_, _19451_);
  not _70685_ (_19454_, \oc8051_golden_model_1.TCON [3]);
  nor _70686_ (_19455_, _05236_, _19454_);
  and _70687_ (_19456_, _12604_, _05236_);
  nor _70688_ (_19457_, _19456_, _19455_);
  nor _70689_ (_19458_, _19457_, _04501_);
  nor _70690_ (_19459_, _09015_, _04843_);
  nor _70691_ (_19461_, _19459_, _19455_);
  and _70692_ (_19462_, _19461_, _07314_);
  and _70693_ (_19463_, _05236_, \oc8051_golden_model_1.ACC [3]);
  nor _70694_ (_19464_, _19463_, _19455_);
  nor _70695_ (_19465_, _19464_, _04427_);
  nor _70696_ (_19466_, _04426_, _19454_);
  or _70697_ (_19467_, _19466_, _19465_);
  and _70698_ (_19468_, _19467_, _04444_);
  nor _70699_ (_19469_, _12486_, _09015_);
  nor _70700_ (_19470_, _19469_, _19455_);
  nor _70701_ (_19472_, _19470_, _04444_);
  or _70702_ (_19473_, _19472_, _19468_);
  and _70703_ (_19474_, _19473_, _03517_);
  nor _70704_ (_19475_, _05799_, _19454_);
  and _70705_ (_19476_, _12490_, _05799_);
  nor _70706_ (_19477_, _19476_, _19475_);
  nor _70707_ (_19478_, _19477_, _03517_);
  or _70708_ (_19479_, _19478_, _03568_);
  or _70709_ (_19480_, _19479_, _19474_);
  nand _70710_ (_19481_, _19461_, _03568_);
  and _70711_ (_19483_, _19481_, _19480_);
  and _70712_ (_19484_, _19483_, _03583_);
  nor _70713_ (_19485_, _19464_, _03583_);
  or _70714_ (_19486_, _19485_, _19484_);
  and _70715_ (_19487_, _19486_, _03513_);
  and _70716_ (_19488_, _12500_, _05799_);
  nor _70717_ (_19489_, _19488_, _19475_);
  nor _70718_ (_19490_, _19489_, _03513_);
  or _70719_ (_19491_, _19490_, _19487_);
  and _70720_ (_19492_, _19491_, _03506_);
  nor _70721_ (_19494_, _19475_, _12507_);
  nor _70722_ (_19495_, _19494_, _19477_);
  and _70723_ (_19496_, _19495_, _03505_);
  or _70724_ (_19497_, _19496_, _19492_);
  and _70725_ (_19498_, _19497_, _03500_);
  nor _70726_ (_19499_, _12525_, _09052_);
  nor _70727_ (_19500_, _19499_, _19475_);
  nor _70728_ (_19501_, _19500_, _03500_);
  nor _70729_ (_19502_, _19501_, _07314_);
  not _70730_ (_19503_, _19502_);
  nor _70731_ (_19505_, _19503_, _19498_);
  nor _70732_ (_19506_, _19505_, _19462_);
  nor _70733_ (_19507_, _19506_, _03479_);
  and _70734_ (_19508_, _06717_, _05236_);
  nor _70735_ (_19509_, _19455_, _06044_);
  not _70736_ (_19510_, _19509_);
  nor _70737_ (_19511_, _19510_, _19508_);
  or _70738_ (_19512_, _19511_, _03221_);
  nor _70739_ (_19513_, _19512_, _19507_);
  nor _70740_ (_19514_, _12583_, _09015_);
  nor _70741_ (_19516_, _19514_, _19455_);
  nor _70742_ (_19517_, _19516_, _03474_);
  or _70743_ (_19518_, _19517_, _03437_);
  or _70744_ (_19519_, _19518_, _19513_);
  and _70745_ (_19520_, _05236_, _06217_);
  nor _70746_ (_19521_, _19520_, _19455_);
  nand _70747_ (_19522_, _19521_, _03437_);
  and _70748_ (_19523_, _19522_, _19519_);
  nor _70749_ (_19524_, _19523_, _03636_);
  and _70750_ (_19525_, _12598_, _05236_);
  or _70751_ (_19527_, _19455_, _04499_);
  nor _70752_ (_19528_, _19527_, _19525_);
  or _70753_ (_19529_, _19528_, _03769_);
  nor _70754_ (_19530_, _19529_, _19524_);
  nor _70755_ (_19531_, _19530_, _19458_);
  nor _70756_ (_19532_, _19531_, _04504_);
  not _70757_ (_19533_, _19455_);
  and _70758_ (_19534_, _19533_, _05520_);
  or _70759_ (_19535_, _19521_, _04505_);
  nor _70760_ (_19536_, _19535_, _19534_);
  nor _70761_ (_19538_, _19536_, _19532_);
  nor _70762_ (_19539_, _19538_, _03752_);
  or _70763_ (_19540_, _19534_, _03753_);
  nor _70764_ (_19541_, _19540_, _19464_);
  or _70765_ (_19542_, _19541_, _19539_);
  and _70766_ (_19543_, _19542_, _03759_);
  nor _70767_ (_19544_, _12597_, _09015_);
  nor _70768_ (_19545_, _19544_, _19455_);
  nor _70769_ (_19546_, _19545_, _03759_);
  or _70770_ (_19547_, _19546_, _19543_);
  and _70771_ (_19549_, _19547_, _04517_);
  nor _70772_ (_19550_, _12603_, _09015_);
  nor _70773_ (_19551_, _19550_, _19455_);
  nor _70774_ (_19552_, _19551_, _04517_);
  or _70775_ (_19553_, _19552_, _19549_);
  and _70776_ (_19554_, _19553_, _04192_);
  nor _70777_ (_19555_, _19470_, _04192_);
  or _70778_ (_19556_, _19555_, _19554_);
  and _70779_ (_19557_, _19556_, _03152_);
  nor _70780_ (_19558_, _19489_, _03152_);
  or _70781_ (_19560_, _19558_, _19557_);
  and _70782_ (_19561_, _19560_, _03521_);
  and _70783_ (_19562_, _12658_, _05236_);
  nor _70784_ (_19563_, _19562_, _19455_);
  nor _70785_ (_19564_, _19563_, _03521_);
  or _70786_ (_19565_, _19564_, _19561_);
  or _70787_ (_19566_, _19565_, _42967_);
  or _70788_ (_19567_, _42963_, \oc8051_golden_model_1.TCON [3]);
  and _70789_ (_19568_, _19567_, _41755_);
  and _70790_ (_43242_, _19568_, _19566_);
  not _70791_ (_19570_, \oc8051_golden_model_1.TCON [4]);
  nor _70792_ (_19571_, _05236_, _19570_);
  and _70793_ (_19572_, _12844_, _05236_);
  nor _70794_ (_19573_, _19572_, _19571_);
  nor _70795_ (_19574_, _19573_, _04501_);
  nor _70796_ (_19575_, _05712_, _09015_);
  nor _70797_ (_19576_, _19575_, _19571_);
  and _70798_ (_19577_, _19576_, _07314_);
  and _70799_ (_19578_, _05236_, \oc8051_golden_model_1.ACC [4]);
  nor _70800_ (_19579_, _19578_, _19571_);
  nor _70801_ (_19581_, _19579_, _04427_);
  nor _70802_ (_19582_, _04426_, _19570_);
  or _70803_ (_19583_, _19582_, _19581_);
  and _70804_ (_19584_, _19583_, _04444_);
  nor _70805_ (_19585_, _12733_, _09015_);
  nor _70806_ (_19586_, _19585_, _19571_);
  nor _70807_ (_19587_, _19586_, _04444_);
  or _70808_ (_19588_, _19587_, _19584_);
  and _70809_ (_19589_, _19588_, _03517_);
  nor _70810_ (_19590_, _05799_, _19570_);
  and _70811_ (_19592_, _12737_, _05799_);
  nor _70812_ (_19593_, _19592_, _19590_);
  nor _70813_ (_19594_, _19593_, _03517_);
  or _70814_ (_19595_, _19594_, _03568_);
  or _70815_ (_19596_, _19595_, _19589_);
  nand _70816_ (_19597_, _19576_, _03568_);
  and _70817_ (_19598_, _19597_, _19596_);
  and _70818_ (_19599_, _19598_, _03583_);
  nor _70819_ (_19600_, _19579_, _03583_);
  or _70820_ (_19601_, _19600_, _19599_);
  and _70821_ (_19603_, _19601_, _03513_);
  and _70822_ (_19604_, _12718_, _05799_);
  nor _70823_ (_19605_, _19604_, _19590_);
  nor _70824_ (_19606_, _19605_, _03513_);
  or _70825_ (_19607_, _19606_, _19603_);
  and _70826_ (_19608_, _19607_, _03506_);
  nor _70827_ (_19609_, _19590_, _12752_);
  nor _70828_ (_19610_, _19609_, _19593_);
  and _70829_ (_19611_, _19610_, _03505_);
  or _70830_ (_19612_, _19611_, _19608_);
  and _70831_ (_19614_, _19612_, _03500_);
  nor _70832_ (_19615_, _12716_, _09052_);
  nor _70833_ (_19616_, _19615_, _19590_);
  nor _70834_ (_19617_, _19616_, _03500_);
  nor _70835_ (_19618_, _19617_, _07314_);
  not _70836_ (_19619_, _19618_);
  nor _70837_ (_19620_, _19619_, _19614_);
  nor _70838_ (_19621_, _19620_, _19577_);
  nor _70839_ (_19622_, _19621_, _03479_);
  and _70840_ (_19623_, _06722_, _05236_);
  nor _70841_ (_19625_, _19571_, _06044_);
  not _70842_ (_19626_, _19625_);
  nor _70843_ (_19627_, _19626_, _19623_);
  or _70844_ (_19628_, _19627_, _03221_);
  nor _70845_ (_19629_, _19628_, _19622_);
  nor _70846_ (_19630_, _12827_, _09015_);
  nor _70847_ (_19631_, _19630_, _19571_);
  nor _70848_ (_19632_, _19631_, _03474_);
  or _70849_ (_19633_, _19632_, _03437_);
  or _70850_ (_19634_, _19633_, _19629_);
  and _70851_ (_19636_, _06233_, _05236_);
  nor _70852_ (_19637_, _19636_, _19571_);
  nand _70853_ (_19638_, _19637_, _03437_);
  and _70854_ (_19639_, _19638_, _19634_);
  nor _70855_ (_19640_, _19639_, _03636_);
  and _70856_ (_19641_, _12711_, _05236_);
  or _70857_ (_19642_, _19571_, _04499_);
  nor _70858_ (_19643_, _19642_, _19641_);
  or _70859_ (_19644_, _19643_, _03769_);
  nor _70860_ (_19645_, _19644_, _19640_);
  nor _70861_ (_19647_, _19645_, _19574_);
  nor _70862_ (_19648_, _19647_, _04504_);
  not _70863_ (_19649_, _19571_);
  and _70864_ (_19650_, _19649_, _05760_);
  or _70865_ (_19651_, _19637_, _04505_);
  nor _70866_ (_19652_, _19651_, _19650_);
  nor _70867_ (_19653_, _19652_, _19648_);
  nor _70868_ (_19654_, _19653_, _03752_);
  or _70869_ (_19655_, _19650_, _03753_);
  nor _70870_ (_19656_, _19655_, _19579_);
  or _70871_ (_19658_, _19656_, _19654_);
  and _70872_ (_19659_, _19658_, _03759_);
  nor _70873_ (_19660_, _12710_, _09015_);
  nor _70874_ (_19661_, _19660_, _19571_);
  nor _70875_ (_19662_, _19661_, _03759_);
  or _70876_ (_19663_, _19662_, _19659_);
  and _70877_ (_19664_, _19663_, _04517_);
  nor _70878_ (_19665_, _12843_, _09015_);
  nor _70879_ (_19666_, _19665_, _19571_);
  nor _70880_ (_19667_, _19666_, _04517_);
  or _70881_ (_19669_, _19667_, _19664_);
  and _70882_ (_19670_, _19669_, _04192_);
  nor _70883_ (_19671_, _19586_, _04192_);
  or _70884_ (_19672_, _19671_, _19670_);
  and _70885_ (_19673_, _19672_, _03152_);
  nor _70886_ (_19674_, _19605_, _03152_);
  or _70887_ (_19675_, _19674_, _19673_);
  and _70888_ (_19676_, _19675_, _03521_);
  and _70889_ (_19677_, _12893_, _05236_);
  nor _70890_ (_19678_, _19677_, _19571_);
  nor _70891_ (_19680_, _19678_, _03521_);
  or _70892_ (_19681_, _19680_, _19676_);
  or _70893_ (_19682_, _19681_, _42967_);
  or _70894_ (_19683_, _42963_, \oc8051_golden_model_1.TCON [4]);
  and _70895_ (_19684_, _19683_, _41755_);
  and _70896_ (_43243_, _19684_, _19682_);
  not _70897_ (_19685_, \oc8051_golden_model_1.TCON [5]);
  nor _70898_ (_19686_, _05236_, _19685_);
  and _70899_ (_19687_, _13042_, _05236_);
  nor _70900_ (_19688_, _19687_, _19686_);
  nor _70901_ (_19690_, _19688_, _04501_);
  nor _70902_ (_19691_, _05422_, _09015_);
  nor _70903_ (_19692_, _19691_, _19686_);
  and _70904_ (_19693_, _19692_, _07314_);
  and _70905_ (_19694_, _05236_, \oc8051_golden_model_1.ACC [5]);
  nor _70906_ (_19695_, _19694_, _19686_);
  nor _70907_ (_19696_, _19695_, _04427_);
  nor _70908_ (_19697_, _04426_, _19685_);
  or _70909_ (_19698_, _19697_, _19696_);
  and _70910_ (_19699_, _19698_, _04444_);
  nor _70911_ (_19701_, _12930_, _09015_);
  nor _70912_ (_19702_, _19701_, _19686_);
  nor _70913_ (_19703_, _19702_, _04444_);
  or _70914_ (_19704_, _19703_, _19699_);
  and _70915_ (_19705_, _19704_, _03517_);
  nor _70916_ (_19706_, _05799_, _19685_);
  and _70917_ (_19707_, _12934_, _05799_);
  nor _70918_ (_19708_, _19707_, _19706_);
  nor _70919_ (_19709_, _19708_, _03517_);
  or _70920_ (_19710_, _19709_, _03568_);
  or _70921_ (_19712_, _19710_, _19705_);
  nand _70922_ (_19713_, _19692_, _03568_);
  and _70923_ (_19714_, _19713_, _19712_);
  and _70924_ (_19715_, _19714_, _03583_);
  nor _70925_ (_19716_, _19695_, _03583_);
  or _70926_ (_19717_, _19716_, _19715_);
  and _70927_ (_19718_, _19717_, _03513_);
  and _70928_ (_19719_, _12914_, _05799_);
  nor _70929_ (_19720_, _19719_, _19706_);
  nor _70930_ (_19721_, _19720_, _03513_);
  or _70931_ (_19723_, _19721_, _03505_);
  or _70932_ (_19724_, _19723_, _19718_);
  nor _70933_ (_19725_, _19706_, _12949_);
  nor _70934_ (_19726_, _19725_, _19708_);
  or _70935_ (_19727_, _19726_, _03506_);
  and _70936_ (_19728_, _19727_, _03500_);
  and _70937_ (_19729_, _19728_, _19724_);
  nor _70938_ (_19730_, _12912_, _09052_);
  nor _70939_ (_19731_, _19730_, _19706_);
  nor _70940_ (_19732_, _19731_, _03500_);
  nor _70941_ (_19734_, _19732_, _07314_);
  not _70942_ (_19735_, _19734_);
  nor _70943_ (_19736_, _19735_, _19729_);
  nor _70944_ (_19737_, _19736_, _19693_);
  nor _70945_ (_19738_, _19737_, _03479_);
  and _70946_ (_19739_, _06721_, _05236_);
  nor _70947_ (_19740_, _19686_, _06044_);
  not _70948_ (_19741_, _19740_);
  nor _70949_ (_19742_, _19741_, _19739_);
  or _70950_ (_19743_, _19742_, _03221_);
  nor _70951_ (_19745_, _19743_, _19738_);
  nor _70952_ (_19746_, _13021_, _09015_);
  nor _70953_ (_19747_, _19746_, _19686_);
  nor _70954_ (_19748_, _19747_, _03474_);
  or _70955_ (_19749_, _19748_, _03437_);
  or _70956_ (_19750_, _19749_, _19745_);
  and _70957_ (_19751_, _06211_, _05236_);
  nor _70958_ (_19752_, _19751_, _19686_);
  nand _70959_ (_19753_, _19752_, _03437_);
  and _70960_ (_19754_, _19753_, _19750_);
  nor _70961_ (_19756_, _19754_, _03636_);
  and _70962_ (_19757_, _13036_, _05236_);
  or _70963_ (_19758_, _19686_, _04499_);
  nor _70964_ (_19759_, _19758_, _19757_);
  or _70965_ (_19760_, _19759_, _03769_);
  nor _70966_ (_19761_, _19760_, _19756_);
  nor _70967_ (_19762_, _19761_, _19690_);
  nor _70968_ (_19763_, _19762_, _04504_);
  not _70969_ (_19764_, _19686_);
  and _70970_ (_19765_, _19764_, _05471_);
  or _70971_ (_19767_, _19752_, _04505_);
  nor _70972_ (_19768_, _19767_, _19765_);
  nor _70973_ (_19769_, _19768_, _19763_);
  nor _70974_ (_19770_, _19769_, _03752_);
  or _70975_ (_19771_, _19765_, _03753_);
  or _70976_ (_19772_, _19771_, _19695_);
  and _70977_ (_19773_, _19772_, _03759_);
  not _70978_ (_19774_, _19773_);
  nor _70979_ (_19775_, _19774_, _19770_);
  nor _70980_ (_19776_, _13035_, _09015_);
  or _70981_ (_19778_, _19686_, _03759_);
  nor _70982_ (_19779_, _19778_, _19776_);
  or _70983_ (_19780_, _19779_, _03760_);
  nor _70984_ (_19781_, _19780_, _19775_);
  nor _70985_ (_19782_, _13041_, _09015_);
  nor _70986_ (_19783_, _19782_, _19686_);
  nor _70987_ (_19784_, _19783_, _04517_);
  or _70988_ (_19785_, _19784_, _19781_);
  and _70989_ (_19786_, _19785_, _04192_);
  nor _70990_ (_19787_, _19702_, _04192_);
  or _70991_ (_19789_, _19787_, _19786_);
  and _70992_ (_19790_, _19789_, _03152_);
  nor _70993_ (_19791_, _19720_, _03152_);
  or _70994_ (_19792_, _19791_, _19790_);
  and _70995_ (_19793_, _19792_, _03521_);
  and _70996_ (_19794_, _13097_, _05236_);
  nor _70997_ (_19795_, _19794_, _19686_);
  nor _70998_ (_19796_, _19795_, _03521_);
  or _70999_ (_19797_, _19796_, _19793_);
  or _71000_ (_19798_, _19797_, _42967_);
  or _71001_ (_19800_, _42963_, \oc8051_golden_model_1.TCON [5]);
  and _71002_ (_19801_, _19800_, _41755_);
  and _71003_ (_43244_, _19801_, _19798_);
  not _71004_ (_19802_, \oc8051_golden_model_1.TCON [6]);
  nor _71005_ (_19803_, _05236_, _19802_);
  and _71006_ (_19804_, _13259_, _05236_);
  nor _71007_ (_19805_, _19804_, _19803_);
  nor _71008_ (_19806_, _19805_, _04501_);
  nor _71009_ (_19807_, _05327_, _09015_);
  nor _71010_ (_19808_, _19807_, _19803_);
  and _71011_ (_19810_, _19808_, _07314_);
  and _71012_ (_19811_, _05236_, \oc8051_golden_model_1.ACC [6]);
  nor _71013_ (_19812_, _19811_, _19803_);
  nor _71014_ (_19813_, _19812_, _04427_);
  nor _71015_ (_19814_, _04426_, _19802_);
  or _71016_ (_19815_, _19814_, _19813_);
  and _71017_ (_19816_, _19815_, _04444_);
  nor _71018_ (_19817_, _13122_, _09015_);
  nor _71019_ (_19818_, _19817_, _19803_);
  nor _71020_ (_19819_, _19818_, _04444_);
  or _71021_ (_19821_, _19819_, _19816_);
  and _71022_ (_19822_, _19821_, _03517_);
  nor _71023_ (_19823_, _05799_, _19802_);
  and _71024_ (_19824_, _13145_, _05799_);
  nor _71025_ (_19825_, _19824_, _19823_);
  nor _71026_ (_19826_, _19825_, _03517_);
  or _71027_ (_19827_, _19826_, _03568_);
  or _71028_ (_19828_, _19827_, _19822_);
  nand _71029_ (_19829_, _19808_, _03568_);
  and _71030_ (_19830_, _19829_, _19828_);
  and _71031_ (_19832_, _19830_, _03583_);
  nor _71032_ (_19833_, _19812_, _03583_);
  or _71033_ (_19834_, _19833_, _19832_);
  and _71034_ (_19835_, _19834_, _03513_);
  and _71035_ (_19836_, _13130_, _05799_);
  nor _71036_ (_19837_, _19836_, _19823_);
  nor _71037_ (_19838_, _19837_, _03513_);
  or _71038_ (_19839_, _19838_, _19835_);
  and _71039_ (_19840_, _19839_, _03506_);
  nor _71040_ (_19841_, _19823_, _13160_);
  nor _71041_ (_19843_, _19841_, _19825_);
  and _71042_ (_19844_, _19843_, _03505_);
  or _71043_ (_19845_, _19844_, _19840_);
  and _71044_ (_19846_, _19845_, _03500_);
  nor _71045_ (_19847_, _13178_, _09052_);
  nor _71046_ (_19848_, _19847_, _19823_);
  nor _71047_ (_19849_, _19848_, _03500_);
  nor _71048_ (_19850_, _19849_, _07314_);
  not _71049_ (_19851_, _19850_);
  nor _71050_ (_19852_, _19851_, _19846_);
  nor _71051_ (_19854_, _19852_, _19810_);
  nor _71052_ (_19855_, _19854_, _03479_);
  and _71053_ (_19856_, _06713_, _05236_);
  nor _71054_ (_19857_, _19803_, _06044_);
  not _71055_ (_19858_, _19857_);
  nor _71056_ (_19859_, _19858_, _19856_);
  or _71057_ (_19860_, _19859_, _03221_);
  nor _71058_ (_19861_, _19860_, _19855_);
  nor _71059_ (_19862_, _13237_, _09015_);
  nor _71060_ (_19863_, _19862_, _19803_);
  nor _71061_ (_19865_, _19863_, _03474_);
  or _71062_ (_19866_, _19865_, _03437_);
  or _71063_ (_19867_, _19866_, _19861_);
  and _71064_ (_19868_, _13244_, _05236_);
  nor _71065_ (_19869_, _19868_, _19803_);
  nand _71066_ (_19870_, _19869_, _03437_);
  and _71067_ (_19871_, _19870_, _19867_);
  nor _71068_ (_19872_, _19871_, _03636_);
  and _71069_ (_19873_, _13253_, _05236_);
  or _71070_ (_19874_, _19803_, _04499_);
  nor _71071_ (_19876_, _19874_, _19873_);
  or _71072_ (_19877_, _19876_, _03769_);
  nor _71073_ (_19878_, _19877_, _19872_);
  nor _71074_ (_19879_, _19878_, _19806_);
  nor _71075_ (_19880_, _19879_, _04504_);
  not _71076_ (_19881_, _19803_);
  and _71077_ (_19882_, _19881_, _05376_);
  or _71078_ (_19883_, _19869_, _04505_);
  nor _71079_ (_19884_, _19883_, _19882_);
  nor _71080_ (_19885_, _19884_, _19880_);
  nor _71081_ (_19887_, _19885_, _03752_);
  or _71082_ (_19888_, _19882_, _03753_);
  or _71083_ (_19889_, _19888_, _19812_);
  and _71084_ (_19890_, _19889_, _03759_);
  not _71085_ (_19891_, _19890_);
  nor _71086_ (_19892_, _19891_, _19887_);
  nor _71087_ (_19893_, _13251_, _09015_);
  or _71088_ (_19894_, _19803_, _03759_);
  nor _71089_ (_19895_, _19894_, _19893_);
  or _71090_ (_19896_, _19895_, _03760_);
  nor _71091_ (_19898_, _19896_, _19892_);
  nor _71092_ (_19899_, _13258_, _09015_);
  nor _71093_ (_19900_, _19899_, _19803_);
  nor _71094_ (_19901_, _19900_, _04517_);
  or _71095_ (_19902_, _19901_, _19898_);
  and _71096_ (_19903_, _19902_, _04192_);
  nor _71097_ (_19904_, _19818_, _04192_);
  or _71098_ (_19905_, _19904_, _19903_);
  and _71099_ (_19906_, _19905_, _03152_);
  nor _71100_ (_19907_, _19837_, _03152_);
  or _71101_ (_19909_, _19907_, _19906_);
  and _71102_ (_19910_, _19909_, _03521_);
  and _71103_ (_19911_, _13312_, _05236_);
  nor _71104_ (_19912_, _19911_, _19803_);
  nor _71105_ (_19913_, _19912_, _03521_);
  or _71106_ (_19914_, _19913_, _19910_);
  or _71107_ (_19915_, _19914_, _42967_);
  or _71108_ (_19916_, _42963_, \oc8051_golden_model_1.TCON [6]);
  and _71109_ (_19917_, _19916_, _41755_);
  and _71110_ (_43245_, _19917_, _19915_);
  not _71111_ (_19919_, \oc8051_golden_model_1.TL0 [0]);
  nor _71112_ (_19920_, _05258_, _19919_);
  and _71113_ (_19921_, _05941_, _05258_);
  nor _71114_ (_19922_, _19921_, _19920_);
  and _71115_ (_19923_, _19922_, _17076_);
  and _71116_ (_19924_, _05258_, \oc8051_golden_model_1.ACC [0]);
  nor _71117_ (_19925_, _19924_, _19920_);
  nor _71118_ (_19926_, _19925_, _03583_);
  nor _71119_ (_19927_, _19926_, _07314_);
  nor _71120_ (_19928_, _19922_, _04444_);
  nor _71121_ (_19930_, _04426_, _19919_);
  nor _71122_ (_19931_, _19925_, _04427_);
  nor _71123_ (_19932_, _19931_, _19930_);
  nor _71124_ (_19933_, _19932_, _03570_);
  or _71125_ (_19934_, _19933_, _03568_);
  nor _71126_ (_19935_, _19934_, _19928_);
  or _71127_ (_19936_, _19935_, _03575_);
  and _71128_ (_19937_, _19936_, _19927_);
  and _71129_ (_19938_, _05258_, _04419_);
  or _71130_ (_19939_, _19920_, _18522_);
  nor _71131_ (_19941_, _19939_, _19938_);
  nor _71132_ (_19942_, _19941_, _19937_);
  nor _71133_ (_19943_, _19942_, _03479_);
  and _71134_ (_19944_, _06715_, _05258_);
  nor _71135_ (_19945_, _19920_, _06044_);
  not _71136_ (_19946_, _19945_);
  nor _71137_ (_19947_, _19946_, _19944_);
  nor _71138_ (_19948_, _19947_, _19943_);
  nor _71139_ (_19949_, _19948_, _03221_);
  nor _71140_ (_19950_, _11975_, _09135_);
  or _71141_ (_19952_, _19920_, _03474_);
  nor _71142_ (_19953_, _19952_, _19950_);
  or _71143_ (_19954_, _19953_, _03437_);
  nor _71144_ (_19955_, _19954_, _19949_);
  and _71145_ (_19956_, _05258_, _06202_);
  nor _71146_ (_19957_, _19956_, _19920_);
  nor _71147_ (_19958_, _19957_, _03438_);
  or _71148_ (_19959_, _19958_, _19955_);
  and _71149_ (_19960_, _19959_, _04499_);
  and _71150_ (_19961_, _11990_, _05258_);
  nor _71151_ (_19963_, _19961_, _19920_);
  nor _71152_ (_19964_, _19963_, _04499_);
  or _71153_ (_19965_, _19964_, _19960_);
  nor _71154_ (_19966_, _19965_, _03769_);
  and _71155_ (_19967_, _11995_, _05258_);
  or _71156_ (_19968_, _19920_, _04501_);
  nor _71157_ (_19969_, _19968_, _19967_);
  or _71158_ (_19970_, _19969_, _04504_);
  nor _71159_ (_19971_, _19970_, _19966_);
  or _71160_ (_19972_, _19957_, _04505_);
  nor _71161_ (_19974_, _19972_, _19921_);
  nor _71162_ (_19975_, _19974_, _19971_);
  nor _71163_ (_19976_, _19975_, _03752_);
  nor _71164_ (_19977_, _19920_, _05617_);
  or _71165_ (_19978_, _19977_, _03753_);
  nor _71166_ (_19979_, _19978_, _19925_);
  or _71167_ (_19980_, _19979_, _19976_);
  and _71168_ (_19981_, _19980_, _03759_);
  nor _71169_ (_19982_, _11988_, _09135_);
  nor _71170_ (_19983_, _19982_, _19920_);
  nor _71171_ (_19985_, _19983_, _03759_);
  or _71172_ (_19986_, _19985_, _19981_);
  and _71173_ (_19987_, _19986_, _04517_);
  nor _71174_ (_19988_, _11870_, _09135_);
  nor _71175_ (_19989_, _19988_, _19920_);
  nor _71176_ (_19990_, _19989_, _04517_);
  nor _71177_ (_19991_, _19990_, _17076_);
  not _71178_ (_19992_, _19991_);
  nor _71179_ (_19993_, _19992_, _19987_);
  nor _71180_ (_19994_, _19993_, _19923_);
  or _71181_ (_19996_, _19994_, _42967_);
  or _71182_ (_19997_, _42963_, \oc8051_golden_model_1.TL0 [0]);
  and _71183_ (_19998_, _19997_, _41755_);
  and _71184_ (_43246_, _19998_, _19996_);
  and _71185_ (_19999_, _06714_, _05258_);
  not _71186_ (_20000_, \oc8051_golden_model_1.TL0 [1]);
  nor _71187_ (_20001_, _05258_, _20000_);
  nor _71188_ (_20002_, _20001_, _06044_);
  not _71189_ (_20003_, _20002_);
  nor _71190_ (_20004_, _20003_, _19999_);
  not _71191_ (_20006_, _20004_);
  nor _71192_ (_20007_, _05258_, \oc8051_golden_model_1.TL0 [1]);
  and _71193_ (_20008_, _05258_, _03233_);
  nor _71194_ (_20009_, _20008_, _20007_);
  and _71195_ (_20010_, _20009_, _03575_);
  nor _71196_ (_20011_, _09135_, _04603_);
  nor _71197_ (_20012_, _20011_, _20001_);
  nor _71198_ (_20013_, _20012_, _03983_);
  and _71199_ (_20014_, _20009_, _04426_);
  nor _71200_ (_20015_, _04426_, _20000_);
  or _71201_ (_20017_, _20015_, _20014_);
  and _71202_ (_20018_, _20017_, _04444_);
  and _71203_ (_20019_, _12252_, _05258_);
  nor _71204_ (_20020_, _20019_, _20007_);
  and _71205_ (_20021_, _20020_, _03570_);
  or _71206_ (_20022_, _20021_, _20018_);
  and _71207_ (_20023_, _20022_, _03983_);
  nor _71208_ (_20024_, _20023_, _20013_);
  nor _71209_ (_20025_, _20024_, _03575_);
  or _71210_ (_20026_, _20025_, _07314_);
  nor _71211_ (_20028_, _20026_, _20010_);
  and _71212_ (_20029_, _20012_, _07314_);
  nor _71213_ (_20030_, _20029_, _20028_);
  nor _71214_ (_20031_, _20030_, _03479_);
  nor _71215_ (_20032_, _20031_, _03221_);
  and _71216_ (_20033_, _20032_, _20006_);
  not _71217_ (_20034_, _20007_);
  and _71218_ (_20035_, _12176_, _05258_);
  nor _71219_ (_20036_, _20035_, _03474_);
  and _71220_ (_20037_, _20036_, _20034_);
  nor _71221_ (_20039_, _20037_, _20033_);
  nor _71222_ (_20040_, _20039_, _03437_);
  and _71223_ (_20041_, _05258_, _04317_);
  not _71224_ (_20042_, _20041_);
  nor _71225_ (_20043_, _20007_, _03438_);
  and _71226_ (_20044_, _20043_, _20042_);
  nor _71227_ (_20045_, _20044_, _20040_);
  nor _71228_ (_20046_, _20045_, _03636_);
  nor _71229_ (_20047_, _12191_, _09135_);
  nor _71230_ (_20048_, _20047_, _04499_);
  and _71231_ (_20050_, _20048_, _20034_);
  nor _71232_ (_20051_, _20050_, _20046_);
  nor _71233_ (_20052_, _20051_, _03769_);
  nor _71234_ (_20053_, _12197_, _09135_);
  nor _71235_ (_20054_, _20053_, _04501_);
  and _71236_ (_20055_, _20054_, _20034_);
  nor _71237_ (_20056_, _20055_, _20052_);
  nor _71238_ (_20057_, _20056_, _04504_);
  nor _71239_ (_20058_, _12190_, _09135_);
  nor _71240_ (_20059_, _20058_, _05769_);
  and _71241_ (_20061_, _20059_, _20034_);
  nor _71242_ (_20062_, _20061_, _20057_);
  nor _71243_ (_20063_, _20062_, _03752_);
  and _71244_ (_20064_, _12195_, _05258_);
  or _71245_ (_20065_, _20064_, _20001_);
  and _71246_ (_20066_, _20065_, _03752_);
  nor _71247_ (_20067_, _20066_, _20063_);
  nor _71248_ (_20068_, _20067_, _03758_);
  and _71249_ (_20069_, _20041_, _05940_);
  nor _71250_ (_20070_, _20069_, _03759_);
  and _71251_ (_20072_, _20070_, _20034_);
  nor _71252_ (_20073_, _20072_, _20068_);
  nor _71253_ (_20074_, _20073_, _03760_);
  and _71254_ (_20075_, _20008_, _05940_);
  nor _71255_ (_20076_, _20075_, _04517_);
  and _71256_ (_20077_, _20076_, _20034_);
  or _71257_ (_20078_, _20077_, _20074_);
  and _71258_ (_20079_, _20078_, _04192_);
  and _71259_ (_20080_, _20020_, _03790_);
  or _71260_ (_20081_, _20080_, _20079_);
  and _71261_ (_20083_, _20081_, _03521_);
  nor _71262_ (_20084_, _20001_, _20019_);
  nor _71263_ (_20085_, _20084_, _03521_);
  or _71264_ (_20086_, _20085_, _20083_);
  or _71265_ (_20087_, _20086_, _42967_);
  or _71266_ (_20088_, _42963_, \oc8051_golden_model_1.TL0 [1]);
  and _71267_ (_20089_, _20088_, _41755_);
  and _71268_ (_43247_, _20089_, _20087_);
  not _71269_ (_20090_, \oc8051_golden_model_1.TL0 [2]);
  nor _71270_ (_20091_, _05258_, _20090_);
  nor _71271_ (_20093_, _12400_, _09135_);
  nor _71272_ (_20094_, _20093_, _20091_);
  nor _71273_ (_20095_, _20094_, _04517_);
  and _71274_ (_20096_, _05258_, \oc8051_golden_model_1.ACC [2]);
  nor _71275_ (_20097_, _20096_, _20091_);
  nor _71276_ (_20098_, _20097_, _03583_);
  nor _71277_ (_20099_, _20097_, _04427_);
  nor _71278_ (_20100_, _04426_, _20090_);
  or _71279_ (_20101_, _20100_, _20099_);
  and _71280_ (_20102_, _20101_, _04444_);
  nor _71281_ (_20104_, _12282_, _09135_);
  nor _71282_ (_20105_, _20104_, _20091_);
  nor _71283_ (_20106_, _20105_, _04444_);
  or _71284_ (_20107_, _20106_, _20102_);
  and _71285_ (_20108_, _20107_, _03983_);
  nor _71286_ (_20109_, _09135_, _05026_);
  nor _71287_ (_20110_, _20109_, _20091_);
  nor _71288_ (_20111_, _20110_, _03983_);
  nor _71289_ (_20112_, _20111_, _20108_);
  nor _71290_ (_20113_, _20112_, _03575_);
  or _71291_ (_20115_, _20113_, _07314_);
  nor _71292_ (_20116_, _20115_, _20098_);
  and _71293_ (_20117_, _20110_, _07314_);
  nor _71294_ (_20118_, _20117_, _20116_);
  nor _71295_ (_20119_, _20118_, _03479_);
  and _71296_ (_20120_, _06718_, _05258_);
  nor _71297_ (_20121_, _20091_, _06044_);
  not _71298_ (_20122_, _20121_);
  nor _71299_ (_20123_, _20122_, _20120_);
  nor _71300_ (_20124_, _20123_, _20119_);
  nor _71301_ (_20126_, _20124_, _03221_);
  nor _71302_ (_20127_, _12384_, _09135_);
  or _71303_ (_20128_, _20091_, _03474_);
  nor _71304_ (_20129_, _20128_, _20127_);
  or _71305_ (_20130_, _20129_, _03437_);
  nor _71306_ (_20131_, _20130_, _20126_);
  and _71307_ (_20132_, _05258_, _06261_);
  nor _71308_ (_20133_, _20132_, _20091_);
  nor _71309_ (_20134_, _20133_, _03438_);
  or _71310_ (_20135_, _20134_, _20131_);
  and _71311_ (_20137_, _20135_, _04499_);
  and _71312_ (_20138_, _12273_, _05258_);
  nor _71313_ (_20139_, _20138_, _20091_);
  nor _71314_ (_20140_, _20139_, _04499_);
  or _71315_ (_20141_, _20140_, _20137_);
  nor _71316_ (_20142_, _20141_, _03769_);
  and _71317_ (_20143_, _12401_, _05258_);
  or _71318_ (_20144_, _20091_, _04501_);
  nor _71319_ (_20145_, _20144_, _20143_);
  or _71320_ (_20146_, _20145_, _04504_);
  nor _71321_ (_20148_, _20146_, _20142_);
  nor _71322_ (_20149_, _20091_, _05665_);
  or _71323_ (_20150_, _20133_, _04505_);
  nor _71324_ (_20151_, _20150_, _20149_);
  nor _71325_ (_20152_, _20151_, _20148_);
  nor _71326_ (_20153_, _20152_, _03752_);
  or _71327_ (_20154_, _20149_, _03753_);
  or _71328_ (_20155_, _20154_, _20097_);
  and _71329_ (_20156_, _20155_, _03759_);
  not _71330_ (_20157_, _20156_);
  nor _71331_ (_20159_, _20157_, _20153_);
  nor _71332_ (_20160_, _12272_, _09135_);
  or _71333_ (_20161_, _20091_, _03759_);
  nor _71334_ (_20162_, _20161_, _20160_);
  or _71335_ (_20163_, _20162_, _03760_);
  nor _71336_ (_20164_, _20163_, _20159_);
  nor _71337_ (_20165_, _20164_, _20095_);
  nor _71338_ (_20166_, _20165_, _03790_);
  nor _71339_ (_20167_, _20105_, _04192_);
  or _71340_ (_20168_, _20167_, _03520_);
  nor _71341_ (_20170_, _20168_, _20166_);
  and _71342_ (_20171_, _12456_, _05258_);
  or _71343_ (_20172_, _20091_, _03521_);
  nor _71344_ (_20173_, _20172_, _20171_);
  nor _71345_ (_20174_, _20173_, _20170_);
  or _71346_ (_20175_, _20174_, _42967_);
  or _71347_ (_20176_, _42963_, \oc8051_golden_model_1.TL0 [2]);
  and _71348_ (_20177_, _20176_, _41755_);
  and _71349_ (_43248_, _20177_, _20175_);
  not _71350_ (_20178_, \oc8051_golden_model_1.TL0 [3]);
  nor _71351_ (_20180_, _05258_, _20178_);
  and _71352_ (_20181_, _12604_, _05258_);
  nor _71353_ (_20182_, _20181_, _20180_);
  nor _71354_ (_20183_, _20182_, _04501_);
  and _71355_ (_20184_, _05258_, \oc8051_golden_model_1.ACC [3]);
  nor _71356_ (_20185_, _20184_, _20180_);
  nor _71357_ (_20186_, _20185_, _03583_);
  nor _71358_ (_20187_, _20185_, _04427_);
  nor _71359_ (_20188_, _04426_, _20178_);
  or _71360_ (_20189_, _20188_, _20187_);
  and _71361_ (_20191_, _20189_, _04444_);
  nor _71362_ (_20192_, _12486_, _09135_);
  nor _71363_ (_20193_, _20192_, _20180_);
  nor _71364_ (_20194_, _20193_, _04444_);
  or _71365_ (_20195_, _20194_, _20191_);
  and _71366_ (_20196_, _20195_, _03983_);
  nor _71367_ (_20197_, _09135_, _04843_);
  nor _71368_ (_20198_, _20197_, _20180_);
  nor _71369_ (_20199_, _20198_, _03983_);
  nor _71370_ (_20200_, _20199_, _20196_);
  nor _71371_ (_20202_, _20200_, _03575_);
  or _71372_ (_20203_, _20202_, _07314_);
  nor _71373_ (_20204_, _20203_, _20186_);
  and _71374_ (_20205_, _20198_, _07314_);
  nor _71375_ (_20206_, _20205_, _20204_);
  nor _71376_ (_20207_, _20206_, _03479_);
  and _71377_ (_20208_, _06717_, _05258_);
  nor _71378_ (_20209_, _20180_, _06044_);
  not _71379_ (_20210_, _20209_);
  nor _71380_ (_20211_, _20210_, _20208_);
  or _71381_ (_20213_, _20211_, _03221_);
  nor _71382_ (_20214_, _20213_, _20207_);
  nor _71383_ (_20215_, _12583_, _09135_);
  nor _71384_ (_20216_, _20215_, _20180_);
  nor _71385_ (_20217_, _20216_, _03474_);
  or _71386_ (_20218_, _20217_, _03437_);
  or _71387_ (_20219_, _20218_, _20214_);
  and _71388_ (_20220_, _05258_, _06217_);
  nor _71389_ (_20221_, _20220_, _20180_);
  nand _71390_ (_20222_, _20221_, _03437_);
  and _71391_ (_20224_, _20222_, _20219_);
  nor _71392_ (_20225_, _20224_, _03636_);
  and _71393_ (_20226_, _12598_, _05258_);
  or _71394_ (_20227_, _20180_, _04499_);
  nor _71395_ (_20228_, _20227_, _20226_);
  or _71396_ (_20229_, _20228_, _03769_);
  nor _71397_ (_20230_, _20229_, _20225_);
  nor _71398_ (_20231_, _20230_, _20183_);
  nor _71399_ (_20232_, _20231_, _04504_);
  not _71400_ (_20233_, _20180_);
  and _71401_ (_20235_, _20233_, _05520_);
  or _71402_ (_20236_, _20221_, _04505_);
  nor _71403_ (_20237_, _20236_, _20235_);
  nor _71404_ (_20238_, _20237_, _20232_);
  nor _71405_ (_20239_, _20238_, _03752_);
  or _71406_ (_20240_, _20235_, _03753_);
  nor _71407_ (_20241_, _20240_, _20185_);
  or _71408_ (_20242_, _20241_, _20239_);
  and _71409_ (_20243_, _20242_, _03759_);
  nor _71410_ (_20244_, _12597_, _09135_);
  nor _71411_ (_20246_, _20244_, _20180_);
  nor _71412_ (_20247_, _20246_, _03759_);
  or _71413_ (_20248_, _20247_, _20243_);
  and _71414_ (_20249_, _20248_, _04517_);
  nor _71415_ (_20250_, _12603_, _09135_);
  nor _71416_ (_20251_, _20250_, _20180_);
  nor _71417_ (_20252_, _20251_, _04517_);
  or _71418_ (_20253_, _20252_, _03790_);
  nor _71419_ (_20254_, _20253_, _20249_);
  and _71420_ (_20255_, _20193_, _03790_);
  or _71421_ (_20257_, _20255_, _03520_);
  nor _71422_ (_20258_, _20257_, _20254_);
  and _71423_ (_20259_, _12658_, _05258_);
  nor _71424_ (_20260_, _20259_, _20180_);
  nor _71425_ (_20261_, _20260_, _03521_);
  or _71426_ (_20262_, _20261_, _20258_);
  or _71427_ (_20263_, _20262_, _42967_);
  or _71428_ (_20264_, _42963_, \oc8051_golden_model_1.TL0 [3]);
  and _71429_ (_20265_, _20264_, _41755_);
  and _71430_ (_43249_, _20265_, _20263_);
  not _71431_ (_20267_, \oc8051_golden_model_1.TL0 [4]);
  nor _71432_ (_20268_, _05258_, _20267_);
  and _71433_ (_20269_, _12844_, _05258_);
  nor _71434_ (_20270_, _20269_, _20268_);
  nor _71435_ (_20271_, _20270_, _04501_);
  and _71436_ (_20272_, _05258_, \oc8051_golden_model_1.ACC [4]);
  nor _71437_ (_20273_, _20272_, _20268_);
  nor _71438_ (_20274_, _20273_, _03583_);
  nor _71439_ (_20275_, _20273_, _04427_);
  nor _71440_ (_20276_, _04426_, _20267_);
  or _71441_ (_20278_, _20276_, _20275_);
  and _71442_ (_20279_, _20278_, _04444_);
  nor _71443_ (_20280_, _12733_, _09135_);
  nor _71444_ (_20281_, _20280_, _20268_);
  nor _71445_ (_20282_, _20281_, _04444_);
  or _71446_ (_20283_, _20282_, _20279_);
  and _71447_ (_20284_, _20283_, _03983_);
  nor _71448_ (_20285_, _05712_, _09135_);
  nor _71449_ (_20286_, _20285_, _20268_);
  nor _71450_ (_20287_, _20286_, _03983_);
  nor _71451_ (_20289_, _20287_, _20284_);
  nor _71452_ (_20290_, _20289_, _03575_);
  or _71453_ (_20291_, _20290_, _07314_);
  nor _71454_ (_20292_, _20291_, _20274_);
  and _71455_ (_20293_, _20286_, _07314_);
  or _71456_ (_20294_, _20293_, _03479_);
  nor _71457_ (_20295_, _20294_, _20292_);
  and _71458_ (_20296_, _06722_, _05258_);
  or _71459_ (_20297_, _20296_, _20268_);
  and _71460_ (_20298_, _20297_, _03479_);
  or _71461_ (_20300_, _20298_, _03221_);
  or _71462_ (_20301_, _20300_, _20295_);
  nor _71463_ (_20302_, _12827_, _09135_);
  or _71464_ (_20303_, _20268_, _03474_);
  or _71465_ (_20304_, _20303_, _20302_);
  and _71466_ (_20305_, _20304_, _03438_);
  and _71467_ (_20306_, _20305_, _20301_);
  and _71468_ (_20307_, _06233_, _05258_);
  nor _71469_ (_20308_, _20307_, _20268_);
  nor _71470_ (_20309_, _20308_, _03438_);
  or _71471_ (_20311_, _20309_, _03636_);
  nor _71472_ (_20312_, _20311_, _20306_);
  and _71473_ (_20313_, _12711_, _05258_);
  or _71474_ (_20314_, _20268_, _04499_);
  nor _71475_ (_20315_, _20314_, _20313_);
  or _71476_ (_20316_, _20315_, _03769_);
  nor _71477_ (_20317_, _20316_, _20312_);
  nor _71478_ (_20318_, _20317_, _20271_);
  nor _71479_ (_20319_, _20318_, _04504_);
  not _71480_ (_20320_, _20268_);
  and _71481_ (_20322_, _20320_, _05760_);
  or _71482_ (_20323_, _20308_, _04505_);
  nor _71483_ (_20324_, _20323_, _20322_);
  nor _71484_ (_20325_, _20324_, _20319_);
  nor _71485_ (_20326_, _20325_, _03752_);
  or _71486_ (_20327_, _20322_, _03753_);
  nor _71487_ (_20328_, _20327_, _20273_);
  or _71488_ (_20329_, _20328_, _20326_);
  and _71489_ (_20330_, _20329_, _03759_);
  nor _71490_ (_20331_, _12710_, _09135_);
  nor _71491_ (_20333_, _20331_, _20268_);
  nor _71492_ (_20334_, _20333_, _03759_);
  or _71493_ (_20335_, _20334_, _20330_);
  and _71494_ (_20336_, _20335_, _04517_);
  nor _71495_ (_20337_, _12843_, _09135_);
  nor _71496_ (_20338_, _20337_, _20268_);
  nor _71497_ (_20339_, _20338_, _04517_);
  or _71498_ (_20340_, _20339_, _03790_);
  nor _71499_ (_20341_, _20340_, _20336_);
  and _71500_ (_20342_, _20281_, _03790_);
  or _71501_ (_20343_, _20342_, _03520_);
  nor _71502_ (_20344_, _20343_, _20341_);
  and _71503_ (_20345_, _12893_, _05258_);
  nor _71504_ (_20346_, _20345_, _20268_);
  nor _71505_ (_20347_, _20346_, _03521_);
  or _71506_ (_20348_, _20347_, _20344_);
  or _71507_ (_20349_, _20348_, _42967_);
  or _71508_ (_20350_, _42963_, \oc8051_golden_model_1.TL0 [4]);
  and _71509_ (_20351_, _20350_, _41755_);
  and _71510_ (_43250_, _20351_, _20349_);
  not _71511_ (_20353_, \oc8051_golden_model_1.TL0 [5]);
  nor _71512_ (_20354_, _05258_, _20353_);
  and _71513_ (_20355_, _13042_, _05258_);
  nor _71514_ (_20356_, _20355_, _20354_);
  nor _71515_ (_20357_, _20356_, _04501_);
  and _71516_ (_20358_, _05258_, \oc8051_golden_model_1.ACC [5]);
  nor _71517_ (_20359_, _20358_, _20354_);
  nor _71518_ (_20360_, _20359_, _03583_);
  nor _71519_ (_20361_, _20359_, _04427_);
  nor _71520_ (_20362_, _04426_, _20353_);
  or _71521_ (_20364_, _20362_, _20361_);
  and _71522_ (_20365_, _20364_, _04444_);
  nor _71523_ (_20366_, _12930_, _09135_);
  nor _71524_ (_20367_, _20366_, _20354_);
  nor _71525_ (_20368_, _20367_, _04444_);
  or _71526_ (_20369_, _20368_, _20365_);
  and _71527_ (_20370_, _20369_, _03983_);
  nor _71528_ (_20371_, _05422_, _09135_);
  nor _71529_ (_20372_, _20371_, _20354_);
  nor _71530_ (_20373_, _20372_, _03983_);
  nor _71531_ (_20375_, _20373_, _20370_);
  nor _71532_ (_20376_, _20375_, _03575_);
  or _71533_ (_20377_, _20376_, _07314_);
  nor _71534_ (_20378_, _20377_, _20360_);
  and _71535_ (_20379_, _20372_, _07314_);
  nor _71536_ (_20380_, _20379_, _20378_);
  nor _71537_ (_20381_, _20380_, _03479_);
  and _71538_ (_20382_, _06721_, _05258_);
  nor _71539_ (_20383_, _20354_, _06044_);
  not _71540_ (_20384_, _20383_);
  nor _71541_ (_20385_, _20384_, _20382_);
  or _71542_ (_20386_, _20385_, _03221_);
  nor _71543_ (_20387_, _20386_, _20381_);
  nor _71544_ (_20388_, _13021_, _09135_);
  nor _71545_ (_20389_, _20388_, _20354_);
  nor _71546_ (_20390_, _20389_, _03474_);
  or _71547_ (_20391_, _20390_, _03437_);
  or _71548_ (_20392_, _20391_, _20387_);
  and _71549_ (_20393_, _06211_, _05258_);
  nor _71550_ (_20394_, _20393_, _20354_);
  nand _71551_ (_20396_, _20394_, _03437_);
  and _71552_ (_20397_, _20396_, _20392_);
  nor _71553_ (_20398_, _20397_, _03636_);
  and _71554_ (_20399_, _13036_, _05258_);
  or _71555_ (_20400_, _20354_, _04499_);
  nor _71556_ (_20401_, _20400_, _20399_);
  or _71557_ (_20402_, _20401_, _03769_);
  nor _71558_ (_20403_, _20402_, _20398_);
  nor _71559_ (_20404_, _20403_, _20357_);
  nor _71560_ (_20405_, _20404_, _04504_);
  not _71561_ (_20406_, _20354_);
  and _71562_ (_20407_, _20406_, _05471_);
  or _71563_ (_20408_, _20394_, _04505_);
  nor _71564_ (_20409_, _20408_, _20407_);
  nor _71565_ (_20410_, _20409_, _20405_);
  nor _71566_ (_20411_, _20410_, _03752_);
  or _71567_ (_20412_, _20407_, _03753_);
  or _71568_ (_20413_, _20412_, _20359_);
  and _71569_ (_20414_, _20413_, _03759_);
  not _71570_ (_20415_, _20414_);
  nor _71571_ (_20417_, _20415_, _20411_);
  nor _71572_ (_20418_, _13035_, _09135_);
  or _71573_ (_20419_, _20354_, _03759_);
  nor _71574_ (_20420_, _20419_, _20418_);
  or _71575_ (_20421_, _20420_, _03760_);
  nor _71576_ (_20422_, _20421_, _20417_);
  nor _71577_ (_20423_, _13041_, _09135_);
  nor _71578_ (_20424_, _20423_, _20354_);
  nor _71579_ (_20425_, _20424_, _04517_);
  or _71580_ (_20426_, _20425_, _03790_);
  nor _71581_ (_20428_, _20426_, _20422_);
  and _71582_ (_20429_, _20367_, _03790_);
  or _71583_ (_20430_, _20429_, _03520_);
  nor _71584_ (_20431_, _20430_, _20428_);
  and _71585_ (_20432_, _13097_, _05258_);
  nor _71586_ (_20433_, _20432_, _20354_);
  nor _71587_ (_20434_, _20433_, _03521_);
  or _71588_ (_20435_, _20434_, _20431_);
  or _71589_ (_20436_, _20435_, _42967_);
  or _71590_ (_20437_, _42963_, \oc8051_golden_model_1.TL0 [5]);
  and _71591_ (_20438_, _20437_, _41755_);
  and _71592_ (_43251_, _20438_, _20436_);
  not _71593_ (_20439_, \oc8051_golden_model_1.TL0 [6]);
  nor _71594_ (_20440_, _05258_, _20439_);
  and _71595_ (_20441_, _13259_, _05258_);
  nor _71596_ (_20442_, _20441_, _20440_);
  nor _71597_ (_20443_, _20442_, _04501_);
  and _71598_ (_20444_, _05258_, \oc8051_golden_model_1.ACC [6]);
  nor _71599_ (_20445_, _20444_, _20440_);
  nor _71600_ (_20446_, _20445_, _03583_);
  nor _71601_ (_20448_, _20445_, _04427_);
  nor _71602_ (_20449_, _04426_, _20439_);
  or _71603_ (_20450_, _20449_, _20448_);
  and _71604_ (_20451_, _20450_, _04444_);
  nor _71605_ (_20452_, _13122_, _09135_);
  nor _71606_ (_20453_, _20452_, _20440_);
  nor _71607_ (_20454_, _20453_, _04444_);
  or _71608_ (_20455_, _20454_, _20451_);
  and _71609_ (_20456_, _20455_, _03983_);
  nor _71610_ (_20457_, _05327_, _09135_);
  nor _71611_ (_20459_, _20457_, _20440_);
  nor _71612_ (_20460_, _20459_, _03983_);
  nor _71613_ (_20461_, _20460_, _20456_);
  nor _71614_ (_20462_, _20461_, _03575_);
  or _71615_ (_20463_, _20462_, _07314_);
  nor _71616_ (_20464_, _20463_, _20446_);
  and _71617_ (_20465_, _20459_, _07314_);
  nor _71618_ (_20466_, _20465_, _20464_);
  nor _71619_ (_20467_, _20466_, _03479_);
  and _71620_ (_20468_, _06713_, _05258_);
  nor _71621_ (_20469_, _20440_, _06044_);
  not _71622_ (_20470_, _20469_);
  nor _71623_ (_20471_, _20470_, _20468_);
  or _71624_ (_20472_, _20471_, _03221_);
  nor _71625_ (_20473_, _20472_, _20467_);
  nor _71626_ (_20474_, _13237_, _09135_);
  nor _71627_ (_20475_, _20474_, _20440_);
  nor _71628_ (_20476_, _20475_, _03474_);
  or _71629_ (_20477_, _20476_, _03437_);
  or _71630_ (_20478_, _20477_, _20473_);
  and _71631_ (_20480_, _13244_, _05258_);
  nor _71632_ (_20481_, _20480_, _20440_);
  nand _71633_ (_20482_, _20481_, _03437_);
  and _71634_ (_20483_, _20482_, _20478_);
  nor _71635_ (_20484_, _20483_, _03636_);
  and _71636_ (_20485_, _13253_, _05258_);
  or _71637_ (_20486_, _20440_, _04499_);
  nor _71638_ (_20487_, _20486_, _20485_);
  or _71639_ (_20488_, _20487_, _03769_);
  nor _71640_ (_20489_, _20488_, _20484_);
  nor _71641_ (_20491_, _20489_, _20443_);
  nor _71642_ (_20492_, _20491_, _04504_);
  not _71643_ (_20493_, _20440_);
  and _71644_ (_20494_, _20493_, _05376_);
  or _71645_ (_20495_, _20481_, _04505_);
  nor _71646_ (_20496_, _20495_, _20494_);
  nor _71647_ (_20497_, _20496_, _20492_);
  nor _71648_ (_20498_, _20497_, _03752_);
  or _71649_ (_20499_, _20494_, _03753_);
  or _71650_ (_20500_, _20499_, _20445_);
  and _71651_ (_20501_, _20500_, _03759_);
  not _71652_ (_20502_, _20501_);
  nor _71653_ (_20503_, _20502_, _20498_);
  nor _71654_ (_20504_, _13251_, _09135_);
  or _71655_ (_20505_, _20440_, _03759_);
  nor _71656_ (_20506_, _20505_, _20504_);
  or _71657_ (_20507_, _20506_, _03760_);
  nor _71658_ (_20508_, _20507_, _20503_);
  nor _71659_ (_20509_, _13258_, _09135_);
  nor _71660_ (_20510_, _20509_, _20440_);
  nor _71661_ (_20512_, _20510_, _04517_);
  or _71662_ (_20513_, _20512_, _03790_);
  nor _71663_ (_20514_, _20513_, _20508_);
  and _71664_ (_20515_, _20453_, _03790_);
  or _71665_ (_20516_, _20515_, _03520_);
  nor _71666_ (_20517_, _20516_, _20514_);
  and _71667_ (_20518_, _13312_, _05258_);
  nor _71668_ (_20519_, _20518_, _20440_);
  nor _71669_ (_20520_, _20519_, _03521_);
  or _71670_ (_20521_, _20520_, _20517_);
  or _71671_ (_20523_, _20521_, _42967_);
  or _71672_ (_20524_, _42963_, \oc8051_golden_model_1.TL0 [6]);
  and _71673_ (_20525_, _20524_, _41755_);
  and _71674_ (_43252_, _20525_, _20523_);
  not _71675_ (_20526_, \oc8051_golden_model_1.TL1 [0]);
  nor _71676_ (_20527_, _05242_, _20526_);
  and _71677_ (_20528_, _05941_, _05444_);
  nor _71678_ (_20529_, _20528_, _20527_);
  and _71679_ (_20530_, _20529_, _17076_);
  and _71680_ (_20531_, _05242_, \oc8051_golden_model_1.ACC [0]);
  nor _71681_ (_20532_, _20531_, _20527_);
  nor _71682_ (_20533_, _20532_, _03583_);
  nor _71683_ (_20534_, _20533_, _07314_);
  nor _71684_ (_20535_, _20529_, _04444_);
  nor _71685_ (_20536_, _04426_, _20526_);
  nor _71686_ (_20537_, _20532_, _04427_);
  nor _71687_ (_20538_, _20537_, _20536_);
  nor _71688_ (_20539_, _20538_, _03570_);
  or _71689_ (_20540_, _20539_, _03568_);
  nor _71690_ (_20541_, _20540_, _20535_);
  or _71691_ (_20543_, _20541_, _03575_);
  and _71692_ (_20544_, _20543_, _20534_);
  or _71693_ (_20545_, _09205_, _04439_);
  nor _71694_ (_20546_, _20527_, _18522_);
  and _71695_ (_20547_, _20546_, _20545_);
  nor _71696_ (_20548_, _20547_, _20544_);
  nor _71697_ (_20549_, _20548_, _03479_);
  nor _71698_ (_20550_, _20527_, _06044_);
  or _71699_ (_20551_, _06478_, _09205_);
  and _71700_ (_20552_, _20551_, _20550_);
  nor _71701_ (_20554_, _20552_, _20549_);
  nor _71702_ (_20555_, _20554_, _03221_);
  or _71703_ (_20556_, _11975_, _09205_);
  nor _71704_ (_20557_, _20527_, _03474_);
  and _71705_ (_20558_, _20557_, _20556_);
  or _71706_ (_20559_, _20558_, _03437_);
  nor _71707_ (_20560_, _20559_, _20555_);
  and _71708_ (_20561_, _05242_, _06202_);
  nor _71709_ (_20562_, _20561_, _20527_);
  nor _71710_ (_20563_, _20562_, _03438_);
  or _71711_ (_20564_, _20563_, _20560_);
  and _71712_ (_20565_, _20564_, _04499_);
  and _71713_ (_20566_, _11990_, _05242_);
  nor _71714_ (_20567_, _20566_, _20527_);
  nor _71715_ (_20568_, _20567_, _04499_);
  or _71716_ (_20569_, _20568_, _20565_);
  nor _71717_ (_20570_, _20569_, _03769_);
  nand _71718_ (_20571_, _11995_, _05444_);
  nor _71719_ (_20572_, _20527_, _04501_);
  and _71720_ (_20573_, _20572_, _20571_);
  or _71721_ (_20575_, _20573_, _04504_);
  nor _71722_ (_20576_, _20575_, _20570_);
  or _71723_ (_20577_, _20562_, _04505_);
  nor _71724_ (_20578_, _20577_, _20528_);
  nor _71725_ (_20579_, _20578_, _20576_);
  nor _71726_ (_20580_, _20579_, _03752_);
  nor _71727_ (_20581_, _20527_, _05617_);
  or _71728_ (_20582_, _20581_, _03753_);
  nor _71729_ (_20583_, _20582_, _20532_);
  or _71730_ (_20584_, _20583_, _20580_);
  and _71731_ (_20586_, _20584_, _03759_);
  nor _71732_ (_20587_, _11988_, _09229_);
  nor _71733_ (_20588_, _20587_, _20527_);
  nor _71734_ (_20589_, _20588_, _03759_);
  or _71735_ (_20590_, _20589_, _20586_);
  and _71736_ (_20591_, _20590_, _04517_);
  nor _71737_ (_20592_, _11870_, _09205_);
  nor _71738_ (_20593_, _20592_, _20527_);
  nor _71739_ (_20594_, _20593_, _04517_);
  nor _71740_ (_20595_, _20594_, _17076_);
  not _71741_ (_20596_, _20595_);
  nor _71742_ (_20597_, _20596_, _20591_);
  nor _71743_ (_20598_, _20597_, _20530_);
  or _71744_ (_20599_, _20598_, _42967_);
  or _71745_ (_20600_, _42963_, \oc8051_golden_model_1.TL1 [0]);
  and _71746_ (_20601_, _20600_, _41755_);
  and _71747_ (_43255_, _20601_, _20599_);
  not _71748_ (_20602_, \oc8051_golden_model_1.TL1 [1]);
  nor _71749_ (_20603_, _05242_, _20602_);
  and _71750_ (_20604_, _05242_, \oc8051_golden_model_1.ACC [1]);
  or _71751_ (_20606_, _20604_, _20603_);
  and _71752_ (_20607_, _20606_, _03575_);
  nor _71753_ (_20608_, _09205_, _04603_);
  nor _71754_ (_20609_, _20608_, _20603_);
  nor _71755_ (_20610_, _20609_, _03983_);
  and _71756_ (_20611_, _20606_, _04426_);
  nor _71757_ (_20612_, _04426_, _20602_);
  or _71758_ (_20613_, _20612_, _20611_);
  and _71759_ (_20614_, _20613_, _04444_);
  nor _71760_ (_20615_, _05242_, \oc8051_golden_model_1.TL1 [1]);
  and _71761_ (_20617_, _12252_, _05242_);
  nor _71762_ (_20618_, _20617_, _20615_);
  and _71763_ (_20619_, _20618_, _03570_);
  or _71764_ (_20620_, _20619_, _20614_);
  and _71765_ (_20621_, _20620_, _03983_);
  nor _71766_ (_20622_, _20621_, _20610_);
  nor _71767_ (_20623_, _20622_, _03575_);
  or _71768_ (_20624_, _20623_, _07314_);
  nor _71769_ (_20625_, _20624_, _20607_);
  and _71770_ (_20626_, _20609_, _07314_);
  nor _71771_ (_20627_, _20626_, _20625_);
  nor _71772_ (_20628_, _20627_, _03479_);
  nor _71773_ (_20629_, _20628_, _03221_);
  nor _71774_ (_20630_, _20603_, _06044_);
  or _71775_ (_20631_, _06433_, _09205_);
  nand _71776_ (_20632_, _20631_, _20630_);
  and _71777_ (_20633_, _20632_, _20629_);
  not _71778_ (_20634_, _20615_);
  nand _71779_ (_20635_, _12176_, _05242_);
  and _71780_ (_20636_, _20635_, _03221_);
  and _71781_ (_20638_, _20636_, _20634_);
  nor _71782_ (_20639_, _20638_, _20633_);
  nor _71783_ (_20640_, _20639_, _03437_);
  nor _71784_ (_20641_, _20615_, _03438_);
  nand _71785_ (_20642_, _05242_, _04317_);
  and _71786_ (_20643_, _20642_, _20641_);
  nor _71787_ (_20644_, _20643_, _20640_);
  nor _71788_ (_20645_, _20644_, _03636_);
  or _71789_ (_20646_, _12191_, _09229_);
  and _71790_ (_20647_, _20646_, _03636_);
  and _71791_ (_20649_, _20647_, _20634_);
  nor _71792_ (_20650_, _20649_, _20645_);
  nor _71793_ (_20651_, _20650_, _03769_);
  or _71794_ (_20652_, _12197_, _09229_);
  and _71795_ (_20653_, _20652_, _03769_);
  and _71796_ (_20654_, _20653_, _20634_);
  nor _71797_ (_20655_, _20654_, _20651_);
  nor _71798_ (_20656_, _20655_, _04504_);
  nor _71799_ (_20657_, _12190_, _09229_);
  nor _71800_ (_20658_, _20657_, _05769_);
  and _71801_ (_20659_, _20658_, _20634_);
  nor _71802_ (_20660_, _20659_, _20656_);
  nor _71803_ (_20661_, _20660_, _03752_);
  nor _71804_ (_20662_, _20603_, _05569_);
  nor _71805_ (_20663_, _20662_, _03753_);
  and _71806_ (_20664_, _20663_, _20606_);
  nor _71807_ (_20665_, _20664_, _20661_);
  nor _71808_ (_20666_, _20665_, _03758_);
  or _71809_ (_20667_, _20642_, _05569_);
  and _71810_ (_20668_, _20667_, _03758_);
  and _71811_ (_20670_, _20668_, _20634_);
  nor _71812_ (_20671_, _20670_, _20666_);
  nor _71813_ (_20672_, _20671_, _03760_);
  and _71814_ (_20673_, _12196_, _05242_);
  nor _71815_ (_20674_, _20673_, _04517_);
  and _71816_ (_20675_, _20674_, _20634_);
  or _71817_ (_20676_, _20675_, _20672_);
  and _71818_ (_20677_, _20676_, _04192_);
  and _71819_ (_20678_, _20618_, _03790_);
  or _71820_ (_20679_, _20678_, _20677_);
  and _71821_ (_20681_, _20679_, _03521_);
  nor _71822_ (_20682_, _20603_, _20617_);
  nor _71823_ (_20683_, _20682_, _03521_);
  or _71824_ (_20684_, _20683_, _20681_);
  or _71825_ (_20685_, _20684_, _42967_);
  or _71826_ (_20686_, _42963_, \oc8051_golden_model_1.TL1 [1]);
  and _71827_ (_20687_, _20686_, _41755_);
  and _71828_ (_43256_, _20687_, _20685_);
  not _71829_ (_20688_, \oc8051_golden_model_1.TL1 [2]);
  nor _71830_ (_20689_, _05242_, _20688_);
  nor _71831_ (_20690_, _12400_, _09205_);
  nor _71832_ (_20691_, _20690_, _20689_);
  nor _71833_ (_20692_, _20691_, _04517_);
  and _71834_ (_20693_, _05242_, \oc8051_golden_model_1.ACC [2]);
  nor _71835_ (_20694_, _20693_, _20689_);
  nor _71836_ (_20695_, _20694_, _03583_);
  nor _71837_ (_20696_, _20694_, _04427_);
  nor _71838_ (_20697_, _04426_, _20688_);
  or _71839_ (_20698_, _20697_, _20696_);
  and _71840_ (_20699_, _20698_, _04444_);
  nor _71841_ (_20701_, _12282_, _09205_);
  nor _71842_ (_20702_, _20701_, _20689_);
  nor _71843_ (_20703_, _20702_, _04444_);
  or _71844_ (_20704_, _20703_, _20699_);
  and _71845_ (_20705_, _20704_, _03983_);
  nor _71846_ (_20706_, _09205_, _05026_);
  nor _71847_ (_20707_, _20706_, _20689_);
  nor _71848_ (_20708_, _20707_, _03983_);
  nor _71849_ (_20709_, _20708_, _20705_);
  nor _71850_ (_20710_, _20709_, _03575_);
  or _71851_ (_20712_, _20710_, _07314_);
  nor _71852_ (_20713_, _20712_, _20695_);
  and _71853_ (_20714_, _20707_, _07314_);
  nor _71854_ (_20715_, _20714_, _20713_);
  nor _71855_ (_20716_, _20715_, _03479_);
  nor _71856_ (_20717_, _20689_, _06044_);
  or _71857_ (_20718_, _06569_, _09205_);
  and _71858_ (_20719_, _20718_, _20717_);
  nor _71859_ (_20720_, _20719_, _20716_);
  nor _71860_ (_20721_, _20720_, _03221_);
  or _71861_ (_20722_, _12384_, _09205_);
  nor _71862_ (_20723_, _20689_, _03474_);
  and _71863_ (_20724_, _20723_, _20722_);
  or _71864_ (_20725_, _20724_, _03437_);
  nor _71865_ (_20726_, _20725_, _20721_);
  and _71866_ (_20727_, _05242_, _06261_);
  nor _71867_ (_20728_, _20727_, _20689_);
  nor _71868_ (_20729_, _20728_, _03438_);
  or _71869_ (_20730_, _20729_, _20726_);
  and _71870_ (_20731_, _20730_, _04499_);
  and _71871_ (_20733_, _12273_, _05242_);
  nor _71872_ (_20734_, _20733_, _20689_);
  nor _71873_ (_20735_, _20734_, _04499_);
  or _71874_ (_20736_, _20735_, _20731_);
  nor _71875_ (_20737_, _20736_, _03769_);
  nand _71876_ (_20738_, _12401_, _05444_);
  nor _71877_ (_20739_, _20689_, _04501_);
  and _71878_ (_20740_, _20739_, _20738_);
  or _71879_ (_20741_, _20740_, _04504_);
  nor _71880_ (_20742_, _20741_, _20737_);
  nor _71881_ (_20744_, _20689_, _05665_);
  or _71882_ (_20745_, _20728_, _04505_);
  nor _71883_ (_20746_, _20745_, _20744_);
  nor _71884_ (_20747_, _20746_, _20742_);
  nor _71885_ (_20748_, _20747_, _03752_);
  or _71886_ (_20749_, _20744_, _03753_);
  or _71887_ (_20750_, _20749_, _20694_);
  and _71888_ (_20751_, _20750_, _03759_);
  not _71889_ (_20752_, _20751_);
  nor _71890_ (_20753_, _20752_, _20748_);
  or _71891_ (_20755_, _12272_, _09205_);
  nor _71892_ (_20756_, _20689_, _03759_);
  and _71893_ (_20757_, _20756_, _20755_);
  or _71894_ (_20758_, _20757_, _03760_);
  nor _71895_ (_20759_, _20758_, _20753_);
  nor _71896_ (_20760_, _20759_, _20692_);
  nor _71897_ (_20761_, _20760_, _03790_);
  nor _71898_ (_20762_, _20702_, _04192_);
  or _71899_ (_20763_, _20762_, _03520_);
  nor _71900_ (_20764_, _20763_, _20761_);
  nand _71901_ (_20765_, _12456_, _05444_);
  nor _71902_ (_20766_, _20689_, _03521_);
  and _71903_ (_20767_, _20766_, _20765_);
  nor _71904_ (_20768_, _20767_, _20764_);
  or _71905_ (_20769_, _20768_, _42967_);
  or _71906_ (_20770_, _42963_, \oc8051_golden_model_1.TL1 [2]);
  and _71907_ (_20771_, _20770_, _41755_);
  and _71908_ (_43257_, _20771_, _20769_);
  not _71909_ (_20772_, \oc8051_golden_model_1.TL1 [3]);
  nor _71910_ (_20773_, _05242_, _20772_);
  and _71911_ (_20775_, _06717_, _05242_);
  nor _71912_ (_20776_, _20775_, _20773_);
  or _71913_ (_20777_, _20776_, _06044_);
  and _71914_ (_20778_, _05242_, \oc8051_golden_model_1.ACC [3]);
  nor _71915_ (_20779_, _20778_, _20773_);
  nor _71916_ (_20780_, _20779_, _04427_);
  nor _71917_ (_20781_, _04426_, _20772_);
  or _71918_ (_20782_, _20781_, _20780_);
  and _71919_ (_20783_, _20782_, _04444_);
  nor _71920_ (_20784_, _12486_, _09205_);
  nor _71921_ (_20786_, _20784_, _20773_);
  nor _71922_ (_20787_, _20786_, _04444_);
  or _71923_ (_20788_, _20787_, _20783_);
  and _71924_ (_20789_, _20788_, _03983_);
  nor _71925_ (_20790_, _09205_, _04843_);
  nor _71926_ (_20791_, _20790_, _20773_);
  nor _71927_ (_20792_, _20791_, _03983_);
  nor _71928_ (_20793_, _20792_, _20789_);
  nor _71929_ (_20794_, _20793_, _03575_);
  nor _71930_ (_20795_, _20779_, _03583_);
  nor _71931_ (_20796_, _20795_, _07314_);
  not _71932_ (_20797_, _20796_);
  nor _71933_ (_20798_, _20797_, _20794_);
  and _71934_ (_20799_, _20791_, _07314_);
  or _71935_ (_20800_, _20799_, _03479_);
  or _71936_ (_20801_, _20800_, _20798_);
  and _71937_ (_20802_, _20801_, _03474_);
  and _71938_ (_20803_, _20802_, _20777_);
  or _71939_ (_20804_, _12583_, _09205_);
  nor _71940_ (_20805_, _20773_, _03474_);
  and _71941_ (_20807_, _20805_, _20804_);
  or _71942_ (_20808_, _20807_, _03437_);
  nor _71943_ (_20809_, _20808_, _20803_);
  and _71944_ (_20810_, _05242_, _06217_);
  nor _71945_ (_20811_, _20810_, _20773_);
  nor _71946_ (_20812_, _20811_, _03438_);
  or _71947_ (_20813_, _20812_, _20809_);
  and _71948_ (_20814_, _20813_, _04499_);
  and _71949_ (_20815_, _12598_, _05242_);
  nor _71950_ (_20816_, _20815_, _20773_);
  nor _71951_ (_20818_, _20816_, _04499_);
  or _71952_ (_20819_, _20818_, _20814_);
  nor _71953_ (_20820_, _20819_, _03769_);
  nand _71954_ (_20821_, _12604_, _05444_);
  nor _71955_ (_20822_, _20773_, _04501_);
  and _71956_ (_20823_, _20822_, _20821_);
  or _71957_ (_20824_, _20823_, _04504_);
  nor _71958_ (_20825_, _20824_, _20820_);
  nor _71959_ (_20826_, _20773_, _05521_);
  or _71960_ (_20827_, _20811_, _04505_);
  nor _71961_ (_20829_, _20827_, _20826_);
  nor _71962_ (_20830_, _20829_, _20825_);
  nor _71963_ (_20831_, _20830_, _03752_);
  or _71964_ (_20832_, _20826_, _03753_);
  or _71965_ (_20833_, _20832_, _20779_);
  and _71966_ (_20834_, _20833_, _03759_);
  not _71967_ (_20835_, _20834_);
  nor _71968_ (_20836_, _20835_, _20831_);
  or _71969_ (_20837_, _12597_, _09205_);
  nor _71970_ (_20838_, _20773_, _03759_);
  and _71971_ (_20839_, _20838_, _20837_);
  or _71972_ (_20840_, _20839_, _03760_);
  nor _71973_ (_20841_, _20840_, _20836_);
  nor _71974_ (_20842_, _12603_, _09205_);
  nor _71975_ (_20843_, _20842_, _20773_);
  nor _71976_ (_20844_, _20843_, _04517_);
  or _71977_ (_20845_, _20844_, _03790_);
  nor _71978_ (_20846_, _20845_, _20841_);
  and _71979_ (_20847_, _20786_, _03790_);
  or _71980_ (_20848_, _20847_, _03520_);
  nor _71981_ (_20850_, _20848_, _20846_);
  and _71982_ (_20851_, _12658_, _05242_);
  nor _71983_ (_20852_, _20851_, _20773_);
  nor _71984_ (_20853_, _20852_, _03521_);
  or _71985_ (_20854_, _20853_, _20850_);
  or _71986_ (_20855_, _20854_, _42967_);
  or _71987_ (_20856_, _42963_, \oc8051_golden_model_1.TL1 [3]);
  and _71988_ (_20857_, _20856_, _41755_);
  and _71989_ (_43258_, _20857_, _20855_);
  not _71990_ (_20858_, \oc8051_golden_model_1.TL1 [4]);
  nor _71991_ (_20860_, _05242_, _20858_);
  and _71992_ (_20861_, _12844_, _05444_);
  nor _71993_ (_20862_, _20861_, _20860_);
  nor _71994_ (_20863_, _20862_, _04501_);
  and _71995_ (_20864_, _05242_, \oc8051_golden_model_1.ACC [4]);
  nor _71996_ (_20865_, _20864_, _20860_);
  nor _71997_ (_20866_, _20865_, _04427_);
  nor _71998_ (_20867_, _04426_, _20858_);
  or _71999_ (_20868_, _20867_, _20866_);
  and _72000_ (_20869_, _20868_, _04444_);
  nor _72001_ (_20870_, _12733_, _09205_);
  nor _72002_ (_20871_, _20870_, _20860_);
  nor _72003_ (_20872_, _20871_, _04444_);
  or _72004_ (_20873_, _20872_, _20869_);
  and _72005_ (_20874_, _20873_, _03983_);
  nor _72006_ (_20875_, _05712_, _09205_);
  nor _72007_ (_20876_, _20875_, _20860_);
  nor _72008_ (_20877_, _20876_, _03983_);
  nor _72009_ (_20878_, _20877_, _20874_);
  nor _72010_ (_20879_, _20878_, _03575_);
  nor _72011_ (_20881_, _20865_, _03583_);
  nor _72012_ (_20882_, _20881_, _07314_);
  not _72013_ (_20883_, _20882_);
  nor _72014_ (_20884_, _20883_, _20879_);
  and _72015_ (_20885_, _20876_, _07314_);
  or _72016_ (_20886_, _20885_, _03479_);
  nor _72017_ (_20887_, _20886_, _20884_);
  and _72018_ (_20888_, _06722_, _05242_);
  or _72019_ (_20889_, _20888_, _20860_);
  and _72020_ (_20890_, _20889_, _03479_);
  or _72021_ (_20892_, _20890_, _03221_);
  or _72022_ (_20893_, _20892_, _20887_);
  nor _72023_ (_20894_, _12827_, _09205_);
  or _72024_ (_20895_, _20860_, _03474_);
  or _72025_ (_20896_, _20895_, _20894_);
  and _72026_ (_20897_, _20896_, _03438_);
  and _72027_ (_20898_, _20897_, _20893_);
  and _72028_ (_20899_, _06233_, _05242_);
  nor _72029_ (_20900_, _20899_, _20860_);
  nor _72030_ (_20901_, _20900_, _03438_);
  or _72031_ (_20903_, _20901_, _03636_);
  nor _72032_ (_20904_, _20903_, _20898_);
  nand _72033_ (_20905_, _12711_, _05444_);
  nor _72034_ (_20906_, _20860_, _04499_);
  and _72035_ (_20907_, _20906_, _20905_);
  or _72036_ (_20908_, _20907_, _03769_);
  nor _72037_ (_20909_, _20908_, _20904_);
  nor _72038_ (_20910_, _20909_, _20863_);
  nor _72039_ (_20911_, _20910_, _04504_);
  not _72040_ (_20912_, _20860_);
  and _72041_ (_20914_, _20912_, _05760_);
  or _72042_ (_20915_, _20900_, _04505_);
  nor _72043_ (_20916_, _20915_, _20914_);
  nor _72044_ (_20917_, _20916_, _20911_);
  nor _72045_ (_20918_, _20917_, _03752_);
  or _72046_ (_20919_, _20914_, _03753_);
  or _72047_ (_20920_, _20919_, _20865_);
  and _72048_ (_20921_, _20920_, _03759_);
  not _72049_ (_20922_, _20921_);
  nor _72050_ (_20923_, _20922_, _20918_);
  or _72051_ (_20925_, _12710_, _09205_);
  nor _72052_ (_20926_, _20860_, _03759_);
  and _72053_ (_20927_, _20926_, _20925_);
  or _72054_ (_20928_, _20927_, _03760_);
  nor _72055_ (_20929_, _20928_, _20923_);
  nor _72056_ (_20930_, _12843_, _09205_);
  nor _72057_ (_20931_, _20930_, _20860_);
  nor _72058_ (_20932_, _20931_, _04517_);
  or _72059_ (_20933_, _20932_, _03790_);
  nor _72060_ (_20934_, _20933_, _20929_);
  and _72061_ (_20936_, _20871_, _03790_);
  or _72062_ (_20937_, _20936_, _03520_);
  nor _72063_ (_20938_, _20937_, _20934_);
  and _72064_ (_20939_, _12893_, _05242_);
  nor _72065_ (_20940_, _20939_, _20860_);
  nor _72066_ (_20941_, _20940_, _03521_);
  or _72067_ (_20942_, _20941_, _20938_);
  or _72068_ (_20943_, _20942_, _42967_);
  or _72069_ (_20944_, _42963_, \oc8051_golden_model_1.TL1 [4]);
  and _72070_ (_20945_, _20944_, _41755_);
  and _72071_ (_43259_, _20945_, _20943_);
  not _72072_ (_20947_, \oc8051_golden_model_1.TL1 [5]);
  nor _72073_ (_20948_, _05242_, _20947_);
  and _72074_ (_20949_, _13042_, _05444_);
  nor _72075_ (_20950_, _20949_, _20948_);
  nor _72076_ (_20951_, _20950_, _04501_);
  nor _72077_ (_20952_, _05422_, _09205_);
  nor _72078_ (_20953_, _20952_, _20948_);
  and _72079_ (_20954_, _20953_, _07314_);
  and _72080_ (_20955_, _05242_, \oc8051_golden_model_1.ACC [5]);
  nor _72081_ (_20957_, _20955_, _20948_);
  nor _72082_ (_20958_, _20957_, _04427_);
  nor _72083_ (_20959_, _04426_, _20947_);
  or _72084_ (_20960_, _20959_, _20958_);
  and _72085_ (_20961_, _20960_, _04444_);
  nor _72086_ (_20962_, _12930_, _09205_);
  nor _72087_ (_20963_, _20962_, _20948_);
  nor _72088_ (_20964_, _20963_, _04444_);
  or _72089_ (_20965_, _20964_, _20961_);
  and _72090_ (_20966_, _20965_, _03983_);
  nor _72091_ (_20968_, _20953_, _03983_);
  nor _72092_ (_20969_, _20968_, _20966_);
  nor _72093_ (_20970_, _20969_, _03575_);
  nor _72094_ (_20971_, _20957_, _03583_);
  nor _72095_ (_20972_, _20971_, _07314_);
  not _72096_ (_20973_, _20972_);
  nor _72097_ (_20974_, _20973_, _20970_);
  nor _72098_ (_20975_, _20974_, _20954_);
  nor _72099_ (_20976_, _20975_, _03479_);
  nor _72100_ (_20977_, _20948_, _06044_);
  or _72101_ (_20978_, _06616_, _09229_);
  and _72102_ (_20979_, _20978_, _20977_);
  or _72103_ (_20980_, _20979_, _03221_);
  nor _72104_ (_20981_, _20980_, _20976_);
  nor _72105_ (_20982_, _13021_, _09229_);
  nor _72106_ (_20983_, _20982_, _20948_);
  nor _72107_ (_20984_, _20983_, _03474_);
  or _72108_ (_20985_, _20984_, _03437_);
  or _72109_ (_20986_, _20985_, _20981_);
  and _72110_ (_20987_, _06211_, _05242_);
  nor _72111_ (_20988_, _20987_, _20948_);
  nand _72112_ (_20989_, _20988_, _03437_);
  and _72113_ (_20990_, _20989_, _20986_);
  nor _72114_ (_20991_, _20990_, _03636_);
  nand _72115_ (_20992_, _13036_, _05444_);
  nor _72116_ (_20993_, _20948_, _04499_);
  and _72117_ (_20994_, _20993_, _20992_);
  or _72118_ (_20995_, _20994_, _03769_);
  nor _72119_ (_20996_, _20995_, _20991_);
  nor _72120_ (_20997_, _20996_, _20951_);
  nor _72121_ (_20999_, _20997_, _04504_);
  not _72122_ (_21000_, _20948_);
  and _72123_ (_21001_, _21000_, _05471_);
  or _72124_ (_21002_, _20988_, _04505_);
  nor _72125_ (_21003_, _21002_, _21001_);
  nor _72126_ (_21004_, _21003_, _20999_);
  nor _72127_ (_21005_, _21004_, _03752_);
  or _72128_ (_21006_, _21001_, _03753_);
  or _72129_ (_21007_, _21006_, _20957_);
  and _72130_ (_21008_, _21007_, _03759_);
  not _72131_ (_21010_, _21008_);
  nor _72132_ (_21011_, _21010_, _21005_);
  or _72133_ (_21012_, _13035_, _09205_);
  nor _72134_ (_21013_, _20948_, _03759_);
  and _72135_ (_21014_, _21013_, _21012_);
  or _72136_ (_21015_, _21014_, _03760_);
  nor _72137_ (_21016_, _21015_, _21011_);
  nor _72138_ (_21017_, _13041_, _09205_);
  nor _72139_ (_21018_, _21017_, _20948_);
  nor _72140_ (_21019_, _21018_, _04517_);
  or _72141_ (_21021_, _21019_, _03790_);
  nor _72142_ (_21022_, _21021_, _21016_);
  and _72143_ (_21023_, _20963_, _03790_);
  or _72144_ (_21024_, _21023_, _03520_);
  nor _72145_ (_21025_, _21024_, _21022_);
  and _72146_ (_21026_, _13097_, _05242_);
  nor _72147_ (_21027_, _21026_, _20948_);
  nor _72148_ (_21028_, _21027_, _03521_);
  or _72149_ (_21029_, _21028_, _21025_);
  or _72150_ (_21030_, _21029_, _42967_);
  or _72151_ (_21032_, _42963_, \oc8051_golden_model_1.TL1 [5]);
  and _72152_ (_21033_, _21032_, _41755_);
  and _72153_ (_43262_, _21033_, _21030_);
  not _72154_ (_21034_, \oc8051_golden_model_1.TL1 [6]);
  nor _72155_ (_21035_, _05242_, _21034_);
  and _72156_ (_21036_, _13259_, _05444_);
  nor _72157_ (_21037_, _21036_, _21035_);
  nor _72158_ (_21038_, _21037_, _04501_);
  nor _72159_ (_21039_, _05327_, _09205_);
  nor _72160_ (_21040_, _21039_, _21035_);
  and _72161_ (_21042_, _21040_, _07314_);
  and _72162_ (_21043_, _05242_, \oc8051_golden_model_1.ACC [6]);
  nor _72163_ (_21044_, _21043_, _21035_);
  nor _72164_ (_21045_, _21044_, _04427_);
  nor _72165_ (_21046_, _04426_, _21034_);
  or _72166_ (_21047_, _21046_, _21045_);
  and _72167_ (_21048_, _21047_, _04444_);
  nor _72168_ (_21049_, _13122_, _09205_);
  nor _72169_ (_21050_, _21049_, _21035_);
  nor _72170_ (_21051_, _21050_, _04444_);
  or _72171_ (_21053_, _21051_, _21048_);
  and _72172_ (_21054_, _21053_, _03983_);
  nor _72173_ (_21055_, _21040_, _03983_);
  nor _72174_ (_21056_, _21055_, _21054_);
  nor _72175_ (_21057_, _21056_, _03575_);
  nor _72176_ (_21058_, _21044_, _03583_);
  nor _72177_ (_21059_, _21058_, _07314_);
  not _72178_ (_21060_, _21059_);
  nor _72179_ (_21061_, _21060_, _21057_);
  nor _72180_ (_21062_, _21061_, _21042_);
  nor _72181_ (_21064_, _21062_, _03479_);
  nor _72182_ (_21065_, _21035_, _06044_);
  or _72183_ (_21066_, _06388_, _09229_);
  and _72184_ (_21067_, _21066_, _21065_);
  or _72185_ (_21068_, _21067_, _03221_);
  nor _72186_ (_21069_, _21068_, _21064_);
  nor _72187_ (_21070_, _13237_, _09229_);
  nor _72188_ (_21071_, _21070_, _21035_);
  nor _72189_ (_21072_, _21071_, _03474_);
  or _72190_ (_21073_, _21072_, _03437_);
  or _72191_ (_21075_, _21073_, _21069_);
  and _72192_ (_21076_, _13244_, _05242_);
  nor _72193_ (_21077_, _21076_, _21035_);
  nand _72194_ (_21078_, _21077_, _03437_);
  and _72195_ (_21079_, _21078_, _21075_);
  nor _72196_ (_21080_, _21079_, _03636_);
  nand _72197_ (_21081_, _13253_, _05444_);
  nor _72198_ (_21082_, _21035_, _04499_);
  and _72199_ (_21083_, _21082_, _21081_);
  or _72200_ (_21084_, _21083_, _03769_);
  nor _72201_ (_21086_, _21084_, _21080_);
  nor _72202_ (_21087_, _21086_, _21038_);
  nor _72203_ (_21088_, _21087_, _04504_);
  not _72204_ (_21089_, _21035_);
  and _72205_ (_21090_, _21089_, _05376_);
  or _72206_ (_21091_, _21077_, _04505_);
  nor _72207_ (_21092_, _21091_, _21090_);
  nor _72208_ (_21093_, _21092_, _21088_);
  nor _72209_ (_21094_, _21093_, _03752_);
  or _72210_ (_21095_, _21090_, _03753_);
  nor _72211_ (_21097_, _21095_, _21044_);
  or _72212_ (_21098_, _21097_, _21094_);
  and _72213_ (_21099_, _21098_, _03759_);
  nor _72214_ (_21100_, _13251_, _09229_);
  nor _72215_ (_21101_, _21100_, _21035_);
  nor _72216_ (_21102_, _21101_, _03759_);
  or _72217_ (_21103_, _21102_, _21099_);
  and _72218_ (_21104_, _21103_, _04517_);
  nor _72219_ (_21105_, _13258_, _09205_);
  nor _72220_ (_21106_, _21105_, _21035_);
  nor _72221_ (_21108_, _21106_, _04517_);
  or _72222_ (_21109_, _21108_, _03790_);
  nor _72223_ (_21110_, _21109_, _21104_);
  and _72224_ (_21111_, _21050_, _03790_);
  or _72225_ (_21112_, _21111_, _03520_);
  nor _72226_ (_21113_, _21112_, _21110_);
  and _72227_ (_21114_, _13312_, _05242_);
  nor _72228_ (_21115_, _21114_, _21035_);
  nor _72229_ (_21116_, _21115_, _03521_);
  or _72230_ (_21117_, _21116_, _21113_);
  or _72231_ (_21119_, _21117_, _42967_);
  or _72232_ (_21120_, _42963_, \oc8051_golden_model_1.TL1 [6]);
  and _72233_ (_21121_, _21120_, _41755_);
  and _72234_ (_43263_, _21121_, _21119_);
  not _72235_ (_21122_, \oc8051_golden_model_1.TH0 [0]);
  nor _72236_ (_21123_, _05234_, _21122_);
  and _72237_ (_21124_, _05941_, _05234_);
  nor _72238_ (_21125_, _21124_, _21123_);
  and _72239_ (_21126_, _21125_, _17076_);
  and _72240_ (_21127_, _05234_, \oc8051_golden_model_1.ACC [0]);
  nor _72241_ (_21129_, _21127_, _21123_);
  nor _72242_ (_21130_, _21129_, _03583_);
  nor _72243_ (_21131_, _21130_, _07314_);
  nor _72244_ (_21132_, _21125_, _04444_);
  nor _72245_ (_21133_, _04426_, _21122_);
  nor _72246_ (_21134_, _21129_, _04427_);
  nor _72247_ (_21135_, _21134_, _21133_);
  nor _72248_ (_21136_, _21135_, _03570_);
  or _72249_ (_21137_, _21136_, _03568_);
  nor _72250_ (_21138_, _21137_, _21132_);
  or _72251_ (_21140_, _21138_, _03575_);
  and _72252_ (_21141_, _21140_, _21131_);
  and _72253_ (_21142_, _05234_, _04419_);
  or _72254_ (_21143_, _21123_, _18522_);
  nor _72255_ (_21144_, _21143_, _21142_);
  nor _72256_ (_21145_, _21144_, _21141_);
  nor _72257_ (_21146_, _21145_, _03479_);
  and _72258_ (_21147_, _06715_, _05234_);
  nor _72259_ (_21148_, _21123_, _06044_);
  not _72260_ (_21149_, _21148_);
  nor _72261_ (_21151_, _21149_, _21147_);
  nor _72262_ (_21152_, _21151_, _21146_);
  nor _72263_ (_21153_, _21152_, _03221_);
  nor _72264_ (_21154_, _11975_, _09299_);
  or _72265_ (_21155_, _21123_, _03474_);
  nor _72266_ (_21156_, _21155_, _21154_);
  or _72267_ (_21157_, _21156_, _03437_);
  nor _72268_ (_21158_, _21157_, _21153_);
  and _72269_ (_21159_, _05234_, _06202_);
  nor _72270_ (_21160_, _21159_, _21123_);
  nor _72271_ (_21162_, _21160_, _03438_);
  or _72272_ (_21163_, _21162_, _21158_);
  and _72273_ (_21164_, _21163_, _04499_);
  and _72274_ (_21165_, _11990_, _05234_);
  nor _72275_ (_21166_, _21165_, _21123_);
  nor _72276_ (_21167_, _21166_, _04499_);
  or _72277_ (_21168_, _21167_, _21164_);
  nor _72278_ (_21169_, _21168_, _03769_);
  and _72279_ (_21170_, _11995_, _05234_);
  or _72280_ (_21171_, _21123_, _04501_);
  nor _72281_ (_21173_, _21171_, _21170_);
  or _72282_ (_21174_, _21173_, _04504_);
  nor _72283_ (_21175_, _21174_, _21169_);
  or _72284_ (_21176_, _21160_, _04505_);
  nor _72285_ (_21177_, _21176_, _21124_);
  nor _72286_ (_21178_, _21177_, _21175_);
  nor _72287_ (_21179_, _21178_, _03752_);
  and _72288_ (_21180_, _11994_, _05234_);
  or _72289_ (_21181_, _21180_, _21123_);
  and _72290_ (_21182_, _21181_, _03752_);
  or _72291_ (_21184_, _21182_, _21179_);
  and _72292_ (_21185_, _21184_, _03759_);
  nor _72293_ (_21186_, _11988_, _09299_);
  nor _72294_ (_21187_, _21186_, _21123_);
  nor _72295_ (_21188_, _21187_, _03759_);
  or _72296_ (_21189_, _21188_, _21185_);
  and _72297_ (_21190_, _21189_, _04517_);
  nor _72298_ (_21191_, _11870_, _09299_);
  nor _72299_ (_21192_, _21191_, _21123_);
  nor _72300_ (_21193_, _21192_, _04517_);
  nor _72301_ (_21195_, _21193_, _17076_);
  not _72302_ (_21196_, _21195_);
  nor _72303_ (_21197_, _21196_, _21190_);
  nor _72304_ (_21198_, _21197_, _21126_);
  or _72305_ (_21199_, _21198_, _42967_);
  or _72306_ (_21200_, _42963_, \oc8051_golden_model_1.TH0 [0]);
  and _72307_ (_21201_, _21200_, _41755_);
  and _72308_ (_43264_, _21201_, _21199_);
  nor _72309_ (_21202_, _05234_, \oc8051_golden_model_1.TH0 [1]);
  and _72310_ (_21203_, _12252_, _05234_);
  nor _72311_ (_21205_, _21203_, _21202_);
  nor _72312_ (_21206_, _21205_, _04192_);
  and _72313_ (_21207_, _06714_, _05234_);
  not _72314_ (_21208_, \oc8051_golden_model_1.TH0 [1]);
  nor _72315_ (_21209_, _05234_, _21208_);
  nor _72316_ (_21210_, _21209_, _06044_);
  not _72317_ (_21211_, _21210_);
  nor _72318_ (_21212_, _21211_, _21207_);
  not _72319_ (_21213_, _21212_);
  and _72320_ (_21214_, _05234_, _03233_);
  nor _72321_ (_21216_, _21214_, _21202_);
  and _72322_ (_21217_, _21216_, _03575_);
  nor _72323_ (_21218_, _09299_, _04603_);
  nor _72324_ (_21219_, _21218_, _21209_);
  nor _72325_ (_21220_, _21219_, _03983_);
  and _72326_ (_21221_, _21216_, _04426_);
  nor _72327_ (_21222_, _04426_, _21208_);
  or _72328_ (_21223_, _21222_, _21221_);
  and _72329_ (_21224_, _21223_, _04444_);
  and _72330_ (_21225_, _21205_, _03570_);
  or _72331_ (_21227_, _21225_, _21224_);
  and _72332_ (_21228_, _21227_, _03983_);
  nor _72333_ (_21229_, _21228_, _21220_);
  nor _72334_ (_21230_, _21229_, _03575_);
  or _72335_ (_21231_, _21230_, _07314_);
  nor _72336_ (_21232_, _21231_, _21217_);
  and _72337_ (_21233_, _21219_, _07314_);
  nor _72338_ (_21234_, _21233_, _21232_);
  nor _72339_ (_21235_, _21234_, _03479_);
  nor _72340_ (_21236_, _21235_, _03221_);
  and _72341_ (_21238_, _21236_, _21213_);
  not _72342_ (_21239_, _21202_);
  and _72343_ (_21240_, _12176_, _05234_);
  nor _72344_ (_21241_, _21240_, _03474_);
  and _72345_ (_21242_, _21241_, _21239_);
  nor _72346_ (_21243_, _21242_, _21238_);
  nor _72347_ (_21244_, _21243_, _03437_);
  and _72348_ (_21245_, _05234_, _04317_);
  not _72349_ (_21246_, _21245_);
  nor _72350_ (_21247_, _21202_, _03438_);
  and _72351_ (_21249_, _21247_, _21246_);
  nor _72352_ (_21250_, _21249_, _21244_);
  nor _72353_ (_21251_, _21250_, _03636_);
  nor _72354_ (_21252_, _12191_, _09299_);
  nor _72355_ (_21253_, _21252_, _04499_);
  and _72356_ (_21254_, _21253_, _21239_);
  nor _72357_ (_21255_, _21254_, _21251_);
  nor _72358_ (_21256_, _21255_, _03769_);
  nor _72359_ (_21257_, _12197_, _09299_);
  nor _72360_ (_21258_, _21257_, _04501_);
  and _72361_ (_21260_, _21258_, _21239_);
  nor _72362_ (_21261_, _21260_, _21256_);
  nor _72363_ (_21262_, _21261_, _04504_);
  nor _72364_ (_21263_, _12190_, _09299_);
  nor _72365_ (_21264_, _21263_, _05769_);
  and _72366_ (_21265_, _21264_, _21239_);
  nor _72367_ (_21266_, _21265_, _21262_);
  nor _72368_ (_21267_, _21266_, _03752_);
  nor _72369_ (_21268_, _21209_, _05569_);
  nor _72370_ (_21269_, _21268_, _03753_);
  and _72371_ (_21271_, _21269_, _21216_);
  nor _72372_ (_21272_, _21271_, _21267_);
  nor _72373_ (_21273_, _21272_, _03758_);
  and _72374_ (_21274_, _21245_, _05940_);
  nor _72375_ (_21275_, _21274_, _03759_);
  and _72376_ (_21276_, _21275_, _21239_);
  nor _72377_ (_21277_, _21276_, _21273_);
  nor _72378_ (_21278_, _21277_, _03760_);
  nand _72379_ (_21279_, _21214_, _05940_);
  nor _72380_ (_21280_, _21202_, _04517_);
  and _72381_ (_21282_, _21280_, _21279_);
  or _72382_ (_21283_, _21282_, _03790_);
  nor _72383_ (_21284_, _21283_, _21278_);
  nor _72384_ (_21285_, _21284_, _21206_);
  and _72385_ (_21286_, _21285_, _03521_);
  nor _72386_ (_21287_, _21209_, _21203_);
  nor _72387_ (_21288_, _21287_, _03521_);
  or _72388_ (_21289_, _21288_, _21286_);
  or _72389_ (_21290_, _21289_, _42967_);
  or _72390_ (_21291_, _42963_, \oc8051_golden_model_1.TH0 [1]);
  and _72391_ (_21293_, _21291_, _41755_);
  and _72392_ (_43265_, _21293_, _21290_);
  not _72393_ (_21294_, \oc8051_golden_model_1.TH0 [2]);
  nor _72394_ (_21295_, _05234_, _21294_);
  nor _72395_ (_21296_, _12400_, _09299_);
  nor _72396_ (_21297_, _21296_, _21295_);
  nor _72397_ (_21298_, _21297_, _04517_);
  and _72398_ (_21299_, _05234_, \oc8051_golden_model_1.ACC [2]);
  nor _72399_ (_21300_, _21299_, _21295_);
  nor _72400_ (_21301_, _21300_, _03583_);
  nor _72401_ (_21303_, _21300_, _04427_);
  nor _72402_ (_21304_, _04426_, _21294_);
  or _72403_ (_21305_, _21304_, _21303_);
  and _72404_ (_21306_, _21305_, _04444_);
  nor _72405_ (_21307_, _12282_, _09299_);
  nor _72406_ (_21308_, _21307_, _21295_);
  nor _72407_ (_21309_, _21308_, _04444_);
  or _72408_ (_21310_, _21309_, _21306_);
  and _72409_ (_21311_, _21310_, _03983_);
  nor _72410_ (_21312_, _09299_, _05026_);
  nor _72411_ (_21314_, _21312_, _21295_);
  nor _72412_ (_21315_, _21314_, _03983_);
  nor _72413_ (_21316_, _21315_, _21311_);
  nor _72414_ (_21317_, _21316_, _03575_);
  or _72415_ (_21318_, _21317_, _07314_);
  nor _72416_ (_21319_, _21318_, _21301_);
  and _72417_ (_21320_, _21314_, _07314_);
  nor _72418_ (_21321_, _21320_, _21319_);
  nor _72419_ (_21322_, _21321_, _03479_);
  and _72420_ (_21323_, _06718_, _05234_);
  nor _72421_ (_21325_, _21295_, _06044_);
  not _72422_ (_21326_, _21325_);
  nor _72423_ (_21327_, _21326_, _21323_);
  nor _72424_ (_21328_, _21327_, _21322_);
  nor _72425_ (_21329_, _21328_, _03221_);
  nor _72426_ (_21330_, _12384_, _09299_);
  or _72427_ (_21331_, _21295_, _03474_);
  nor _72428_ (_21332_, _21331_, _21330_);
  or _72429_ (_21333_, _21332_, _03437_);
  nor _72430_ (_21334_, _21333_, _21329_);
  and _72431_ (_21336_, _05234_, _06261_);
  nor _72432_ (_21337_, _21336_, _21295_);
  nor _72433_ (_21338_, _21337_, _03438_);
  or _72434_ (_21339_, _21338_, _21334_);
  and _72435_ (_21340_, _21339_, _04499_);
  and _72436_ (_21341_, _12273_, _05234_);
  nor _72437_ (_21342_, _21341_, _21295_);
  nor _72438_ (_21343_, _21342_, _04499_);
  or _72439_ (_21344_, _21343_, _21340_);
  nor _72440_ (_21345_, _21344_, _03769_);
  and _72441_ (_21347_, _12401_, _05234_);
  or _72442_ (_21348_, _21295_, _04501_);
  nor _72443_ (_21349_, _21348_, _21347_);
  or _72444_ (_21350_, _21349_, _04504_);
  nor _72445_ (_21351_, _21350_, _21345_);
  nor _72446_ (_21352_, _21295_, _05665_);
  or _72447_ (_21353_, _21337_, _04505_);
  nor _72448_ (_21354_, _21353_, _21352_);
  nor _72449_ (_21355_, _21354_, _21351_);
  nor _72450_ (_21356_, _21355_, _03752_);
  or _72451_ (_21358_, _21352_, _03753_);
  nor _72452_ (_21359_, _21358_, _21300_);
  or _72453_ (_21360_, _21359_, _21356_);
  and _72454_ (_21361_, _21360_, _03759_);
  nor _72455_ (_21362_, _12272_, _09299_);
  nor _72456_ (_21363_, _21362_, _21295_);
  nor _72457_ (_21364_, _21363_, _03759_);
  or _72458_ (_21365_, _21364_, _21361_);
  and _72459_ (_21366_, _21365_, _04517_);
  nor _72460_ (_21367_, _21366_, _21298_);
  nor _72461_ (_21369_, _21367_, _03790_);
  nor _72462_ (_21370_, _21308_, _04192_);
  or _72463_ (_21371_, _21370_, _03520_);
  nor _72464_ (_21372_, _21371_, _21369_);
  and _72465_ (_21373_, _12456_, _05234_);
  or _72466_ (_21374_, _21295_, _03521_);
  nor _72467_ (_21375_, _21374_, _21373_);
  nor _72468_ (_21376_, _21375_, _21372_);
  or _72469_ (_21377_, _21376_, _42967_);
  or _72470_ (_21378_, _42963_, \oc8051_golden_model_1.TH0 [2]);
  and _72471_ (_21380_, _21378_, _41755_);
  and _72472_ (_43266_, _21380_, _21377_);
  not _72473_ (_21381_, \oc8051_golden_model_1.TH0 [3]);
  nor _72474_ (_21382_, _05234_, _21381_);
  and _72475_ (_21383_, _12604_, _05234_);
  nor _72476_ (_21384_, _21383_, _21382_);
  nor _72477_ (_21385_, _21384_, _04501_);
  and _72478_ (_21386_, _05234_, \oc8051_golden_model_1.ACC [3]);
  nor _72479_ (_21387_, _21386_, _21382_);
  nor _72480_ (_21388_, _21387_, _03583_);
  nor _72481_ (_21390_, _21387_, _04427_);
  nor _72482_ (_21391_, _04426_, _21381_);
  or _72483_ (_21392_, _21391_, _21390_);
  and _72484_ (_21393_, _21392_, _04444_);
  nor _72485_ (_21394_, _12486_, _09299_);
  nor _72486_ (_21395_, _21394_, _21382_);
  nor _72487_ (_21396_, _21395_, _04444_);
  or _72488_ (_21397_, _21396_, _21393_);
  and _72489_ (_21398_, _21397_, _03983_);
  nor _72490_ (_21399_, _09299_, _04843_);
  nor _72491_ (_21401_, _21399_, _21382_);
  nor _72492_ (_21402_, _21401_, _03983_);
  nor _72493_ (_21403_, _21402_, _21398_);
  nor _72494_ (_21404_, _21403_, _03575_);
  or _72495_ (_21405_, _21404_, _07314_);
  nor _72496_ (_21406_, _21405_, _21388_);
  and _72497_ (_21407_, _21401_, _07314_);
  nor _72498_ (_21408_, _21407_, _21406_);
  nor _72499_ (_21409_, _21408_, _03479_);
  and _72500_ (_21410_, _06717_, _05234_);
  nor _72501_ (_21412_, _21382_, _06044_);
  not _72502_ (_21413_, _21412_);
  nor _72503_ (_21414_, _21413_, _21410_);
  or _72504_ (_21415_, _21414_, _03221_);
  nor _72505_ (_21416_, _21415_, _21409_);
  nor _72506_ (_21417_, _12583_, _09299_);
  nor _72507_ (_21418_, _21417_, _21382_);
  nor _72508_ (_21419_, _21418_, _03474_);
  or _72509_ (_21420_, _21419_, _03437_);
  or _72510_ (_21421_, _21420_, _21416_);
  and _72511_ (_21423_, _05234_, _06217_);
  nor _72512_ (_21424_, _21423_, _21382_);
  nand _72513_ (_21425_, _21424_, _03437_);
  and _72514_ (_21426_, _21425_, _21421_);
  nor _72515_ (_21427_, _21426_, _03636_);
  and _72516_ (_21428_, _12598_, _05234_);
  or _72517_ (_21429_, _21382_, _04499_);
  nor _72518_ (_21430_, _21429_, _21428_);
  or _72519_ (_21431_, _21430_, _03769_);
  nor _72520_ (_21432_, _21431_, _21427_);
  nor _72521_ (_21434_, _21432_, _21385_);
  nor _72522_ (_21435_, _21434_, _04504_);
  not _72523_ (_21436_, _21382_);
  and _72524_ (_21437_, _21436_, _05520_);
  or _72525_ (_21438_, _21424_, _04505_);
  nor _72526_ (_21439_, _21438_, _21437_);
  nor _72527_ (_21440_, _21439_, _21435_);
  nor _72528_ (_21441_, _21440_, _03752_);
  or _72529_ (_21442_, _21437_, _03753_);
  or _72530_ (_21443_, _21442_, _21387_);
  and _72531_ (_21445_, _21443_, _03759_);
  not _72532_ (_21446_, _21445_);
  nor _72533_ (_21447_, _21446_, _21441_);
  nor _72534_ (_21448_, _12597_, _09299_);
  or _72535_ (_21449_, _21382_, _03759_);
  nor _72536_ (_21450_, _21449_, _21448_);
  or _72537_ (_21451_, _21450_, _03760_);
  nor _72538_ (_21452_, _21451_, _21447_);
  nor _72539_ (_21453_, _12603_, _09299_);
  nor _72540_ (_21454_, _21453_, _21382_);
  nor _72541_ (_21456_, _21454_, _04517_);
  or _72542_ (_21457_, _21456_, _03790_);
  nor _72543_ (_21458_, _21457_, _21452_);
  and _72544_ (_21459_, _21395_, _03790_);
  or _72545_ (_21460_, _21459_, _03520_);
  nor _72546_ (_21461_, _21460_, _21458_);
  and _72547_ (_21462_, _12658_, _05234_);
  nor _72548_ (_21463_, _21462_, _21382_);
  nor _72549_ (_21464_, _21463_, _03521_);
  or _72550_ (_21465_, _21464_, _21461_);
  or _72551_ (_21467_, _21465_, _42967_);
  or _72552_ (_21468_, _42963_, \oc8051_golden_model_1.TH0 [3]);
  and _72553_ (_21469_, _21468_, _41755_);
  and _72554_ (_43267_, _21469_, _21467_);
  not _72555_ (_21470_, \oc8051_golden_model_1.TH0 [4]);
  nor _72556_ (_21471_, _05234_, _21470_);
  and _72557_ (_21472_, _12844_, _05234_);
  nor _72558_ (_21473_, _21472_, _21471_);
  nor _72559_ (_21474_, _21473_, _04501_);
  and _72560_ (_21475_, _05234_, \oc8051_golden_model_1.ACC [4]);
  nor _72561_ (_21477_, _21475_, _21471_);
  nor _72562_ (_21478_, _21477_, _03583_);
  nor _72563_ (_21479_, _21477_, _04427_);
  nor _72564_ (_21480_, _04426_, _21470_);
  or _72565_ (_21481_, _21480_, _21479_);
  and _72566_ (_21482_, _21481_, _04444_);
  nor _72567_ (_21483_, _12733_, _09299_);
  nor _72568_ (_21484_, _21483_, _21471_);
  nor _72569_ (_21485_, _21484_, _04444_);
  or _72570_ (_21486_, _21485_, _21482_);
  and _72571_ (_21488_, _21486_, _03983_);
  nor _72572_ (_21489_, _05712_, _09299_);
  nor _72573_ (_21490_, _21489_, _21471_);
  nor _72574_ (_21491_, _21490_, _03983_);
  nor _72575_ (_21492_, _21491_, _21488_);
  nor _72576_ (_21493_, _21492_, _03575_);
  or _72577_ (_21494_, _21493_, _07314_);
  nor _72578_ (_21495_, _21494_, _21478_);
  and _72579_ (_21496_, _21490_, _07314_);
  or _72580_ (_21497_, _21496_, _03479_);
  nor _72581_ (_21500_, _21497_, _21495_);
  and _72582_ (_21501_, _06722_, _05234_);
  or _72583_ (_21502_, _21501_, _21471_);
  and _72584_ (_21503_, _21502_, _03479_);
  or _72585_ (_21504_, _21503_, _03221_);
  or _72586_ (_21505_, _21504_, _21500_);
  nor _72587_ (_21506_, _12827_, _09299_);
  or _72588_ (_21507_, _21471_, _03474_);
  or _72589_ (_21508_, _21507_, _21506_);
  and _72590_ (_21509_, _21508_, _03438_);
  and _72591_ (_21512_, _21509_, _21505_);
  and _72592_ (_21513_, _06233_, _05234_);
  nor _72593_ (_21514_, _21513_, _21471_);
  nor _72594_ (_21515_, _21514_, _03438_);
  or _72595_ (_21516_, _21515_, _03636_);
  nor _72596_ (_21517_, _21516_, _21512_);
  and _72597_ (_21518_, _12711_, _05234_);
  or _72598_ (_21519_, _21471_, _04499_);
  nor _72599_ (_21520_, _21519_, _21518_);
  or _72600_ (_21521_, _21520_, _03769_);
  nor _72601_ (_21524_, _21521_, _21517_);
  nor _72602_ (_21525_, _21524_, _21474_);
  nor _72603_ (_21526_, _21525_, _04504_);
  not _72604_ (_21527_, _21471_);
  and _72605_ (_21528_, _21527_, _05760_);
  or _72606_ (_21529_, _21514_, _04505_);
  nor _72607_ (_21530_, _21529_, _21528_);
  nor _72608_ (_21531_, _21530_, _21526_);
  nor _72609_ (_21532_, _21531_, _03752_);
  or _72610_ (_21533_, _21528_, _03753_);
  or _72611_ (_21536_, _21533_, _21477_);
  and _72612_ (_21537_, _21536_, _03759_);
  not _72613_ (_21538_, _21537_);
  nor _72614_ (_21539_, _21538_, _21532_);
  nor _72615_ (_21540_, _12710_, _09299_);
  or _72616_ (_21541_, _21471_, _03759_);
  nor _72617_ (_21542_, _21541_, _21540_);
  or _72618_ (_21543_, _21542_, _03760_);
  nor _72619_ (_21544_, _21543_, _21539_);
  nor _72620_ (_21545_, _12843_, _09299_);
  nor _72621_ (_21548_, _21545_, _21471_);
  nor _72622_ (_21549_, _21548_, _04517_);
  or _72623_ (_21550_, _21549_, _03790_);
  nor _72624_ (_21551_, _21550_, _21544_);
  and _72625_ (_21552_, _21484_, _03790_);
  or _72626_ (_21553_, _21552_, _03520_);
  nor _72627_ (_21554_, _21553_, _21551_);
  and _72628_ (_21555_, _12893_, _05234_);
  nor _72629_ (_21556_, _21555_, _21471_);
  nor _72630_ (_21557_, _21556_, _03521_);
  or _72631_ (_21560_, _21557_, _21554_);
  or _72632_ (_21561_, _21560_, _42967_);
  or _72633_ (_21562_, _42963_, \oc8051_golden_model_1.TH0 [4]);
  and _72634_ (_21563_, _21562_, _41755_);
  and _72635_ (_43268_, _21563_, _21561_);
  not _72636_ (_21564_, \oc8051_golden_model_1.TH0 [5]);
  nor _72637_ (_21565_, _05234_, _21564_);
  and _72638_ (_21566_, _13042_, _05234_);
  nor _72639_ (_21567_, _21566_, _21565_);
  nor _72640_ (_21568_, _21567_, _04501_);
  and _72641_ (_21570_, _05234_, \oc8051_golden_model_1.ACC [5]);
  nor _72642_ (_21571_, _21570_, _21565_);
  nor _72643_ (_21572_, _21571_, _03583_);
  nor _72644_ (_21573_, _21571_, _04427_);
  nor _72645_ (_21574_, _04426_, _21564_);
  or _72646_ (_21575_, _21574_, _21573_);
  and _72647_ (_21576_, _21575_, _04444_);
  nor _72648_ (_21577_, _12930_, _09299_);
  nor _72649_ (_21578_, _21577_, _21565_);
  nor _72650_ (_21579_, _21578_, _04444_);
  or _72651_ (_21581_, _21579_, _21576_);
  and _72652_ (_21582_, _21581_, _03983_);
  nor _72653_ (_21583_, _05422_, _09299_);
  nor _72654_ (_21584_, _21583_, _21565_);
  nor _72655_ (_21585_, _21584_, _03983_);
  nor _72656_ (_21586_, _21585_, _21582_);
  nor _72657_ (_21587_, _21586_, _03575_);
  or _72658_ (_21588_, _21587_, _07314_);
  nor _72659_ (_21589_, _21588_, _21572_);
  and _72660_ (_21590_, _21584_, _07314_);
  nor _72661_ (_21592_, _21590_, _21589_);
  nor _72662_ (_21593_, _21592_, _03479_);
  and _72663_ (_21594_, _06721_, _05234_);
  nor _72664_ (_21595_, _21565_, _06044_);
  not _72665_ (_21596_, _21595_);
  nor _72666_ (_21597_, _21596_, _21594_);
  or _72667_ (_21598_, _21597_, _03221_);
  nor _72668_ (_21599_, _21598_, _21593_);
  nor _72669_ (_21600_, _13021_, _09299_);
  nor _72670_ (_21601_, _21600_, _21565_);
  nor _72671_ (_21603_, _21601_, _03474_);
  or _72672_ (_21604_, _21603_, _03437_);
  or _72673_ (_21605_, _21604_, _21599_);
  and _72674_ (_21606_, _06211_, _05234_);
  nor _72675_ (_21607_, _21606_, _21565_);
  nand _72676_ (_21608_, _21607_, _03437_);
  and _72677_ (_21609_, _21608_, _21605_);
  nor _72678_ (_21610_, _21609_, _03636_);
  and _72679_ (_21611_, _13036_, _05234_);
  or _72680_ (_21612_, _21565_, _04499_);
  nor _72681_ (_21614_, _21612_, _21611_);
  or _72682_ (_21615_, _21614_, _03769_);
  nor _72683_ (_21616_, _21615_, _21610_);
  nor _72684_ (_21617_, _21616_, _21568_);
  nor _72685_ (_21618_, _21617_, _04504_);
  not _72686_ (_21619_, _21565_);
  and _72687_ (_21620_, _21619_, _05471_);
  or _72688_ (_21621_, _21607_, _04505_);
  nor _72689_ (_21622_, _21621_, _21620_);
  nor _72690_ (_21623_, _21622_, _21618_);
  nor _72691_ (_21625_, _21623_, _03752_);
  or _72692_ (_21626_, _21620_, _03753_);
  nor _72693_ (_21627_, _21626_, _21571_);
  or _72694_ (_21628_, _21627_, _21625_);
  and _72695_ (_21629_, _21628_, _03759_);
  nor _72696_ (_21630_, _13035_, _09299_);
  nor _72697_ (_21631_, _21630_, _21565_);
  nor _72698_ (_21632_, _21631_, _03759_);
  or _72699_ (_21633_, _21632_, _21629_);
  and _72700_ (_21634_, _21633_, _04517_);
  nor _72701_ (_21636_, _13041_, _09299_);
  nor _72702_ (_21637_, _21636_, _21565_);
  nor _72703_ (_21638_, _21637_, _04517_);
  or _72704_ (_21639_, _21638_, _03790_);
  nor _72705_ (_21640_, _21639_, _21634_);
  and _72706_ (_21641_, _21578_, _03790_);
  or _72707_ (_21642_, _21641_, _03520_);
  nor _72708_ (_21643_, _21642_, _21640_);
  and _72709_ (_21644_, _13097_, _05234_);
  nor _72710_ (_21645_, _21644_, _21565_);
  nor _72711_ (_21647_, _21645_, _03521_);
  or _72712_ (_21648_, _21647_, _21643_);
  or _72713_ (_21649_, _21648_, _42967_);
  or _72714_ (_21650_, _42963_, \oc8051_golden_model_1.TH0 [5]);
  and _72715_ (_21651_, _21650_, _41755_);
  and _72716_ (_43269_, _21651_, _21649_);
  not _72717_ (_21652_, \oc8051_golden_model_1.TH0 [6]);
  nor _72718_ (_21653_, _05234_, _21652_);
  and _72719_ (_21654_, _13259_, _05234_);
  nor _72720_ (_21655_, _21654_, _21653_);
  nor _72721_ (_21657_, _21655_, _04501_);
  and _72722_ (_21658_, _05234_, \oc8051_golden_model_1.ACC [6]);
  nor _72723_ (_21659_, _21658_, _21653_);
  nor _72724_ (_21660_, _21659_, _03583_);
  nor _72725_ (_21661_, _21659_, _04427_);
  nor _72726_ (_21662_, _04426_, _21652_);
  or _72727_ (_21663_, _21662_, _21661_);
  and _72728_ (_21664_, _21663_, _04444_);
  nor _72729_ (_21665_, _13122_, _09299_);
  nor _72730_ (_21666_, _21665_, _21653_);
  nor _72731_ (_21668_, _21666_, _04444_);
  or _72732_ (_21669_, _21668_, _21664_);
  and _72733_ (_21670_, _21669_, _03983_);
  nor _72734_ (_21671_, _05327_, _09299_);
  nor _72735_ (_21672_, _21671_, _21653_);
  nor _72736_ (_21673_, _21672_, _03983_);
  nor _72737_ (_21674_, _21673_, _21670_);
  nor _72738_ (_21675_, _21674_, _03575_);
  or _72739_ (_21676_, _21675_, _07314_);
  nor _72740_ (_21677_, _21676_, _21660_);
  and _72741_ (_21679_, _21672_, _07314_);
  nor _72742_ (_21680_, _21679_, _21677_);
  nor _72743_ (_21681_, _21680_, _03479_);
  and _72744_ (_21682_, _06713_, _05234_);
  nor _72745_ (_21683_, _21653_, _06044_);
  not _72746_ (_21684_, _21683_);
  nor _72747_ (_21685_, _21684_, _21682_);
  or _72748_ (_21686_, _21685_, _03221_);
  nor _72749_ (_21687_, _21686_, _21681_);
  nor _72750_ (_21688_, _13237_, _09299_);
  nor _72751_ (_21690_, _21688_, _21653_);
  nor _72752_ (_21691_, _21690_, _03474_);
  or _72753_ (_21692_, _21691_, _03437_);
  or _72754_ (_21693_, _21692_, _21687_);
  and _72755_ (_21694_, _13244_, _05234_);
  nor _72756_ (_21695_, _21694_, _21653_);
  nand _72757_ (_21696_, _21695_, _03437_);
  and _72758_ (_21697_, _21696_, _21693_);
  nor _72759_ (_21698_, _21697_, _03636_);
  and _72760_ (_21699_, _13253_, _05234_);
  or _72761_ (_21701_, _21653_, _04499_);
  nor _72762_ (_21702_, _21701_, _21699_);
  or _72763_ (_21703_, _21702_, _03769_);
  nor _72764_ (_21704_, _21703_, _21698_);
  nor _72765_ (_21705_, _21704_, _21657_);
  nor _72766_ (_21706_, _21705_, _04504_);
  not _72767_ (_21707_, _21653_);
  and _72768_ (_21708_, _21707_, _05376_);
  or _72769_ (_21709_, _21695_, _04505_);
  nor _72770_ (_21710_, _21709_, _21708_);
  nor _72771_ (_21712_, _21710_, _21706_);
  nor _72772_ (_21713_, _21712_, _03752_);
  or _72773_ (_21714_, _21708_, _03753_);
  or _72774_ (_21715_, _21714_, _21659_);
  and _72775_ (_21716_, _21715_, _03759_);
  not _72776_ (_21717_, _21716_);
  nor _72777_ (_21718_, _21717_, _21713_);
  nor _72778_ (_21719_, _13251_, _09299_);
  or _72779_ (_21720_, _21653_, _03759_);
  nor _72780_ (_21721_, _21720_, _21719_);
  or _72781_ (_21723_, _21721_, _03760_);
  nor _72782_ (_21724_, _21723_, _21718_);
  nor _72783_ (_21725_, _13258_, _09299_);
  nor _72784_ (_21726_, _21725_, _21653_);
  nor _72785_ (_21727_, _21726_, _04517_);
  or _72786_ (_21728_, _21727_, _03790_);
  nor _72787_ (_21729_, _21728_, _21724_);
  and _72788_ (_21730_, _21666_, _03790_);
  or _72789_ (_21731_, _21730_, _03520_);
  nor _72790_ (_21732_, _21731_, _21729_);
  and _72791_ (_21734_, _13312_, _05234_);
  nor _72792_ (_21735_, _21734_, _21653_);
  nor _72793_ (_21736_, _21735_, _03521_);
  or _72794_ (_21737_, _21736_, _21732_);
  or _72795_ (_21738_, _21737_, _42967_);
  or _72796_ (_21739_, _42963_, \oc8051_golden_model_1.TH0 [6]);
  and _72797_ (_21740_, _21739_, _41755_);
  and _72798_ (_43270_, _21740_, _21738_);
  not _72799_ (_21741_, \oc8051_golden_model_1.TH1 [0]);
  nor _72800_ (_21742_, _05251_, _21741_);
  and _72801_ (_21744_, _05941_, _05251_);
  nor _72802_ (_21745_, _21744_, _21742_);
  and _72803_ (_21746_, _21745_, _17076_);
  and _72804_ (_21747_, _05251_, \oc8051_golden_model_1.ACC [0]);
  nor _72805_ (_21748_, _21747_, _21742_);
  nor _72806_ (_21749_, _21748_, _03583_);
  nor _72807_ (_21750_, _21748_, _04427_);
  nor _72808_ (_21751_, _04426_, _21741_);
  or _72809_ (_21752_, _21751_, _21750_);
  and _72810_ (_21753_, _21752_, _04444_);
  nor _72811_ (_21755_, _21745_, _04444_);
  or _72812_ (_21756_, _21755_, _21753_);
  and _72813_ (_21757_, _21756_, _03983_);
  and _72814_ (_21758_, _05251_, _04419_);
  nor _72815_ (_21759_, _21758_, _21742_);
  nor _72816_ (_21760_, _21759_, _03983_);
  nor _72817_ (_21761_, _21760_, _21757_);
  nor _72818_ (_21762_, _21761_, _03575_);
  or _72819_ (_21763_, _21762_, _07314_);
  nor _72820_ (_21764_, _21763_, _21749_);
  and _72821_ (_21766_, _21759_, _07314_);
  nor _72822_ (_21767_, _21766_, _21764_);
  nor _72823_ (_21768_, _21767_, _03479_);
  and _72824_ (_21769_, _06715_, _05251_);
  nor _72825_ (_21770_, _21742_, _06044_);
  not _72826_ (_21771_, _21770_);
  nor _72827_ (_21772_, _21771_, _21769_);
  nor _72828_ (_21773_, _21772_, _21768_);
  nor _72829_ (_21774_, _21773_, _03221_);
  nor _72830_ (_21775_, _11975_, _09381_);
  or _72831_ (_21777_, _21742_, _03474_);
  nor _72832_ (_21778_, _21777_, _21775_);
  or _72833_ (_21779_, _21778_, _03437_);
  nor _72834_ (_21780_, _21779_, _21774_);
  and _72835_ (_21781_, _05251_, _06202_);
  nor _72836_ (_21782_, _21781_, _21742_);
  nor _72837_ (_21783_, _21782_, _03438_);
  or _72838_ (_21784_, _21783_, _21780_);
  and _72839_ (_21785_, _21784_, _04499_);
  and _72840_ (_21786_, _11990_, _05251_);
  nor _72841_ (_21788_, _21786_, _21742_);
  nor _72842_ (_21789_, _21788_, _04499_);
  or _72843_ (_21790_, _21789_, _21785_);
  nor _72844_ (_21791_, _21790_, _03769_);
  and _72845_ (_21792_, _11995_, _05251_);
  or _72846_ (_21793_, _21742_, _04501_);
  nor _72847_ (_21794_, _21793_, _21792_);
  or _72848_ (_21795_, _21794_, _04504_);
  nor _72849_ (_21796_, _21795_, _21791_);
  or _72850_ (_21797_, _21782_, _04505_);
  nor _72851_ (_21799_, _21797_, _21744_);
  nor _72852_ (_21800_, _21799_, _21796_);
  nor _72853_ (_21801_, _21800_, _03752_);
  nor _72854_ (_21802_, _21742_, _05617_);
  or _72855_ (_21803_, _21802_, _03753_);
  nor _72856_ (_21804_, _21803_, _21748_);
  or _72857_ (_21805_, _21804_, _21801_);
  and _72858_ (_21806_, _21805_, _03759_);
  nor _72859_ (_21807_, _11988_, _09381_);
  nor _72860_ (_21808_, _21807_, _21742_);
  nor _72861_ (_21810_, _21808_, _03759_);
  or _72862_ (_21811_, _21810_, _21806_);
  and _72863_ (_21812_, _21811_, _04517_);
  nor _72864_ (_21813_, _11870_, _09381_);
  nor _72865_ (_21814_, _21813_, _21742_);
  nor _72866_ (_21815_, _21814_, _04517_);
  nor _72867_ (_21816_, _21815_, _17076_);
  not _72868_ (_21817_, _21816_);
  nor _72869_ (_21818_, _21817_, _21812_);
  nor _72870_ (_21819_, _21818_, _21746_);
  or _72871_ (_21821_, _21819_, _42967_);
  or _72872_ (_21822_, _42963_, \oc8051_golden_model_1.TH1 [0]);
  and _72873_ (_21823_, _21822_, _41755_);
  and _72874_ (_43273_, _21823_, _21821_);
  and _72875_ (_21824_, _06714_, _05251_);
  not _72876_ (_21825_, \oc8051_golden_model_1.TH1 [1]);
  nor _72877_ (_21826_, _05251_, _21825_);
  nor _72878_ (_21827_, _21826_, _06044_);
  not _72879_ (_21828_, _21827_);
  nor _72880_ (_21829_, _21828_, _21824_);
  not _72881_ (_21831_, _21829_);
  nor _72882_ (_21832_, _09381_, _04603_);
  nor _72883_ (_21833_, _21832_, _21826_);
  and _72884_ (_21834_, _21833_, _07314_);
  nor _72885_ (_21835_, _05251_, \oc8051_golden_model_1.TH1 [1]);
  and _72886_ (_21836_, _05251_, _03233_);
  nor _72887_ (_21837_, _21836_, _21835_);
  and _72888_ (_21838_, _21837_, _03575_);
  nor _72889_ (_21839_, _21833_, _03983_);
  and _72890_ (_21840_, _21837_, _04426_);
  nor _72891_ (_21842_, _04426_, _21825_);
  or _72892_ (_21843_, _21842_, _21840_);
  and _72893_ (_21844_, _21843_, _04444_);
  and _72894_ (_21845_, _12252_, _05251_);
  nor _72895_ (_21846_, _21845_, _21835_);
  and _72896_ (_21847_, _21846_, _03570_);
  or _72897_ (_21848_, _21847_, _21844_);
  and _72898_ (_21849_, _21848_, _03983_);
  nor _72899_ (_21850_, _21849_, _21839_);
  nor _72900_ (_21851_, _21850_, _03575_);
  or _72901_ (_21853_, _21851_, _07314_);
  nor _72902_ (_21854_, _21853_, _21838_);
  nor _72903_ (_21855_, _21854_, _21834_);
  nor _72904_ (_21856_, _21855_, _03479_);
  nor _72905_ (_21857_, _21856_, _03221_);
  and _72906_ (_21858_, _21857_, _21831_);
  not _72907_ (_21859_, _21835_);
  and _72908_ (_21860_, _12176_, _05251_);
  nor _72909_ (_21861_, _21860_, _03474_);
  and _72910_ (_21862_, _21861_, _21859_);
  nor _72911_ (_21864_, _21862_, _21858_);
  nor _72912_ (_21865_, _21864_, _03437_);
  and _72913_ (_21866_, _05251_, _04317_);
  not _72914_ (_21867_, _21866_);
  nor _72915_ (_21868_, _21835_, _03438_);
  and _72916_ (_21869_, _21868_, _21867_);
  nor _72917_ (_21870_, _21869_, _21865_);
  nor _72918_ (_21871_, _21870_, _03636_);
  nor _72919_ (_21872_, _12191_, _09381_);
  nor _72920_ (_21873_, _21872_, _04499_);
  and _72921_ (_21875_, _21873_, _21859_);
  nor _72922_ (_21876_, _21875_, _21871_);
  nor _72923_ (_21877_, _21876_, _03769_);
  nor _72924_ (_21878_, _12197_, _09381_);
  nor _72925_ (_21879_, _21878_, _04501_);
  and _72926_ (_21880_, _21879_, _21859_);
  nor _72927_ (_21881_, _21880_, _21877_);
  nor _72928_ (_21882_, _21881_, _04504_);
  nor _72929_ (_21883_, _12190_, _09381_);
  nor _72930_ (_21884_, _21883_, _05769_);
  and _72931_ (_21886_, _21884_, _21859_);
  nor _72932_ (_21887_, _21886_, _21882_);
  nor _72933_ (_21888_, _21887_, _03752_);
  nor _72934_ (_21889_, _21826_, _05569_);
  nor _72935_ (_21890_, _21889_, _03753_);
  and _72936_ (_21891_, _21890_, _21837_);
  nor _72937_ (_21892_, _21891_, _21888_);
  nor _72938_ (_21893_, _21892_, _03758_);
  and _72939_ (_21894_, _21866_, _05940_);
  nor _72940_ (_21895_, _21894_, _03759_);
  and _72941_ (_21897_, _21895_, _21859_);
  nor _72942_ (_21898_, _21897_, _21893_);
  nor _72943_ (_21899_, _21898_, _03760_);
  nand _72944_ (_21900_, _21836_, _05940_);
  nor _72945_ (_21901_, _21835_, _04517_);
  and _72946_ (_21902_, _21901_, _21900_);
  or _72947_ (_21903_, _21902_, _21899_);
  and _72948_ (_21904_, _21903_, _04192_);
  and _72949_ (_21905_, _21846_, _03790_);
  or _72950_ (_21906_, _21905_, _21904_);
  and _72951_ (_21908_, _21906_, _03521_);
  nor _72952_ (_21909_, _21826_, _21845_);
  nor _72953_ (_21910_, _21909_, _03521_);
  or _72954_ (_21911_, _21910_, _21908_);
  or _72955_ (_21912_, _21911_, _42967_);
  or _72956_ (_21913_, _42963_, \oc8051_golden_model_1.TH1 [1]);
  and _72957_ (_21914_, _21913_, _41755_);
  and _72958_ (_43274_, _21914_, _21912_);
  not _72959_ (_21915_, \oc8051_golden_model_1.TH1 [2]);
  nor _72960_ (_21916_, _05251_, _21915_);
  nor _72961_ (_21918_, _12400_, _09381_);
  nor _72962_ (_21919_, _21918_, _21916_);
  nor _72963_ (_21920_, _21919_, _04517_);
  and _72964_ (_21921_, _05251_, \oc8051_golden_model_1.ACC [2]);
  nor _72965_ (_21922_, _21921_, _21916_);
  nor _72966_ (_21923_, _21922_, _03583_);
  nor _72967_ (_21924_, _21922_, _04427_);
  nor _72968_ (_21925_, _04426_, _21915_);
  or _72969_ (_21926_, _21925_, _21924_);
  and _72970_ (_21927_, _21926_, _04444_);
  nor _72971_ (_21929_, _12282_, _09381_);
  nor _72972_ (_21930_, _21929_, _21916_);
  nor _72973_ (_21931_, _21930_, _04444_);
  or _72974_ (_21932_, _21931_, _21927_);
  and _72975_ (_21933_, _21932_, _03983_);
  nor _72976_ (_21934_, _09381_, _05026_);
  nor _72977_ (_21935_, _21934_, _21916_);
  nor _72978_ (_21936_, _21935_, _03983_);
  nor _72979_ (_21937_, _21936_, _21933_);
  nor _72980_ (_21938_, _21937_, _03575_);
  or _72981_ (_21940_, _21938_, _07314_);
  nor _72982_ (_21941_, _21940_, _21923_);
  and _72983_ (_21942_, _21935_, _07314_);
  nor _72984_ (_21943_, _21942_, _21941_);
  nor _72985_ (_21944_, _21943_, _03479_);
  and _72986_ (_21945_, _06718_, _05251_);
  nor _72987_ (_21946_, _21916_, _06044_);
  not _72988_ (_21947_, _21946_);
  nor _72989_ (_21948_, _21947_, _21945_);
  nor _72990_ (_21949_, _21948_, _21944_);
  nor _72991_ (_21951_, _21949_, _03221_);
  nor _72992_ (_21952_, _12384_, _09381_);
  or _72993_ (_21953_, _21916_, _03474_);
  nor _72994_ (_21954_, _21953_, _21952_);
  or _72995_ (_21955_, _21954_, _03437_);
  nor _72996_ (_21956_, _21955_, _21951_);
  and _72997_ (_21957_, _05251_, _06261_);
  nor _72998_ (_21958_, _21957_, _21916_);
  nor _72999_ (_21959_, _21958_, _03438_);
  or _73000_ (_21960_, _21959_, _21956_);
  and _73001_ (_21962_, _21960_, _04499_);
  and _73002_ (_21963_, _12273_, _05251_);
  nor _73003_ (_21964_, _21963_, _21916_);
  nor _73004_ (_21965_, _21964_, _04499_);
  or _73005_ (_21966_, _21965_, _21962_);
  nor _73006_ (_21967_, _21966_, _03769_);
  and _73007_ (_21968_, _12401_, _05251_);
  or _73008_ (_21969_, _21916_, _04501_);
  nor _73009_ (_21970_, _21969_, _21968_);
  or _73010_ (_21971_, _21970_, _04504_);
  nor _73011_ (_21973_, _21971_, _21967_);
  nor _73012_ (_21974_, _21916_, _05665_);
  or _73013_ (_21975_, _21958_, _04505_);
  nor _73014_ (_21976_, _21975_, _21974_);
  nor _73015_ (_21977_, _21976_, _21973_);
  nor _73016_ (_21978_, _21977_, _03752_);
  or _73017_ (_21979_, _21974_, _03753_);
  nor _73018_ (_21980_, _21979_, _21922_);
  or _73019_ (_21981_, _21980_, _21978_);
  and _73020_ (_21982_, _21981_, _03759_);
  nor _73021_ (_21984_, _12272_, _09381_);
  nor _73022_ (_21985_, _21984_, _21916_);
  nor _73023_ (_21986_, _21985_, _03759_);
  or _73024_ (_21987_, _21986_, _21982_);
  and _73025_ (_21988_, _21987_, _04517_);
  nor _73026_ (_21989_, _21988_, _21920_);
  nor _73027_ (_21990_, _21989_, _03790_);
  nor _73028_ (_21991_, _21930_, _04192_);
  or _73029_ (_21992_, _21991_, _03520_);
  nor _73030_ (_21993_, _21992_, _21990_);
  and _73031_ (_21995_, _12456_, _05251_);
  or _73032_ (_21996_, _21916_, _03521_);
  nor _73033_ (_21997_, _21996_, _21995_);
  nor _73034_ (_21998_, _21997_, _21993_);
  or _73035_ (_21999_, _21998_, _42967_);
  or _73036_ (_22000_, _42963_, \oc8051_golden_model_1.TH1 [2]);
  and _73037_ (_22001_, _22000_, _41755_);
  and _73038_ (_43275_, _22001_, _21999_);
  not _73039_ (_22002_, \oc8051_golden_model_1.TH1 [3]);
  nor _73040_ (_22003_, _05251_, _22002_);
  and _73041_ (_22005_, _12604_, _05251_);
  nor _73042_ (_22006_, _22005_, _22003_);
  nor _73043_ (_22007_, _22006_, _04501_);
  nor _73044_ (_22008_, _09381_, _04843_);
  nor _73045_ (_22009_, _22008_, _22003_);
  and _73046_ (_22010_, _22009_, _07314_);
  and _73047_ (_22011_, _05251_, \oc8051_golden_model_1.ACC [3]);
  nor _73048_ (_22012_, _22011_, _22003_);
  nor _73049_ (_22013_, _22012_, _03583_);
  nor _73050_ (_22014_, _22012_, _04427_);
  nor _73051_ (_22016_, _04426_, _22002_);
  or _73052_ (_22017_, _22016_, _22014_);
  and _73053_ (_22018_, _22017_, _04444_);
  nor _73054_ (_22019_, _12486_, _09381_);
  nor _73055_ (_22020_, _22019_, _22003_);
  nor _73056_ (_22021_, _22020_, _04444_);
  or _73057_ (_22022_, _22021_, _22018_);
  and _73058_ (_22023_, _22022_, _03983_);
  nor _73059_ (_22024_, _22009_, _03983_);
  nor _73060_ (_22025_, _22024_, _22023_);
  nor _73061_ (_22027_, _22025_, _03575_);
  or _73062_ (_22028_, _22027_, _07314_);
  nor _73063_ (_22029_, _22028_, _22013_);
  nor _73064_ (_22030_, _22029_, _22010_);
  nor _73065_ (_22031_, _22030_, _03479_);
  and _73066_ (_22032_, _06717_, _05251_);
  nor _73067_ (_22033_, _22003_, _06044_);
  not _73068_ (_22034_, _22033_);
  nor _73069_ (_22035_, _22034_, _22032_);
  or _73070_ (_22036_, _22035_, _03221_);
  nor _73071_ (_22038_, _22036_, _22031_);
  nor _73072_ (_22039_, _12583_, _09381_);
  nor _73073_ (_22040_, _22039_, _22003_);
  nor _73074_ (_22041_, _22040_, _03474_);
  or _73075_ (_22042_, _22041_, _03437_);
  or _73076_ (_22043_, _22042_, _22038_);
  and _73077_ (_22044_, _05251_, _06217_);
  nor _73078_ (_22045_, _22044_, _22003_);
  nand _73079_ (_22046_, _22045_, _03437_);
  and _73080_ (_22047_, _22046_, _22043_);
  nor _73081_ (_22049_, _22047_, _03636_);
  and _73082_ (_22050_, _12598_, _05251_);
  or _73083_ (_22051_, _22003_, _04499_);
  nor _73084_ (_22052_, _22051_, _22050_);
  or _73085_ (_22053_, _22052_, _03769_);
  nor _73086_ (_22054_, _22053_, _22049_);
  nor _73087_ (_22055_, _22054_, _22007_);
  nor _73088_ (_22056_, _22055_, _04504_);
  not _73089_ (_22057_, _22003_);
  and _73090_ (_22058_, _22057_, _05520_);
  or _73091_ (_22059_, _22045_, _04505_);
  nor _73092_ (_22060_, _22059_, _22058_);
  nor _73093_ (_22061_, _22060_, _22056_);
  nor _73094_ (_22062_, _22061_, _03752_);
  or _73095_ (_22063_, _22058_, _03753_);
  nor _73096_ (_22064_, _22063_, _22012_);
  or _73097_ (_22065_, _22064_, _22062_);
  and _73098_ (_22066_, _22065_, _03759_);
  nor _73099_ (_22067_, _12597_, _09381_);
  nor _73100_ (_22068_, _22067_, _22003_);
  nor _73101_ (_22071_, _22068_, _03759_);
  or _73102_ (_22072_, _22071_, _22066_);
  and _73103_ (_22073_, _22072_, _04517_);
  nor _73104_ (_22074_, _12603_, _09381_);
  nor _73105_ (_22075_, _22074_, _22003_);
  nor _73106_ (_22076_, _22075_, _04517_);
  or _73107_ (_22077_, _22076_, _03790_);
  nor _73108_ (_22078_, _22077_, _22073_);
  and _73109_ (_22079_, _22020_, _03790_);
  or _73110_ (_22080_, _22079_, _03520_);
  nor _73111_ (_22082_, _22080_, _22078_);
  and _73112_ (_22083_, _12658_, _05251_);
  nor _73113_ (_22084_, _22083_, _22003_);
  nor _73114_ (_22085_, _22084_, _03521_);
  or _73115_ (_22086_, _22085_, _22082_);
  or _73116_ (_22087_, _22086_, _42967_);
  or _73117_ (_22088_, _42963_, \oc8051_golden_model_1.TH1 [3]);
  and _73118_ (_22089_, _22088_, _41755_);
  and _73119_ (_43276_, _22089_, _22087_);
  not _73120_ (_22090_, \oc8051_golden_model_1.TH1 [4]);
  nor _73121_ (_22092_, _05251_, _22090_);
  and _73122_ (_22093_, _12844_, _05251_);
  nor _73123_ (_22094_, _22093_, _22092_);
  nor _73124_ (_22095_, _22094_, _04501_);
  and _73125_ (_22096_, _05251_, \oc8051_golden_model_1.ACC [4]);
  nor _73126_ (_22097_, _22096_, _22092_);
  nor _73127_ (_22098_, _22097_, _03583_);
  nor _73128_ (_22099_, _22097_, _04427_);
  nor _73129_ (_22100_, _04426_, _22090_);
  or _73130_ (_22101_, _22100_, _22099_);
  and _73131_ (_22103_, _22101_, _04444_);
  nor _73132_ (_22104_, _12733_, _09381_);
  nor _73133_ (_22105_, _22104_, _22092_);
  nor _73134_ (_22106_, _22105_, _04444_);
  or _73135_ (_22107_, _22106_, _22103_);
  and _73136_ (_22108_, _22107_, _03983_);
  nor _73137_ (_22109_, _05712_, _09381_);
  nor _73138_ (_22110_, _22109_, _22092_);
  nor _73139_ (_22111_, _22110_, _03983_);
  nor _73140_ (_22112_, _22111_, _22108_);
  nor _73141_ (_22114_, _22112_, _03575_);
  or _73142_ (_22115_, _22114_, _07314_);
  nor _73143_ (_22116_, _22115_, _22098_);
  and _73144_ (_22117_, _22110_, _07314_);
  or _73145_ (_22118_, _22117_, _03479_);
  nor _73146_ (_22119_, _22118_, _22116_);
  and _73147_ (_22120_, _06722_, _05251_);
  or _73148_ (_22121_, _22120_, _22092_);
  and _73149_ (_22122_, _22121_, _03479_);
  or _73150_ (_22123_, _22122_, _03221_);
  or _73151_ (_22125_, _22123_, _22119_);
  nor _73152_ (_22126_, _12827_, _09381_);
  or _73153_ (_22127_, _22092_, _03474_);
  or _73154_ (_22128_, _22127_, _22126_);
  and _73155_ (_22129_, _22128_, _03438_);
  and _73156_ (_22130_, _22129_, _22125_);
  and _73157_ (_22131_, _06233_, _05251_);
  nor _73158_ (_22132_, _22131_, _22092_);
  nor _73159_ (_22133_, _22132_, _03438_);
  or _73160_ (_22134_, _22133_, _03636_);
  nor _73161_ (_22136_, _22134_, _22130_);
  and _73162_ (_22137_, _12711_, _05251_);
  or _73163_ (_22138_, _22092_, _04499_);
  nor _73164_ (_22139_, _22138_, _22137_);
  or _73165_ (_22140_, _22139_, _03769_);
  nor _73166_ (_22141_, _22140_, _22136_);
  nor _73167_ (_22142_, _22141_, _22095_);
  nor _73168_ (_22143_, _22142_, _04504_);
  not _73169_ (_22144_, _22092_);
  and _73170_ (_22145_, _22144_, _05760_);
  or _73171_ (_22147_, _22132_, _04505_);
  nor _73172_ (_22148_, _22147_, _22145_);
  nor _73173_ (_22149_, _22148_, _22143_);
  nor _73174_ (_22150_, _22149_, _03752_);
  or _73175_ (_22151_, _22145_, _03753_);
  or _73176_ (_22152_, _22151_, _22097_);
  and _73177_ (_22153_, _22152_, _03759_);
  not _73178_ (_22154_, _22153_);
  nor _73179_ (_22155_, _22154_, _22150_);
  nor _73180_ (_22156_, _12710_, _09381_);
  or _73181_ (_22158_, _22092_, _03759_);
  nor _73182_ (_22159_, _22158_, _22156_);
  or _73183_ (_22160_, _22159_, _03760_);
  nor _73184_ (_22161_, _22160_, _22155_);
  nor _73185_ (_22162_, _12843_, _09381_);
  nor _73186_ (_22163_, _22162_, _22092_);
  nor _73187_ (_22164_, _22163_, _04517_);
  or _73188_ (_22165_, _22164_, _03790_);
  nor _73189_ (_22166_, _22165_, _22161_);
  and _73190_ (_22167_, _22105_, _03790_);
  or _73191_ (_22169_, _22167_, _03520_);
  nor _73192_ (_22170_, _22169_, _22166_);
  and _73193_ (_22171_, _12893_, _05251_);
  nor _73194_ (_22172_, _22171_, _22092_);
  nor _73195_ (_22173_, _22172_, _03521_);
  or _73196_ (_22174_, _22173_, _22170_);
  or _73197_ (_22175_, _22174_, _42967_);
  or _73198_ (_22176_, _42963_, \oc8051_golden_model_1.TH1 [4]);
  and _73199_ (_22177_, _22176_, _41755_);
  and _73200_ (_43277_, _22177_, _22175_);
  not _73201_ (_22179_, \oc8051_golden_model_1.TH1 [5]);
  nor _73202_ (_22180_, _05251_, _22179_);
  and _73203_ (_22181_, _13042_, _05251_);
  nor _73204_ (_22182_, _22181_, _22180_);
  nor _73205_ (_22183_, _22182_, _04501_);
  and _73206_ (_22184_, _05251_, \oc8051_golden_model_1.ACC [5]);
  nor _73207_ (_22185_, _22184_, _22180_);
  nor _73208_ (_22186_, _22185_, _03583_);
  nor _73209_ (_22187_, _22185_, _04427_);
  nor _73210_ (_22188_, _04426_, _22179_);
  or _73211_ (_22190_, _22188_, _22187_);
  and _73212_ (_22191_, _22190_, _04444_);
  nor _73213_ (_22192_, _12930_, _09381_);
  nor _73214_ (_22193_, _22192_, _22180_);
  nor _73215_ (_22194_, _22193_, _04444_);
  or _73216_ (_22195_, _22194_, _22191_);
  and _73217_ (_22196_, _22195_, _03983_);
  nor _73218_ (_22197_, _05422_, _09381_);
  nor _73219_ (_22198_, _22197_, _22180_);
  nor _73220_ (_22199_, _22198_, _03983_);
  nor _73221_ (_22201_, _22199_, _22196_);
  nor _73222_ (_22202_, _22201_, _03575_);
  or _73223_ (_22203_, _22202_, _07314_);
  nor _73224_ (_22204_, _22203_, _22186_);
  and _73225_ (_22205_, _22198_, _07314_);
  nor _73226_ (_22206_, _22205_, _22204_);
  nor _73227_ (_22207_, _22206_, _03479_);
  and _73228_ (_22208_, _06721_, _05251_);
  nor _73229_ (_22209_, _22180_, _06044_);
  not _73230_ (_22210_, _22209_);
  nor _73231_ (_22212_, _22210_, _22208_);
  or _73232_ (_22213_, _22212_, _03221_);
  nor _73233_ (_22214_, _22213_, _22207_);
  nor _73234_ (_22215_, _13021_, _09381_);
  nor _73235_ (_22216_, _22215_, _22180_);
  nor _73236_ (_22217_, _22216_, _03474_);
  or _73237_ (_22218_, _22217_, _03437_);
  or _73238_ (_22219_, _22218_, _22214_);
  and _73239_ (_22220_, _06211_, _05251_);
  nor _73240_ (_22221_, _22220_, _22180_);
  nand _73241_ (_22223_, _22221_, _03437_);
  and _73242_ (_22224_, _22223_, _22219_);
  nor _73243_ (_22225_, _22224_, _03636_);
  and _73244_ (_22226_, _13036_, _05251_);
  or _73245_ (_22227_, _22180_, _04499_);
  nor _73246_ (_22228_, _22227_, _22226_);
  or _73247_ (_22229_, _22228_, _03769_);
  nor _73248_ (_22230_, _22229_, _22225_);
  nor _73249_ (_22231_, _22230_, _22183_);
  nor _73250_ (_22232_, _22231_, _04504_);
  not _73251_ (_22234_, _22180_);
  and _73252_ (_22235_, _22234_, _05471_);
  or _73253_ (_22236_, _22221_, _04505_);
  nor _73254_ (_22237_, _22236_, _22235_);
  nor _73255_ (_22238_, _22237_, _22232_);
  nor _73256_ (_22239_, _22238_, _03752_);
  or _73257_ (_22240_, _22235_, _03753_);
  or _73258_ (_22241_, _22240_, _22185_);
  and _73259_ (_22242_, _22241_, _03759_);
  not _73260_ (_22243_, _22242_);
  nor _73261_ (_22245_, _22243_, _22239_);
  nor _73262_ (_22246_, _13035_, _09381_);
  or _73263_ (_22247_, _22180_, _03759_);
  nor _73264_ (_22248_, _22247_, _22246_);
  or _73265_ (_22249_, _22248_, _03760_);
  nor _73266_ (_22250_, _22249_, _22245_);
  nor _73267_ (_22251_, _13041_, _09381_);
  nor _73268_ (_22252_, _22251_, _22180_);
  nor _73269_ (_22253_, _22252_, _04517_);
  or _73270_ (_22254_, _22253_, _03790_);
  nor _73271_ (_22256_, _22254_, _22250_);
  and _73272_ (_22257_, _22193_, _03790_);
  or _73273_ (_22258_, _22257_, _03520_);
  nor _73274_ (_22259_, _22258_, _22256_);
  and _73275_ (_22260_, _13097_, _05251_);
  nor _73276_ (_22261_, _22260_, _22180_);
  nor _73277_ (_22262_, _22261_, _03521_);
  or _73278_ (_22263_, _22262_, _22259_);
  or _73279_ (_22264_, _22263_, _42967_);
  or _73280_ (_22265_, _42963_, \oc8051_golden_model_1.TH1 [5]);
  and _73281_ (_22267_, _22265_, _41755_);
  and _73282_ (_43278_, _22267_, _22264_);
  not _73283_ (_22268_, \oc8051_golden_model_1.TH1 [6]);
  nor _73284_ (_22269_, _05251_, _22268_);
  and _73285_ (_22270_, _13259_, _05251_);
  nor _73286_ (_22271_, _22270_, _22269_);
  nor _73287_ (_22272_, _22271_, _04501_);
  and _73288_ (_22273_, _05251_, \oc8051_golden_model_1.ACC [6]);
  nor _73289_ (_22274_, _22273_, _22269_);
  nor _73290_ (_22275_, _22274_, _03583_);
  nor _73291_ (_22277_, _22274_, _04427_);
  nor _73292_ (_22278_, _04426_, _22268_);
  or _73293_ (_22279_, _22278_, _22277_);
  and _73294_ (_22280_, _22279_, _04444_);
  nor _73295_ (_22281_, _13122_, _09381_);
  nor _73296_ (_22282_, _22281_, _22269_);
  nor _73297_ (_22283_, _22282_, _04444_);
  or _73298_ (_22284_, _22283_, _22280_);
  and _73299_ (_22285_, _22284_, _03983_);
  nor _73300_ (_22286_, _05327_, _09381_);
  nor _73301_ (_22288_, _22286_, _22269_);
  nor _73302_ (_22289_, _22288_, _03983_);
  nor _73303_ (_22290_, _22289_, _22285_);
  nor _73304_ (_22291_, _22290_, _03575_);
  or _73305_ (_22292_, _22291_, _07314_);
  nor _73306_ (_22293_, _22292_, _22275_);
  and _73307_ (_22294_, _22288_, _07314_);
  nor _73308_ (_22295_, _22294_, _22293_);
  nor _73309_ (_22296_, _22295_, _03479_);
  and _73310_ (_22297_, _06713_, _05251_);
  nor _73311_ (_22299_, _22269_, _06044_);
  not _73312_ (_22300_, _22299_);
  nor _73313_ (_22301_, _22300_, _22297_);
  or _73314_ (_22302_, _22301_, _03221_);
  nor _73315_ (_22303_, _22302_, _22296_);
  nor _73316_ (_22304_, _13237_, _09381_);
  nor _73317_ (_22305_, _22304_, _22269_);
  nor _73318_ (_22306_, _22305_, _03474_);
  or _73319_ (_22307_, _22306_, _03437_);
  or _73320_ (_22308_, _22307_, _22303_);
  and _73321_ (_22310_, _13244_, _05251_);
  nor _73322_ (_22311_, _22310_, _22269_);
  nand _73323_ (_22312_, _22311_, _03437_);
  and _73324_ (_22313_, _22312_, _22308_);
  nor _73325_ (_22314_, _22313_, _03636_);
  and _73326_ (_22315_, _13253_, _05251_);
  or _73327_ (_22316_, _22269_, _04499_);
  nor _73328_ (_22317_, _22316_, _22315_);
  or _73329_ (_22318_, _22317_, _03769_);
  nor _73330_ (_22319_, _22318_, _22314_);
  nor _73331_ (_22321_, _22319_, _22272_);
  nor _73332_ (_22322_, _22321_, _04504_);
  not _73333_ (_22323_, _22269_);
  and _73334_ (_22324_, _22323_, _05376_);
  or _73335_ (_22325_, _22311_, _04505_);
  nor _73336_ (_22326_, _22325_, _22324_);
  nor _73337_ (_22327_, _22326_, _22322_);
  nor _73338_ (_22328_, _22327_, _03752_);
  or _73339_ (_22329_, _22324_, _03753_);
  nor _73340_ (_22330_, _22329_, _22274_);
  or _73341_ (_22333_, _22330_, _22328_);
  and _73342_ (_22334_, _22333_, _03759_);
  nor _73343_ (_22335_, _13251_, _09381_);
  nor _73344_ (_22336_, _22335_, _22269_);
  nor _73345_ (_22337_, _22336_, _03759_);
  or _73346_ (_22338_, _22337_, _22334_);
  and _73347_ (_22339_, _22338_, _04517_);
  nor _73348_ (_22340_, _13258_, _09381_);
  nor _73349_ (_22341_, _22340_, _22269_);
  nor _73350_ (_22342_, _22341_, _04517_);
  or _73351_ (_22344_, _22342_, _03790_);
  nor _73352_ (_22345_, _22344_, _22339_);
  and _73353_ (_22346_, _22282_, _03790_);
  or _73354_ (_22347_, _22346_, _03520_);
  nor _73355_ (_22348_, _22347_, _22345_);
  and _73356_ (_22349_, _13312_, _05251_);
  nor _73357_ (_22350_, _22349_, _22269_);
  nor _73358_ (_22351_, _22350_, _03521_);
  or _73359_ (_22352_, _22351_, _22348_);
  or _73360_ (_22353_, _22352_, _42967_);
  or _73361_ (_22355_, _42963_, \oc8051_golden_model_1.TH1 [6]);
  and _73362_ (_22356_, _22355_, _41755_);
  and _73363_ (_43279_, _22356_, _22353_);
  not _73364_ (_22357_, \oc8051_golden_model_1.TMOD [0]);
  nor _73365_ (_22358_, _05254_, _22357_);
  and _73366_ (_22359_, _05941_, _05254_);
  nor _73367_ (_22360_, _22359_, _22358_);
  and _73368_ (_22361_, _22360_, _17076_);
  and _73369_ (_22362_, _05254_, \oc8051_golden_model_1.ACC [0]);
  nor _73370_ (_22363_, _22362_, _22358_);
  nor _73371_ (_22365_, _22363_, _03583_);
  nor _73372_ (_22366_, _22363_, _04427_);
  nor _73373_ (_22367_, _04426_, _22357_);
  or _73374_ (_22368_, _22367_, _22366_);
  and _73375_ (_22369_, _22368_, _04444_);
  nor _73376_ (_22370_, _22360_, _04444_);
  or _73377_ (_22371_, _22370_, _22369_);
  and _73378_ (_22372_, _22371_, _03983_);
  and _73379_ (_22373_, _05254_, _04419_);
  nor _73380_ (_22374_, _22373_, _22358_);
  nor _73381_ (_22376_, _22374_, _03983_);
  nor _73382_ (_22377_, _22376_, _22372_);
  nor _73383_ (_22378_, _22377_, _03575_);
  or _73384_ (_22379_, _22378_, _07314_);
  nor _73385_ (_22380_, _22379_, _22365_);
  and _73386_ (_22381_, _22374_, _07314_);
  nor _73387_ (_22382_, _22381_, _22380_);
  nor _73388_ (_22383_, _22382_, _03479_);
  and _73389_ (_22384_, _06715_, _05254_);
  nor _73390_ (_22385_, _22358_, _06044_);
  not _73391_ (_22387_, _22385_);
  nor _73392_ (_22388_, _22387_, _22384_);
  nor _73393_ (_22389_, _22388_, _22383_);
  nor _73394_ (_22390_, _22389_, _03221_);
  nor _73395_ (_22391_, _11975_, _09462_);
  or _73396_ (_22392_, _22358_, _03474_);
  nor _73397_ (_22393_, _22392_, _22391_);
  or _73398_ (_22394_, _22393_, _03437_);
  nor _73399_ (_22395_, _22394_, _22390_);
  and _73400_ (_22396_, _05254_, _06202_);
  nor _73401_ (_22398_, _22396_, _22358_);
  nor _73402_ (_22399_, _22398_, _03438_);
  or _73403_ (_22400_, _22399_, _22395_);
  and _73404_ (_22401_, _22400_, _04499_);
  and _73405_ (_22402_, _11990_, _05254_);
  nor _73406_ (_22403_, _22402_, _22358_);
  nor _73407_ (_22404_, _22403_, _04499_);
  or _73408_ (_22405_, _22404_, _22401_);
  nor _73409_ (_22406_, _22405_, _03769_);
  and _73410_ (_22407_, _11995_, _05254_);
  or _73411_ (_22409_, _22358_, _04501_);
  nor _73412_ (_22410_, _22409_, _22407_);
  or _73413_ (_22411_, _22410_, _04504_);
  nor _73414_ (_22412_, _22411_, _22406_);
  or _73415_ (_22413_, _22398_, _04505_);
  nor _73416_ (_22414_, _22413_, _22359_);
  nor _73417_ (_22415_, _22414_, _22412_);
  nor _73418_ (_22416_, _22415_, _03752_);
  and _73419_ (_22417_, _11994_, _05254_);
  or _73420_ (_22418_, _22417_, _22358_);
  and _73421_ (_22420_, _22418_, _03752_);
  or _73422_ (_22421_, _22420_, _22416_);
  and _73423_ (_22422_, _22421_, _03759_);
  nor _73424_ (_22423_, _11988_, _09462_);
  nor _73425_ (_22424_, _22423_, _22358_);
  nor _73426_ (_22425_, _22424_, _03759_);
  or _73427_ (_22426_, _22425_, _22422_);
  and _73428_ (_22427_, _22426_, _04517_);
  nor _73429_ (_22428_, _11870_, _09462_);
  nor _73430_ (_22429_, _22428_, _22358_);
  nor _73431_ (_22431_, _22429_, _04517_);
  nor _73432_ (_22432_, _22431_, _17076_);
  not _73433_ (_22433_, _22432_);
  nor _73434_ (_22434_, _22433_, _22427_);
  nor _73435_ (_22435_, _22434_, _22361_);
  or _73436_ (_22436_, _22435_, _42967_);
  or _73437_ (_22437_, _42963_, \oc8051_golden_model_1.TMOD [0]);
  and _73438_ (_22438_, _22437_, _41755_);
  and _73439_ (_43282_, _22438_, _22436_);
  nor _73440_ (_22439_, _05254_, \oc8051_golden_model_1.TMOD [1]);
  and _73441_ (_22442_, _12252_, _05254_);
  nor _73442_ (_22443_, _22442_, _22439_);
  nor _73443_ (_22444_, _22443_, _04192_);
  and _73444_ (_22445_, _06714_, _05254_);
  not _73445_ (_22446_, \oc8051_golden_model_1.TMOD [1]);
  nor _73446_ (_22447_, _05254_, _22446_);
  nor _73447_ (_22448_, _22447_, _06044_);
  not _73448_ (_22449_, _22448_);
  nor _73449_ (_22450_, _22449_, _22445_);
  not _73450_ (_22451_, _22450_);
  nor _73451_ (_22453_, _09462_, _04603_);
  nor _73452_ (_22454_, _22453_, _22447_);
  and _73453_ (_22455_, _22454_, _07314_);
  nor _73454_ (_22456_, _22454_, _03983_);
  and _73455_ (_22457_, _05254_, _03233_);
  nor _73456_ (_22458_, _22457_, _22439_);
  and _73457_ (_22459_, _22458_, _04426_);
  nor _73458_ (_22460_, _04426_, _22446_);
  or _73459_ (_22461_, _22460_, _22459_);
  and _73460_ (_22462_, _22461_, _04444_);
  and _73461_ (_22464_, _22443_, _03570_);
  or _73462_ (_22465_, _22464_, _22462_);
  and _73463_ (_22466_, _22465_, _03983_);
  nor _73464_ (_22467_, _22466_, _22456_);
  nor _73465_ (_22468_, _22467_, _03575_);
  and _73466_ (_22469_, _22458_, _03575_);
  nor _73467_ (_22470_, _22469_, _07314_);
  not _73468_ (_22471_, _22470_);
  nor _73469_ (_22472_, _22471_, _22468_);
  nor _73470_ (_22473_, _22472_, _22455_);
  nor _73471_ (_22475_, _22473_, _03479_);
  nor _73472_ (_22476_, _22475_, _03221_);
  and _73473_ (_22477_, _22476_, _22451_);
  not _73474_ (_22478_, _22439_);
  and _73475_ (_22479_, _12176_, _05254_);
  nor _73476_ (_22480_, _22479_, _03474_);
  and _73477_ (_22481_, _22480_, _22478_);
  nor _73478_ (_22482_, _22481_, _22477_);
  nor _73479_ (_22483_, _22482_, _03437_);
  and _73480_ (_22484_, _05254_, _04317_);
  not _73481_ (_22486_, _22484_);
  nor _73482_ (_22487_, _22439_, _03438_);
  and _73483_ (_22488_, _22487_, _22486_);
  nor _73484_ (_22489_, _22488_, _22483_);
  nor _73485_ (_22490_, _22489_, _03636_);
  nor _73486_ (_22491_, _12191_, _09462_);
  nor _73487_ (_22492_, _22491_, _04499_);
  and _73488_ (_22493_, _22492_, _22478_);
  nor _73489_ (_22494_, _22493_, _22490_);
  nor _73490_ (_22495_, _22494_, _03769_);
  nor _73491_ (_22497_, _12197_, _09462_);
  nor _73492_ (_22498_, _22497_, _04501_);
  and _73493_ (_22499_, _22498_, _22478_);
  nor _73494_ (_22500_, _22499_, _22495_);
  nor _73495_ (_22501_, _22500_, _04504_);
  nor _73496_ (_22502_, _12190_, _09462_);
  nor _73497_ (_22503_, _22502_, _05769_);
  and _73498_ (_22504_, _22503_, _22478_);
  nor _73499_ (_22505_, _22504_, _22501_);
  nor _73500_ (_22506_, _22505_, _03752_);
  nor _73501_ (_22508_, _22447_, _05569_);
  nor _73502_ (_22509_, _22508_, _03753_);
  and _73503_ (_22510_, _22509_, _22458_);
  nor _73504_ (_22511_, _22510_, _22506_);
  nor _73505_ (_22512_, _22511_, _03758_);
  and _73506_ (_22513_, _22484_, _05940_);
  nor _73507_ (_22514_, _22513_, _03759_);
  and _73508_ (_22515_, _22514_, _22478_);
  nor _73509_ (_22516_, _22515_, _22512_);
  nor _73510_ (_22517_, _22516_, _03760_);
  nand _73511_ (_22519_, _22457_, _05940_);
  nor _73512_ (_22520_, _22439_, _04517_);
  and _73513_ (_22521_, _22520_, _22519_);
  or _73514_ (_22522_, _22521_, _03790_);
  nor _73515_ (_22523_, _22522_, _22517_);
  nor _73516_ (_22524_, _22523_, _22444_);
  and _73517_ (_22525_, _22524_, _03521_);
  nor _73518_ (_22526_, _22447_, _22442_);
  nor _73519_ (_22527_, _22526_, _03521_);
  or _73520_ (_22528_, _22527_, _22525_);
  or _73521_ (_22530_, _22528_, _42967_);
  or _73522_ (_22531_, _42963_, \oc8051_golden_model_1.TMOD [1]);
  and _73523_ (_22532_, _22531_, _41755_);
  and _73524_ (_43283_, _22532_, _22530_);
  not _73525_ (_22533_, \oc8051_golden_model_1.TMOD [2]);
  nor _73526_ (_22534_, _05254_, _22533_);
  nor _73527_ (_22535_, _12400_, _09462_);
  nor _73528_ (_22536_, _22535_, _22534_);
  nor _73529_ (_22537_, _22536_, _04517_);
  and _73530_ (_22538_, _05254_, \oc8051_golden_model_1.ACC [2]);
  nor _73531_ (_22540_, _22538_, _22534_);
  nor _73532_ (_22541_, _22540_, _03583_);
  nor _73533_ (_22542_, _22540_, _04427_);
  nor _73534_ (_22543_, _04426_, _22533_);
  or _73535_ (_22544_, _22543_, _22542_);
  and _73536_ (_22545_, _22544_, _04444_);
  nor _73537_ (_22546_, _12282_, _09462_);
  nor _73538_ (_22547_, _22546_, _22534_);
  nor _73539_ (_22548_, _22547_, _04444_);
  or _73540_ (_22549_, _22548_, _22545_);
  and _73541_ (_22551_, _22549_, _03983_);
  nor _73542_ (_22552_, _09462_, _05026_);
  nor _73543_ (_22553_, _22552_, _22534_);
  nor _73544_ (_22554_, _22553_, _03983_);
  nor _73545_ (_22555_, _22554_, _22551_);
  nor _73546_ (_22556_, _22555_, _03575_);
  or _73547_ (_22557_, _22556_, _07314_);
  nor _73548_ (_22558_, _22557_, _22541_);
  and _73549_ (_22559_, _22553_, _07314_);
  nor _73550_ (_22560_, _22559_, _22558_);
  nor _73551_ (_22562_, _22560_, _03479_);
  and _73552_ (_22563_, _06718_, _05254_);
  nor _73553_ (_22564_, _22534_, _06044_);
  not _73554_ (_22565_, _22564_);
  nor _73555_ (_22566_, _22565_, _22563_);
  nor _73556_ (_22567_, _22566_, _22562_);
  nor _73557_ (_22568_, _22567_, _03221_);
  nor _73558_ (_22569_, _12384_, _09462_);
  or _73559_ (_22570_, _22534_, _03474_);
  nor _73560_ (_22571_, _22570_, _22569_);
  or _73561_ (_22573_, _22571_, _03437_);
  nor _73562_ (_22574_, _22573_, _22568_);
  and _73563_ (_22575_, _05254_, _06261_);
  nor _73564_ (_22576_, _22575_, _22534_);
  nor _73565_ (_22577_, _22576_, _03438_);
  or _73566_ (_22578_, _22577_, _22574_);
  and _73567_ (_22579_, _22578_, _04499_);
  and _73568_ (_22580_, _12273_, _05254_);
  nor _73569_ (_22581_, _22580_, _22534_);
  nor _73570_ (_22582_, _22581_, _04499_);
  or _73571_ (_22584_, _22582_, _22579_);
  nor _73572_ (_22585_, _22584_, _03769_);
  and _73573_ (_22586_, _12401_, _05254_);
  or _73574_ (_22587_, _22534_, _04501_);
  nor _73575_ (_22588_, _22587_, _22586_);
  or _73576_ (_22589_, _22588_, _04504_);
  nor _73577_ (_22590_, _22589_, _22585_);
  nor _73578_ (_22591_, _22534_, _05665_);
  or _73579_ (_22592_, _22576_, _04505_);
  nor _73580_ (_22593_, _22592_, _22591_);
  nor _73581_ (_22595_, _22593_, _22590_);
  nor _73582_ (_22596_, _22595_, _03752_);
  or _73583_ (_22597_, _22591_, _03753_);
  or _73584_ (_22598_, _22597_, _22540_);
  and _73585_ (_22599_, _22598_, _03759_);
  not _73586_ (_22600_, _22599_);
  nor _73587_ (_22601_, _22600_, _22596_);
  nor _73588_ (_22602_, _12272_, _09462_);
  or _73589_ (_22603_, _22534_, _03759_);
  nor _73590_ (_22604_, _22603_, _22602_);
  or _73591_ (_22606_, _22604_, _03760_);
  nor _73592_ (_22607_, _22606_, _22601_);
  nor _73593_ (_22608_, _22607_, _22537_);
  nor _73594_ (_22609_, _22608_, _03790_);
  nor _73595_ (_22610_, _22547_, _04192_);
  or _73596_ (_22611_, _22610_, _03520_);
  nor _73597_ (_22612_, _22611_, _22609_);
  and _73598_ (_22613_, _12456_, _05254_);
  or _73599_ (_22614_, _22534_, _03521_);
  nor _73600_ (_22615_, _22614_, _22613_);
  nor _73601_ (_22617_, _22615_, _22612_);
  or _73602_ (_22618_, _22617_, _42967_);
  or _73603_ (_22619_, _42963_, \oc8051_golden_model_1.TMOD [2]);
  and _73604_ (_22620_, _22619_, _41755_);
  and _73605_ (_43284_, _22620_, _22618_);
  not _73606_ (_22621_, \oc8051_golden_model_1.TMOD [3]);
  nor _73607_ (_22622_, _05254_, _22621_);
  and _73608_ (_22623_, _06717_, _05254_);
  nor _73609_ (_22624_, _22623_, _22622_);
  or _73610_ (_22625_, _22624_, _06044_);
  and _73611_ (_22627_, _05254_, \oc8051_golden_model_1.ACC [3]);
  nor _73612_ (_22628_, _22627_, _22622_);
  nor _73613_ (_22629_, _22628_, _04427_);
  nor _73614_ (_22630_, _04426_, _22621_);
  or _73615_ (_22631_, _22630_, _22629_);
  and _73616_ (_22632_, _22631_, _04444_);
  nor _73617_ (_22633_, _12486_, _09462_);
  nor _73618_ (_22634_, _22633_, _22622_);
  nor _73619_ (_22635_, _22634_, _04444_);
  or _73620_ (_22636_, _22635_, _22632_);
  and _73621_ (_22638_, _22636_, _03983_);
  nor _73622_ (_22639_, _09462_, _04843_);
  nor _73623_ (_22640_, _22639_, _22622_);
  nor _73624_ (_22641_, _22640_, _03983_);
  nor _73625_ (_22642_, _22641_, _22638_);
  nor _73626_ (_22643_, _22642_, _03575_);
  nor _73627_ (_22644_, _22628_, _03583_);
  nor _73628_ (_22645_, _22644_, _07314_);
  not _73629_ (_22646_, _22645_);
  nor _73630_ (_22647_, _22646_, _22643_);
  and _73631_ (_22649_, _22640_, _07314_);
  or _73632_ (_22650_, _22649_, _03479_);
  or _73633_ (_22651_, _22650_, _22647_);
  and _73634_ (_22652_, _22651_, _03474_);
  and _73635_ (_22653_, _22652_, _22625_);
  nor _73636_ (_22654_, _12583_, _09462_);
  or _73637_ (_22655_, _22622_, _03474_);
  nor _73638_ (_22656_, _22655_, _22654_);
  or _73639_ (_22657_, _22656_, _03437_);
  nor _73640_ (_22658_, _22657_, _22653_);
  and _73641_ (_22660_, _05254_, _06217_);
  nor _73642_ (_22661_, _22660_, _22622_);
  nor _73643_ (_22662_, _22661_, _03438_);
  or _73644_ (_22663_, _22662_, _22658_);
  and _73645_ (_22664_, _22663_, _04499_);
  and _73646_ (_22665_, _12598_, _05254_);
  nor _73647_ (_22666_, _22665_, _22622_);
  nor _73648_ (_22667_, _22666_, _04499_);
  or _73649_ (_22668_, _22667_, _22664_);
  nor _73650_ (_22669_, _22668_, _03769_);
  and _73651_ (_22671_, _12604_, _05254_);
  or _73652_ (_22672_, _22622_, _04501_);
  nor _73653_ (_22673_, _22672_, _22671_);
  or _73654_ (_22674_, _22673_, _04504_);
  nor _73655_ (_22675_, _22674_, _22669_);
  nor _73656_ (_22676_, _22622_, _05521_);
  or _73657_ (_22677_, _22661_, _04505_);
  nor _73658_ (_22678_, _22677_, _22676_);
  nor _73659_ (_22679_, _22678_, _22675_);
  nor _73660_ (_22680_, _22679_, _03752_);
  or _73661_ (_22682_, _22676_, _03753_);
  nor _73662_ (_22683_, _22682_, _22628_);
  or _73663_ (_22684_, _22683_, _22680_);
  and _73664_ (_22685_, _22684_, _03759_);
  nor _73665_ (_22686_, _12597_, _09462_);
  nor _73666_ (_22687_, _22686_, _22622_);
  nor _73667_ (_22688_, _22687_, _03759_);
  or _73668_ (_22689_, _22688_, _22685_);
  and _73669_ (_22690_, _22689_, _04517_);
  nor _73670_ (_22691_, _12603_, _09462_);
  nor _73671_ (_22693_, _22691_, _22622_);
  nor _73672_ (_22694_, _22693_, _04517_);
  or _73673_ (_22695_, _22694_, _03790_);
  nor _73674_ (_22696_, _22695_, _22690_);
  and _73675_ (_22697_, _22634_, _03790_);
  or _73676_ (_22698_, _22697_, _03520_);
  nor _73677_ (_22699_, _22698_, _22696_);
  and _73678_ (_22700_, _12658_, _05254_);
  nor _73679_ (_22701_, _22700_, _22622_);
  nor _73680_ (_22702_, _22701_, _03521_);
  or _73681_ (_22704_, _22702_, _22699_);
  or _73682_ (_22705_, _22704_, _42967_);
  or _73683_ (_22706_, _42963_, \oc8051_golden_model_1.TMOD [3]);
  and _73684_ (_22707_, _22706_, _41755_);
  and _73685_ (_43285_, _22707_, _22705_);
  not _73686_ (_22708_, \oc8051_golden_model_1.TMOD [4]);
  nor _73687_ (_22709_, _05254_, _22708_);
  and _73688_ (_22710_, _12844_, _05254_);
  nor _73689_ (_22711_, _22710_, _22709_);
  nor _73690_ (_22712_, _22711_, _04501_);
  and _73691_ (_22714_, _05254_, \oc8051_golden_model_1.ACC [4]);
  nor _73692_ (_22715_, _22714_, _22709_);
  nor _73693_ (_22716_, _22715_, _04427_);
  nor _73694_ (_22717_, _04426_, _22708_);
  or _73695_ (_22718_, _22717_, _22716_);
  and _73696_ (_22719_, _22718_, _04444_);
  nor _73697_ (_22720_, _12733_, _09462_);
  nor _73698_ (_22721_, _22720_, _22709_);
  nor _73699_ (_22722_, _22721_, _04444_);
  or _73700_ (_22723_, _22722_, _22719_);
  and _73701_ (_22725_, _22723_, _03983_);
  nor _73702_ (_22726_, _05712_, _09462_);
  nor _73703_ (_22727_, _22726_, _22709_);
  nor _73704_ (_22728_, _22727_, _03983_);
  nor _73705_ (_22729_, _22728_, _22725_);
  nor _73706_ (_22730_, _22729_, _03575_);
  nor _73707_ (_22731_, _22715_, _03583_);
  nor _73708_ (_22732_, _22731_, _07314_);
  not _73709_ (_22733_, _22732_);
  nor _73710_ (_22734_, _22733_, _22730_);
  and _73711_ (_22736_, _22727_, _07314_);
  or _73712_ (_22737_, _22736_, _03479_);
  nor _73713_ (_22738_, _22737_, _22734_);
  and _73714_ (_22739_, _06722_, _05254_);
  or _73715_ (_22740_, _22739_, _22709_);
  and _73716_ (_22741_, _22740_, _03479_);
  or _73717_ (_22742_, _22741_, _03221_);
  or _73718_ (_22743_, _22742_, _22738_);
  nor _73719_ (_22744_, _12827_, _09462_);
  or _73720_ (_22745_, _22709_, _03474_);
  or _73721_ (_22747_, _22745_, _22744_);
  and _73722_ (_22748_, _22747_, _03438_);
  and _73723_ (_22749_, _22748_, _22743_);
  and _73724_ (_22750_, _06233_, _05254_);
  nor _73725_ (_22751_, _22750_, _22709_);
  nor _73726_ (_22752_, _22751_, _03438_);
  or _73727_ (_22753_, _22752_, _03636_);
  nor _73728_ (_22754_, _22753_, _22749_);
  and _73729_ (_22755_, _12711_, _05254_);
  or _73730_ (_22756_, _22709_, _04499_);
  nor _73731_ (_22758_, _22756_, _22755_);
  or _73732_ (_22759_, _22758_, _03769_);
  nor _73733_ (_22760_, _22759_, _22754_);
  nor _73734_ (_22761_, _22760_, _22712_);
  nor _73735_ (_22762_, _22761_, _04504_);
  not _73736_ (_22763_, _22709_);
  and _73737_ (_22764_, _22763_, _05760_);
  or _73738_ (_22765_, _22751_, _04505_);
  nor _73739_ (_22766_, _22765_, _22764_);
  nor _73740_ (_22767_, _22766_, _22762_);
  nor _73741_ (_22769_, _22767_, _03752_);
  or _73742_ (_22770_, _22764_, _03753_);
  or _73743_ (_22771_, _22770_, _22715_);
  and _73744_ (_22772_, _22771_, _03759_);
  not _73745_ (_22773_, _22772_);
  nor _73746_ (_22774_, _22773_, _22769_);
  nor _73747_ (_22775_, _12710_, _09462_);
  or _73748_ (_22776_, _22709_, _03759_);
  nor _73749_ (_22777_, _22776_, _22775_);
  or _73750_ (_22778_, _22777_, _03760_);
  nor _73751_ (_22780_, _22778_, _22774_);
  nor _73752_ (_22781_, _12843_, _09462_);
  nor _73753_ (_22782_, _22781_, _22709_);
  nor _73754_ (_22783_, _22782_, _04517_);
  or _73755_ (_22784_, _22783_, _03790_);
  nor _73756_ (_22785_, _22784_, _22780_);
  and _73757_ (_22786_, _22721_, _03790_);
  or _73758_ (_22787_, _22786_, _03520_);
  nor _73759_ (_22788_, _22787_, _22785_);
  and _73760_ (_22789_, _12893_, _05254_);
  nor _73761_ (_22791_, _22789_, _22709_);
  nor _73762_ (_22792_, _22791_, _03521_);
  or _73763_ (_22793_, _22792_, _22788_);
  or _73764_ (_22794_, _22793_, _42967_);
  or _73765_ (_22795_, _42963_, \oc8051_golden_model_1.TMOD [4]);
  and _73766_ (_22796_, _22795_, _41755_);
  and _73767_ (_43286_, _22796_, _22794_);
  not _73768_ (_22797_, \oc8051_golden_model_1.TMOD [5]);
  nor _73769_ (_22798_, _05254_, _22797_);
  and _73770_ (_22799_, _13042_, _05254_);
  nor _73771_ (_22801_, _22799_, _22798_);
  nor _73772_ (_22802_, _22801_, _04501_);
  nor _73773_ (_22803_, _05422_, _09462_);
  nor _73774_ (_22804_, _22803_, _22798_);
  and _73775_ (_22805_, _22804_, _07314_);
  and _73776_ (_22806_, _05254_, \oc8051_golden_model_1.ACC [5]);
  nor _73777_ (_22807_, _22806_, _22798_);
  nor _73778_ (_22808_, _22807_, _04427_);
  nor _73779_ (_22809_, _04426_, _22797_);
  or _73780_ (_22810_, _22809_, _22808_);
  and _73781_ (_22812_, _22810_, _04444_);
  nor _73782_ (_22813_, _12930_, _09462_);
  nor _73783_ (_22814_, _22813_, _22798_);
  nor _73784_ (_22815_, _22814_, _04444_);
  or _73785_ (_22816_, _22815_, _22812_);
  and _73786_ (_22817_, _22816_, _03983_);
  nor _73787_ (_22818_, _22804_, _03983_);
  nor _73788_ (_22819_, _22818_, _22817_);
  nor _73789_ (_22820_, _22819_, _03575_);
  nor _73790_ (_22821_, _22807_, _03583_);
  nor _73791_ (_22823_, _22821_, _07314_);
  not _73792_ (_22824_, _22823_);
  nor _73793_ (_22825_, _22824_, _22820_);
  nor _73794_ (_22826_, _22825_, _22805_);
  nor _73795_ (_22827_, _22826_, _03479_);
  and _73796_ (_22828_, _06721_, _05254_);
  nor _73797_ (_22829_, _22798_, _06044_);
  not _73798_ (_22830_, _22829_);
  nor _73799_ (_22831_, _22830_, _22828_);
  or _73800_ (_22832_, _22831_, _03221_);
  nor _73801_ (_22834_, _22832_, _22827_);
  nor _73802_ (_22835_, _13021_, _09462_);
  nor _73803_ (_22836_, _22835_, _22798_);
  nor _73804_ (_22837_, _22836_, _03474_);
  or _73805_ (_22838_, _22837_, _03437_);
  or _73806_ (_22839_, _22838_, _22834_);
  and _73807_ (_22840_, _06211_, _05254_);
  nor _73808_ (_22841_, _22840_, _22798_);
  nand _73809_ (_22842_, _22841_, _03437_);
  and _73810_ (_22843_, _22842_, _22839_);
  nor _73811_ (_22845_, _22843_, _03636_);
  and _73812_ (_22846_, _13036_, _05254_);
  or _73813_ (_22847_, _22798_, _04499_);
  nor _73814_ (_22848_, _22847_, _22846_);
  or _73815_ (_22849_, _22848_, _03769_);
  nor _73816_ (_22850_, _22849_, _22845_);
  nor _73817_ (_22851_, _22850_, _22802_);
  nor _73818_ (_22852_, _22851_, _04504_);
  not _73819_ (_22853_, _22798_);
  and _73820_ (_22854_, _22853_, _05471_);
  or _73821_ (_22856_, _22841_, _04505_);
  nor _73822_ (_22857_, _22856_, _22854_);
  nor _73823_ (_22858_, _22857_, _22852_);
  nor _73824_ (_22859_, _22858_, _03752_);
  or _73825_ (_22860_, _22854_, _03753_);
  nor _73826_ (_22861_, _22860_, _22807_);
  or _73827_ (_22862_, _22861_, _22859_);
  and _73828_ (_22863_, _22862_, _03759_);
  nor _73829_ (_22864_, _13035_, _09462_);
  nor _73830_ (_22865_, _22864_, _22798_);
  nor _73831_ (_22867_, _22865_, _03759_);
  or _73832_ (_22868_, _22867_, _22863_);
  and _73833_ (_22869_, _22868_, _04517_);
  nor _73834_ (_22870_, _13041_, _09462_);
  nor _73835_ (_22871_, _22870_, _22798_);
  nor _73836_ (_22872_, _22871_, _04517_);
  or _73837_ (_22873_, _22872_, _03790_);
  nor _73838_ (_22874_, _22873_, _22869_);
  and _73839_ (_22875_, _22814_, _03790_);
  or _73840_ (_22876_, _22875_, _03520_);
  nor _73841_ (_22878_, _22876_, _22874_);
  and _73842_ (_22879_, _13097_, _05254_);
  nor _73843_ (_22880_, _22879_, _22798_);
  nor _73844_ (_22881_, _22880_, _03521_);
  or _73845_ (_22882_, _22881_, _22878_);
  or _73846_ (_22883_, _22882_, _42967_);
  or _73847_ (_22884_, _42963_, \oc8051_golden_model_1.TMOD [5]);
  and _73848_ (_22885_, _22884_, _41755_);
  and _73849_ (_43287_, _22885_, _22883_);
  not _73850_ (_22886_, \oc8051_golden_model_1.TMOD [6]);
  nor _73851_ (_22888_, _05254_, _22886_);
  and _73852_ (_22889_, _13259_, _05254_);
  nor _73853_ (_22890_, _22889_, _22888_);
  nor _73854_ (_22891_, _22890_, _04501_);
  and _73855_ (_22892_, _05254_, \oc8051_golden_model_1.ACC [6]);
  nor _73856_ (_22893_, _22892_, _22888_);
  nor _73857_ (_22894_, _22893_, _03583_);
  nor _73858_ (_22895_, _22893_, _04427_);
  nor _73859_ (_22896_, _04426_, _22886_);
  or _73860_ (_22897_, _22896_, _22895_);
  and _73861_ (_22899_, _22897_, _04444_);
  nor _73862_ (_22900_, _13122_, _09462_);
  nor _73863_ (_22901_, _22900_, _22888_);
  nor _73864_ (_22902_, _22901_, _04444_);
  or _73865_ (_22903_, _22902_, _22899_);
  and _73866_ (_22904_, _22903_, _03983_);
  nor _73867_ (_22905_, _05327_, _09462_);
  nor _73868_ (_22906_, _22905_, _22888_);
  nor _73869_ (_22907_, _22906_, _03983_);
  nor _73870_ (_22908_, _22907_, _22904_);
  nor _73871_ (_22910_, _22908_, _03575_);
  or _73872_ (_22911_, _22910_, _07314_);
  nor _73873_ (_22912_, _22911_, _22894_);
  and _73874_ (_22913_, _22906_, _07314_);
  nor _73875_ (_22914_, _22913_, _22912_);
  nor _73876_ (_22915_, _22914_, _03479_);
  and _73877_ (_22916_, _06713_, _05254_);
  nor _73878_ (_22917_, _22888_, _06044_);
  not _73879_ (_22918_, _22917_);
  nor _73880_ (_22919_, _22918_, _22916_);
  or _73881_ (_22921_, _22919_, _03221_);
  nor _73882_ (_22922_, _22921_, _22915_);
  nor _73883_ (_22923_, _13237_, _09462_);
  nor _73884_ (_22924_, _22923_, _22888_);
  nor _73885_ (_22925_, _22924_, _03474_);
  or _73886_ (_22926_, _22925_, _03437_);
  or _73887_ (_22927_, _22926_, _22922_);
  and _73888_ (_22928_, _13244_, _05254_);
  nor _73889_ (_22929_, _22928_, _22888_);
  nand _73890_ (_22930_, _22929_, _03437_);
  and _73891_ (_22932_, _22930_, _22927_);
  nor _73892_ (_22933_, _22932_, _03636_);
  and _73893_ (_22934_, _13253_, _05254_);
  or _73894_ (_22935_, _22888_, _04499_);
  nor _73895_ (_22936_, _22935_, _22934_);
  or _73896_ (_22937_, _22936_, _03769_);
  nor _73897_ (_22938_, _22937_, _22933_);
  nor _73898_ (_22939_, _22938_, _22891_);
  nor _73899_ (_22940_, _22939_, _04504_);
  not _73900_ (_22941_, _22888_);
  and _73901_ (_22943_, _22941_, _05376_);
  or _73902_ (_22944_, _22929_, _04505_);
  nor _73903_ (_22945_, _22944_, _22943_);
  nor _73904_ (_22946_, _22945_, _22940_);
  nor _73905_ (_22947_, _22946_, _03752_);
  or _73906_ (_22948_, _22943_, _03753_);
  nor _73907_ (_22949_, _22948_, _22893_);
  or _73908_ (_22950_, _22949_, _22947_);
  and _73909_ (_22951_, _22950_, _03759_);
  nor _73910_ (_22952_, _13251_, _09462_);
  nor _73911_ (_22954_, _22952_, _22888_);
  nor _73912_ (_22955_, _22954_, _03759_);
  or _73913_ (_22956_, _22955_, _22951_);
  and _73914_ (_22957_, _22956_, _04517_);
  nor _73915_ (_22958_, _13258_, _09462_);
  nor _73916_ (_22959_, _22958_, _22888_);
  nor _73917_ (_22960_, _22959_, _04517_);
  or _73918_ (_22961_, _22960_, _03790_);
  nor _73919_ (_22962_, _22961_, _22957_);
  and _73920_ (_22963_, _22901_, _03790_);
  or _73921_ (_22965_, _22963_, _03520_);
  nor _73922_ (_22966_, _22965_, _22962_);
  and _73923_ (_22967_, _13312_, _05254_);
  nor _73924_ (_22968_, _22967_, _22888_);
  nor _73925_ (_22969_, _22968_, _03521_);
  or _73926_ (_22970_, _22969_, _22966_);
  or _73927_ (_22971_, _22970_, _42967_);
  or _73928_ (_22972_, _42963_, \oc8051_golden_model_1.TMOD [6]);
  and _73929_ (_22973_, _22972_, _41755_);
  and _73930_ (_43288_, _22973_, _22971_);
  not _73931_ (_22975_, \oc8051_golden_model_1.IE [0]);
  nor _73932_ (_22976_, _05193_, _22975_);
  and _73933_ (_22977_, _11995_, _05193_);
  nor _73934_ (_22978_, _22977_, _22976_);
  nor _73935_ (_22979_, _22978_, _04501_);
  and _73936_ (_22980_, _05941_, _05193_);
  nor _73937_ (_22981_, _22980_, _22976_);
  nor _73938_ (_22982_, _22981_, _04444_);
  nor _73939_ (_22983_, _04426_, _22975_);
  and _73940_ (_22984_, _05193_, \oc8051_golden_model_1.ACC [0]);
  nor _73941_ (_22986_, _22984_, _22976_);
  nor _73942_ (_22987_, _22986_, _04427_);
  nor _73943_ (_22988_, _22987_, _22983_);
  nor _73944_ (_22989_, _22988_, _03570_);
  or _73945_ (_22990_, _22989_, _03516_);
  nor _73946_ (_22991_, _22990_, _22982_);
  and _73947_ (_22992_, _11887_, _05807_);
  nor _73948_ (_22993_, _05807_, _22975_);
  or _73949_ (_22994_, _22993_, _03517_);
  nor _73950_ (_22995_, _22994_, _22992_);
  or _73951_ (_22996_, _22995_, _03568_);
  nor _73952_ (_22997_, _22996_, _22991_);
  and _73953_ (_22998_, _05193_, _04419_);
  nor _73954_ (_22999_, _22998_, _22976_);
  nor _73955_ (_23000_, _22999_, _03983_);
  or _73956_ (_23001_, _23000_, _22997_);
  and _73957_ (_23002_, _23001_, _03583_);
  nor _73958_ (_23003_, _22986_, _03583_);
  or _73959_ (_23004_, _23003_, _23002_);
  and _73960_ (_23005_, _23004_, _03513_);
  and _73961_ (_23008_, _22976_, _03512_);
  or _73962_ (_23009_, _23008_, _23005_);
  and _73963_ (_23010_, _23009_, _03506_);
  nor _73964_ (_23011_, _22981_, _03506_);
  or _73965_ (_23012_, _23011_, _23010_);
  and _73966_ (_23013_, _23012_, _03500_);
  nor _73967_ (_23014_, _11916_, _09570_);
  nor _73968_ (_23015_, _23014_, _22993_);
  nor _73969_ (_23016_, _23015_, _03500_);
  or _73970_ (_23017_, _23016_, _07314_);
  nor _73971_ (_23019_, _23017_, _23013_);
  and _73972_ (_23020_, _22999_, _07314_);
  or _73973_ (_23021_, _23020_, _03479_);
  nor _73974_ (_23022_, _23021_, _23019_);
  and _73975_ (_23023_, _06715_, _05193_);
  or _73976_ (_23024_, _23023_, _22976_);
  and _73977_ (_23025_, _23024_, _03479_);
  or _73978_ (_23026_, _23025_, _03221_);
  or _73979_ (_23027_, _23026_, _23022_);
  nor _73980_ (_23028_, _11975_, _09531_);
  or _73981_ (_23029_, _22976_, _03474_);
  or _73982_ (_23030_, _23029_, _23028_);
  and _73983_ (_23031_, _23030_, _03438_);
  and _73984_ (_23032_, _23031_, _23027_);
  and _73985_ (_23033_, _05193_, _06202_);
  nor _73986_ (_23034_, _23033_, _22976_);
  nor _73987_ (_23035_, _23034_, _03438_);
  or _73988_ (_23036_, _23035_, _03636_);
  nor _73989_ (_23037_, _23036_, _23032_);
  and _73990_ (_23038_, _11990_, _05193_);
  or _73991_ (_23041_, _22976_, _04499_);
  nor _73992_ (_23042_, _23041_, _23038_);
  or _73993_ (_23043_, _23042_, _03769_);
  nor _73994_ (_23044_, _23043_, _23037_);
  nor _73995_ (_23045_, _23044_, _22979_);
  nor _73996_ (_23046_, _23045_, _04504_);
  or _73997_ (_23047_, _23034_, _04505_);
  nor _73998_ (_23048_, _23047_, _22980_);
  nor _73999_ (_23049_, _23048_, _23046_);
  nor _74000_ (_23050_, _23049_, _03752_);
  and _74001_ (_23052_, _11994_, _05193_);
  or _74002_ (_23053_, _23052_, _22976_);
  and _74003_ (_23054_, _23053_, _03752_);
  or _74004_ (_23055_, _23054_, _23050_);
  and _74005_ (_23056_, _23055_, _03759_);
  nor _74006_ (_23057_, _11988_, _09531_);
  nor _74007_ (_23058_, _23057_, _22976_);
  nor _74008_ (_23059_, _23058_, _03759_);
  or _74009_ (_23060_, _23059_, _23056_);
  and _74010_ (_23061_, _23060_, _04517_);
  nor _74011_ (_23062_, _11870_, _09531_);
  nor _74012_ (_23063_, _23062_, _22976_);
  nor _74013_ (_23064_, _23063_, _04517_);
  or _74014_ (_23065_, _23064_, _23061_);
  and _74015_ (_23066_, _23065_, _04192_);
  nor _74016_ (_23067_, _22981_, _04192_);
  or _74017_ (_23068_, _23067_, _23066_);
  and _74018_ (_23069_, _23068_, _03152_);
  and _74019_ (_23070_, _22976_, _03151_);
  or _74020_ (_23071_, _23070_, _23069_);
  and _74021_ (_23074_, _23071_, _03521_);
  nor _74022_ (_23075_, _22981_, _03521_);
  or _74023_ (_23076_, _23075_, _23074_);
  or _74024_ (_23077_, _23076_, _42967_);
  or _74025_ (_23078_, _42963_, \oc8051_golden_model_1.IE [0]);
  and _74026_ (_23079_, _23078_, _41755_);
  and _74027_ (_43291_, _23079_, _23077_);
  or _74028_ (_23080_, _06714_, _09531_);
  nor _74029_ (_23081_, _05193_, \oc8051_golden_model_1.IE [1]);
  nor _74030_ (_23082_, _23081_, _06044_);
  and _74031_ (_23084_, _23082_, _23080_);
  not _74032_ (_23085_, \oc8051_golden_model_1.IE [1]);
  nor _74033_ (_23086_, _05193_, _23085_);
  nor _74034_ (_23087_, _09531_, _04603_);
  nor _74035_ (_23088_, _23087_, _23086_);
  nor _74036_ (_23089_, _23088_, _03983_);
  nor _74037_ (_23090_, _05807_, _23085_);
  and _74038_ (_23091_, _12083_, _05807_);
  nor _74039_ (_23092_, _23091_, _23090_);
  and _74040_ (_23093_, _23092_, _03516_);
  and _74041_ (_23094_, _12252_, _05193_);
  nor _74042_ (_23095_, _23094_, _23081_);
  and _74043_ (_23096_, _23095_, _03570_);
  and _74044_ (_23097_, _05193_, _03233_);
  nor _74045_ (_23098_, _23097_, _23081_);
  and _74046_ (_23099_, _23098_, _04426_);
  nor _74047_ (_23100_, _04426_, _23085_);
  nor _74048_ (_23101_, _23100_, _23099_);
  nor _74049_ (_23102_, _23101_, _03570_);
  or _74050_ (_23103_, _23102_, _03516_);
  nor _74051_ (_23106_, _23103_, _23096_);
  nor _74052_ (_23107_, _23106_, _23093_);
  and _74053_ (_23108_, _23107_, _03983_);
  or _74054_ (_23109_, _23108_, _23089_);
  and _74055_ (_23110_, _23109_, _03583_);
  and _74056_ (_23111_, _23098_, _03575_);
  or _74057_ (_23112_, _23111_, _23110_);
  and _74058_ (_23113_, _23112_, _03513_);
  and _74059_ (_23114_, _12069_, _05807_);
  nor _74060_ (_23115_, _23114_, _23090_);
  nor _74061_ (_23117_, _23115_, _03513_);
  or _74062_ (_23118_, _23117_, _03505_);
  or _74063_ (_23119_, _23118_, _23113_);
  nor _74064_ (_23120_, _23090_, _12098_);
  nor _74065_ (_23121_, _23120_, _23092_);
  or _74066_ (_23122_, _23121_, _03506_);
  and _74067_ (_23123_, _23122_, _03500_);
  and _74068_ (_23124_, _23123_, _23119_);
  nor _74069_ (_23125_, _12116_, _09570_);
  nor _74070_ (_23126_, _23125_, _23090_);
  nor _74071_ (_23127_, _23126_, _03500_);
  nor _74072_ (_23128_, _23127_, _07314_);
  not _74073_ (_23129_, _23128_);
  nor _74074_ (_23130_, _23129_, _23124_);
  and _74075_ (_23131_, _23088_, _07314_);
  or _74076_ (_23132_, _23131_, _03479_);
  nor _74077_ (_23133_, _23132_, _23130_);
  or _74078_ (_23134_, _23133_, _23084_);
  and _74079_ (_23135_, _23134_, _03474_);
  nor _74080_ (_23136_, _12176_, _09531_);
  or _74081_ (_23139_, _23136_, _23086_);
  and _74082_ (_23140_, _23139_, _03221_);
  nor _74083_ (_23141_, _23140_, _23135_);
  nor _74084_ (_23142_, _23141_, _03437_);
  and _74085_ (_23143_, _05193_, _04317_);
  not _74086_ (_23144_, _23143_);
  nor _74087_ (_23145_, _23081_, _03438_);
  and _74088_ (_23146_, _23145_, _23144_);
  nor _74089_ (_23147_, _23146_, _23142_);
  nor _74090_ (_23148_, _23147_, _03636_);
  not _74091_ (_23150_, _23081_);
  nor _74092_ (_23151_, _12191_, _09531_);
  nor _74093_ (_23152_, _23151_, _04499_);
  and _74094_ (_23153_, _23152_, _23150_);
  nor _74095_ (_23154_, _23153_, _23148_);
  nor _74096_ (_23155_, _23154_, _03769_);
  nor _74097_ (_23156_, _12197_, _09531_);
  nor _74098_ (_23157_, _23156_, _04501_);
  and _74099_ (_23158_, _23157_, _23150_);
  nor _74100_ (_23159_, _23158_, _23155_);
  nor _74101_ (_23160_, _23159_, _04504_);
  nor _74102_ (_23161_, _12190_, _09531_);
  nor _74103_ (_23162_, _23161_, _05769_);
  and _74104_ (_23163_, _23162_, _23150_);
  nor _74105_ (_23164_, _23163_, _23160_);
  nor _74106_ (_23165_, _23164_, _03752_);
  nor _74107_ (_23166_, _23086_, _05569_);
  nor _74108_ (_23167_, _23166_, _03753_);
  and _74109_ (_23168_, _23167_, _23098_);
  nor _74110_ (_23169_, _23168_, _23165_);
  nor _74111_ (_23171_, _23169_, _03758_);
  and _74112_ (_23172_, _23143_, _05940_);
  nor _74113_ (_23173_, _23172_, _03759_);
  and _74114_ (_23174_, _23173_, _23150_);
  nor _74115_ (_23175_, _23174_, _23171_);
  nor _74116_ (_23176_, _23175_, _03760_);
  and _74117_ (_23177_, _23097_, _05940_);
  nor _74118_ (_23178_, _23177_, _04517_);
  and _74119_ (_23179_, _23178_, _23150_);
  or _74120_ (_23180_, _23179_, _03790_);
  nor _74121_ (_23182_, _23180_, _23176_);
  nor _74122_ (_23183_, _23095_, _04192_);
  or _74123_ (_23184_, _23183_, _03151_);
  nor _74124_ (_23185_, _23184_, _23182_);
  nor _74125_ (_23186_, _23115_, _03152_);
  or _74126_ (_23187_, _23186_, _03520_);
  nor _74127_ (_23188_, _23187_, _23185_);
  or _74128_ (_23189_, _23086_, _03521_);
  nor _74129_ (_23190_, _23189_, _23094_);
  nor _74130_ (_23191_, _23190_, _23188_);
  or _74131_ (_23192_, _23191_, _42967_);
  or _74132_ (_23193_, _42963_, \oc8051_golden_model_1.IE [1]);
  and _74133_ (_23194_, _23193_, _41755_);
  and _74134_ (_43292_, _23194_, _23192_);
  not _74135_ (_23195_, \oc8051_golden_model_1.IE [2]);
  nor _74136_ (_23196_, _05193_, _23195_);
  and _74137_ (_23197_, _12401_, _05193_);
  nor _74138_ (_23198_, _23197_, _23196_);
  nor _74139_ (_23199_, _23198_, _04501_);
  nor _74140_ (_23200_, _09531_, _05026_);
  nor _74141_ (_23202_, _23200_, _23196_);
  and _74142_ (_23203_, _23202_, _07314_);
  and _74143_ (_23204_, _05193_, \oc8051_golden_model_1.ACC [2]);
  nor _74144_ (_23205_, _23204_, _23196_);
  nor _74145_ (_23206_, _23205_, _04427_);
  nor _74146_ (_23207_, _04426_, _23195_);
  or _74147_ (_23208_, _23207_, _23206_);
  and _74148_ (_23209_, _23208_, _04444_);
  nor _74149_ (_23210_, _12282_, _09531_);
  nor _74150_ (_23211_, _23210_, _23196_);
  nor _74151_ (_23212_, _23211_, _04444_);
  or _74152_ (_23213_, _23212_, _23209_);
  and _74153_ (_23214_, _23213_, _03517_);
  nor _74154_ (_23215_, _05807_, _23195_);
  and _74155_ (_23216_, _12278_, _05807_);
  nor _74156_ (_23217_, _23216_, _23215_);
  nor _74157_ (_23218_, _23217_, _03517_);
  or _74158_ (_23219_, _23218_, _23214_);
  and _74159_ (_23220_, _23219_, _03983_);
  nor _74160_ (_23221_, _23202_, _03983_);
  or _74161_ (_23222_, _23221_, _23220_);
  and _74162_ (_23223_, _23222_, _03583_);
  nor _74163_ (_23224_, _23205_, _03583_);
  or _74164_ (_23225_, _23224_, _23223_);
  and _74165_ (_23226_, _23225_, _03513_);
  and _74166_ (_23227_, _12276_, _05807_);
  nor _74167_ (_23228_, _23227_, _23215_);
  nor _74168_ (_23229_, _23228_, _03513_);
  or _74169_ (_23230_, _23229_, _03505_);
  or _74170_ (_23231_, _23230_, _23226_);
  and _74171_ (_23232_, _23216_, _12309_);
  or _74172_ (_23233_, _23215_, _03506_);
  or _74173_ (_23234_, _23233_, _23232_);
  and _74174_ (_23235_, _23234_, _03500_);
  and _74175_ (_23236_, _23235_, _23231_);
  nor _74176_ (_23237_, _12326_, _09570_);
  nor _74177_ (_23238_, _23237_, _23215_);
  nor _74178_ (_23239_, _23238_, _03500_);
  nor _74179_ (_23240_, _23239_, _07314_);
  not _74180_ (_23241_, _23240_);
  nor _74181_ (_23242_, _23241_, _23236_);
  nor _74182_ (_23243_, _23242_, _23203_);
  nor _74183_ (_23244_, _23243_, _03479_);
  and _74184_ (_23245_, _06718_, _05193_);
  nor _74185_ (_23246_, _23196_, _06044_);
  not _74186_ (_23247_, _23246_);
  nor _74187_ (_23248_, _23247_, _23245_);
  or _74188_ (_23249_, _23248_, _03221_);
  nor _74189_ (_23250_, _23249_, _23244_);
  nor _74190_ (_23251_, _12384_, _09531_);
  nor _74191_ (_23253_, _23251_, _23196_);
  nor _74192_ (_23254_, _23253_, _03474_);
  or _74193_ (_23255_, _23254_, _03437_);
  or _74194_ (_23256_, _23255_, _23250_);
  and _74195_ (_23257_, _05193_, _06261_);
  nor _74196_ (_23258_, _23257_, _23196_);
  nand _74197_ (_23259_, _23258_, _03437_);
  and _74198_ (_23260_, _23259_, _23256_);
  nor _74199_ (_23261_, _23260_, _03636_);
  and _74200_ (_23262_, _12273_, _05193_);
  or _74201_ (_23264_, _23196_, _04499_);
  nor _74202_ (_23265_, _23264_, _23262_);
  or _74203_ (_23266_, _23265_, _03769_);
  nor _74204_ (_23267_, _23266_, _23261_);
  nor _74205_ (_23268_, _23267_, _23199_);
  nor _74206_ (_23269_, _23268_, _04504_);
  not _74207_ (_23270_, _23196_);
  and _74208_ (_23271_, _23270_, _05664_);
  or _74209_ (_23272_, _23258_, _04505_);
  nor _74210_ (_23273_, _23272_, _23271_);
  nor _74211_ (_23274_, _23273_, _23269_);
  nor _74212_ (_23275_, _23274_, _03752_);
  or _74213_ (_23276_, _23271_, _03753_);
  nor _74214_ (_23277_, _23276_, _23205_);
  or _74215_ (_23278_, _23277_, _23275_);
  and _74216_ (_23279_, _23278_, _03759_);
  nor _74217_ (_23280_, _12272_, _09531_);
  nor _74218_ (_23281_, _23280_, _23196_);
  nor _74219_ (_23282_, _23281_, _03759_);
  or _74220_ (_23283_, _23282_, _23279_);
  and _74221_ (_23285_, _23283_, _04517_);
  nor _74222_ (_23286_, _12400_, _09531_);
  nor _74223_ (_23287_, _23286_, _23196_);
  nor _74224_ (_23288_, _23287_, _04517_);
  or _74225_ (_23289_, _23288_, _23285_);
  and _74226_ (_23290_, _23289_, _04192_);
  nor _74227_ (_23291_, _23211_, _04192_);
  or _74228_ (_23292_, _23291_, _23290_);
  and _74229_ (_23293_, _23292_, _03152_);
  nor _74230_ (_23294_, _23228_, _03152_);
  or _74231_ (_23296_, _23294_, _23293_);
  and _74232_ (_23297_, _23296_, _03521_);
  and _74233_ (_23298_, _12456_, _05193_);
  nor _74234_ (_23299_, _23298_, _23196_);
  nor _74235_ (_23300_, _23299_, _03521_);
  or _74236_ (_23301_, _23300_, _23297_);
  or _74237_ (_23302_, _23301_, _42967_);
  or _74238_ (_23303_, _42963_, \oc8051_golden_model_1.IE [2]);
  and _74239_ (_23304_, _23303_, _41755_);
  and _74240_ (_43293_, _23304_, _23302_);
  not _74241_ (_23306_, \oc8051_golden_model_1.IE [3]);
  nor _74242_ (_23307_, _05193_, _23306_);
  and _74243_ (_23308_, _12604_, _05193_);
  nor _74244_ (_23309_, _23308_, _23307_);
  nor _74245_ (_23310_, _23309_, _04501_);
  nor _74246_ (_23311_, _09531_, _04843_);
  nor _74247_ (_23312_, _23311_, _23307_);
  and _74248_ (_23313_, _23312_, _07314_);
  and _74249_ (_23314_, _05193_, \oc8051_golden_model_1.ACC [3]);
  nor _74250_ (_23315_, _23314_, _23307_);
  nor _74251_ (_23317_, _23315_, _04427_);
  nor _74252_ (_23318_, _04426_, _23306_);
  or _74253_ (_23319_, _23318_, _23317_);
  and _74254_ (_23320_, _23319_, _04444_);
  nor _74255_ (_23321_, _12486_, _09531_);
  nor _74256_ (_23322_, _23321_, _23307_);
  nor _74257_ (_23323_, _23322_, _04444_);
  or _74258_ (_23324_, _23323_, _23320_);
  and _74259_ (_23325_, _23324_, _03517_);
  nor _74260_ (_23326_, _05807_, _23306_);
  and _74261_ (_23327_, _12490_, _05807_);
  nor _74262_ (_23328_, _23327_, _23326_);
  nor _74263_ (_23329_, _23328_, _03517_);
  or _74264_ (_23330_, _23329_, _03568_);
  or _74265_ (_23331_, _23330_, _23325_);
  nand _74266_ (_23332_, _23312_, _03568_);
  and _74267_ (_23333_, _23332_, _23331_);
  and _74268_ (_23334_, _23333_, _03583_);
  nor _74269_ (_23335_, _23315_, _03583_);
  or _74270_ (_23336_, _23335_, _23334_);
  and _74271_ (_23338_, _23336_, _03513_);
  and _74272_ (_23339_, _12500_, _05807_);
  nor _74273_ (_23340_, _23339_, _23326_);
  nor _74274_ (_23341_, _23340_, _03513_);
  or _74275_ (_23342_, _23341_, _03505_);
  or _74276_ (_23343_, _23342_, _23338_);
  nor _74277_ (_23344_, _23326_, _12507_);
  nor _74278_ (_23345_, _23344_, _23328_);
  or _74279_ (_23346_, _23345_, _03506_);
  and _74280_ (_23347_, _23346_, _03500_);
  and _74281_ (_23349_, _23347_, _23343_);
  nor _74282_ (_23350_, _12525_, _09570_);
  nor _74283_ (_23351_, _23350_, _23326_);
  nor _74284_ (_23352_, _23351_, _03500_);
  nor _74285_ (_23353_, _23352_, _07314_);
  not _74286_ (_23354_, _23353_);
  nor _74287_ (_23355_, _23354_, _23349_);
  nor _74288_ (_23356_, _23355_, _23313_);
  nor _74289_ (_23357_, _23356_, _03479_);
  and _74290_ (_23358_, _06717_, _05193_);
  nor _74291_ (_23360_, _23307_, _06044_);
  not _74292_ (_23361_, _23360_);
  nor _74293_ (_23362_, _23361_, _23358_);
  or _74294_ (_23363_, _23362_, _03221_);
  nor _74295_ (_23364_, _23363_, _23357_);
  nor _74296_ (_23365_, _12583_, _09531_);
  nor _74297_ (_23366_, _23365_, _23307_);
  nor _74298_ (_23367_, _23366_, _03474_);
  or _74299_ (_23368_, _23367_, _03437_);
  or _74300_ (_23369_, _23368_, _23364_);
  and _74301_ (_23371_, _05193_, _06217_);
  nor _74302_ (_23372_, _23371_, _23307_);
  nand _74303_ (_23373_, _23372_, _03437_);
  and _74304_ (_23374_, _23373_, _23369_);
  nor _74305_ (_23375_, _23374_, _03636_);
  and _74306_ (_23376_, _12598_, _05193_);
  or _74307_ (_23377_, _23307_, _04499_);
  nor _74308_ (_23378_, _23377_, _23376_);
  or _74309_ (_23379_, _23378_, _03769_);
  nor _74310_ (_23380_, _23379_, _23375_);
  nor _74311_ (_23382_, _23380_, _23310_);
  nor _74312_ (_23383_, _23382_, _04504_);
  not _74313_ (_23384_, _23307_);
  and _74314_ (_23385_, _23384_, _05520_);
  or _74315_ (_23386_, _23372_, _04505_);
  nor _74316_ (_23387_, _23386_, _23385_);
  nor _74317_ (_23388_, _23387_, _23383_);
  nor _74318_ (_23389_, _23388_, _03752_);
  or _74319_ (_23390_, _23385_, _03753_);
  or _74320_ (_23391_, _23390_, _23315_);
  and _74321_ (_23392_, _23391_, _03759_);
  not _74322_ (_23393_, _23392_);
  nor _74323_ (_23394_, _23393_, _23389_);
  nor _74324_ (_23395_, _12597_, _09531_);
  or _74325_ (_23396_, _23307_, _03759_);
  nor _74326_ (_23397_, _23396_, _23395_);
  or _74327_ (_23398_, _23397_, _03760_);
  nor _74328_ (_23399_, _23398_, _23394_);
  nor _74329_ (_23400_, _12603_, _09531_);
  nor _74330_ (_23401_, _23400_, _23307_);
  nor _74331_ (_23403_, _23401_, _04517_);
  or _74332_ (_23404_, _23403_, _23399_);
  and _74333_ (_23405_, _23404_, _04192_);
  nor _74334_ (_23406_, _23322_, _04192_);
  or _74335_ (_23407_, _23406_, _23405_);
  and _74336_ (_23408_, _23407_, _03152_);
  nor _74337_ (_23409_, _23340_, _03152_);
  or _74338_ (_23410_, _23409_, _23408_);
  and _74339_ (_23411_, _23410_, _03521_);
  and _74340_ (_23412_, _12658_, _05193_);
  nor _74341_ (_23414_, _23412_, _23307_);
  nor _74342_ (_23415_, _23414_, _03521_);
  or _74343_ (_23416_, _23415_, _23411_);
  or _74344_ (_23417_, _23416_, _42967_);
  or _74345_ (_23418_, _42963_, \oc8051_golden_model_1.IE [3]);
  and _74346_ (_23419_, _23418_, _41755_);
  and _74347_ (_43294_, _23419_, _23417_);
  not _74348_ (_23420_, \oc8051_golden_model_1.IE [4]);
  nor _74349_ (_23421_, _05193_, _23420_);
  and _74350_ (_23422_, _12844_, _05193_);
  nor _74351_ (_23424_, _23422_, _23421_);
  nor _74352_ (_23425_, _23424_, _04501_);
  nor _74353_ (_23426_, _05712_, _09531_);
  nor _74354_ (_23427_, _23426_, _23421_);
  and _74355_ (_23428_, _23427_, _07314_);
  and _74356_ (_23429_, _05193_, \oc8051_golden_model_1.ACC [4]);
  nor _74357_ (_23430_, _23429_, _23421_);
  nor _74358_ (_23431_, _23430_, _04427_);
  nor _74359_ (_23432_, _04426_, _23420_);
  or _74360_ (_23433_, _23432_, _23431_);
  and _74361_ (_23435_, _23433_, _04444_);
  nor _74362_ (_23436_, _12733_, _09531_);
  nor _74363_ (_23437_, _23436_, _23421_);
  nor _74364_ (_23438_, _23437_, _04444_);
  or _74365_ (_23439_, _23438_, _23435_);
  and _74366_ (_23440_, _23439_, _03517_);
  nor _74367_ (_23441_, _05807_, _23420_);
  and _74368_ (_23442_, _12737_, _05807_);
  nor _74369_ (_23443_, _23442_, _23441_);
  nor _74370_ (_23444_, _23443_, _03517_);
  or _74371_ (_23446_, _23444_, _03568_);
  or _74372_ (_23447_, _23446_, _23440_);
  nand _74373_ (_23448_, _23427_, _03568_);
  and _74374_ (_23449_, _23448_, _23447_);
  and _74375_ (_23450_, _23449_, _03583_);
  nor _74376_ (_23451_, _23430_, _03583_);
  or _74377_ (_23452_, _23451_, _23450_);
  and _74378_ (_23453_, _23452_, _03513_);
  and _74379_ (_23454_, _12718_, _05807_);
  nor _74380_ (_23455_, _23454_, _23441_);
  nor _74381_ (_23456_, _23455_, _03513_);
  or _74382_ (_23457_, _23456_, _03505_);
  or _74383_ (_23458_, _23457_, _23453_);
  nor _74384_ (_23459_, _23441_, _12752_);
  nor _74385_ (_23460_, _23459_, _23443_);
  or _74386_ (_23461_, _23460_, _03506_);
  and _74387_ (_23462_, _23461_, _03500_);
  and _74388_ (_23463_, _23462_, _23458_);
  nor _74389_ (_23464_, _12716_, _09570_);
  nor _74390_ (_23465_, _23464_, _23441_);
  nor _74391_ (_23467_, _23465_, _03500_);
  nor _74392_ (_23468_, _23467_, _07314_);
  not _74393_ (_23469_, _23468_);
  nor _74394_ (_23470_, _23469_, _23463_);
  nor _74395_ (_23471_, _23470_, _23428_);
  nor _74396_ (_23472_, _23471_, _03479_);
  and _74397_ (_23473_, _06722_, _05193_);
  nor _74398_ (_23474_, _23421_, _06044_);
  not _74399_ (_23475_, _23474_);
  nor _74400_ (_23476_, _23475_, _23473_);
  or _74401_ (_23478_, _23476_, _03221_);
  nor _74402_ (_23479_, _23478_, _23472_);
  nor _74403_ (_23480_, _12827_, _09531_);
  nor _74404_ (_23481_, _23480_, _23421_);
  nor _74405_ (_23482_, _23481_, _03474_);
  or _74406_ (_23483_, _23482_, _03437_);
  or _74407_ (_23484_, _23483_, _23479_);
  and _74408_ (_23485_, _06233_, _05193_);
  nor _74409_ (_23486_, _23485_, _23421_);
  nand _74410_ (_23487_, _23486_, _03437_);
  and _74411_ (_23489_, _23487_, _23484_);
  nor _74412_ (_23490_, _23489_, _03636_);
  and _74413_ (_23491_, _12711_, _05193_);
  or _74414_ (_23492_, _23421_, _04499_);
  nor _74415_ (_23493_, _23492_, _23491_);
  or _74416_ (_23494_, _23493_, _03769_);
  nor _74417_ (_23495_, _23494_, _23490_);
  nor _74418_ (_23496_, _23495_, _23425_);
  nor _74419_ (_23497_, _23496_, _04504_);
  not _74420_ (_23498_, _23421_);
  and _74421_ (_23500_, _23498_, _05760_);
  or _74422_ (_23501_, _23486_, _04505_);
  nor _74423_ (_23502_, _23501_, _23500_);
  nor _74424_ (_23503_, _23502_, _23497_);
  nor _74425_ (_23504_, _23503_, _03752_);
  or _74426_ (_23505_, _23500_, _03753_);
  nor _74427_ (_23506_, _23505_, _23430_);
  or _74428_ (_23507_, _23506_, _23504_);
  and _74429_ (_23508_, _23507_, _03759_);
  nor _74430_ (_23509_, _12710_, _09531_);
  nor _74431_ (_23511_, _23509_, _23421_);
  nor _74432_ (_23512_, _23511_, _03759_);
  or _74433_ (_23513_, _23512_, _23508_);
  and _74434_ (_23514_, _23513_, _04517_);
  nor _74435_ (_23515_, _12843_, _09531_);
  nor _74436_ (_23516_, _23515_, _23421_);
  nor _74437_ (_23517_, _23516_, _04517_);
  or _74438_ (_23518_, _23517_, _23514_);
  and _74439_ (_23519_, _23518_, _04192_);
  nor _74440_ (_23520_, _23437_, _04192_);
  or _74441_ (_23521_, _23520_, _23519_);
  and _74442_ (_23522_, _23521_, _03152_);
  nor _74443_ (_23523_, _23455_, _03152_);
  or _74444_ (_23524_, _23523_, _23522_);
  and _74445_ (_23525_, _23524_, _03521_);
  and _74446_ (_23526_, _12893_, _05193_);
  nor _74447_ (_23527_, _23526_, _23421_);
  nor _74448_ (_23528_, _23527_, _03521_);
  or _74449_ (_23529_, _23528_, _23525_);
  or _74450_ (_23530_, _23529_, _42967_);
  or _74451_ (_23532_, _42963_, \oc8051_golden_model_1.IE [4]);
  and _74452_ (_23533_, _23532_, _41755_);
  and _74453_ (_43295_, _23533_, _23530_);
  not _74454_ (_23534_, \oc8051_golden_model_1.IE [5]);
  nor _74455_ (_23535_, _05193_, _23534_);
  and _74456_ (_23536_, _13042_, _05193_);
  nor _74457_ (_23537_, _23536_, _23535_);
  nor _74458_ (_23538_, _23537_, _04501_);
  nor _74459_ (_23539_, _05422_, _09531_);
  nor _74460_ (_23540_, _23539_, _23535_);
  and _74461_ (_23542_, _23540_, _07314_);
  and _74462_ (_23543_, _05193_, \oc8051_golden_model_1.ACC [5]);
  nor _74463_ (_23544_, _23543_, _23535_);
  nor _74464_ (_23545_, _23544_, _04427_);
  nor _74465_ (_23546_, _04426_, _23534_);
  or _74466_ (_23547_, _23546_, _23545_);
  and _74467_ (_23548_, _23547_, _04444_);
  nor _74468_ (_23549_, _12930_, _09531_);
  nor _74469_ (_23550_, _23549_, _23535_);
  nor _74470_ (_23551_, _23550_, _04444_);
  or _74471_ (_23553_, _23551_, _23548_);
  and _74472_ (_23554_, _23553_, _03517_);
  nor _74473_ (_23555_, _05807_, _23534_);
  and _74474_ (_23556_, _12934_, _05807_);
  nor _74475_ (_23557_, _23556_, _23555_);
  nor _74476_ (_23558_, _23557_, _03517_);
  or _74477_ (_23559_, _23558_, _03568_);
  or _74478_ (_23560_, _23559_, _23554_);
  nand _74479_ (_23561_, _23540_, _03568_);
  and _74480_ (_23562_, _23561_, _23560_);
  and _74481_ (_23564_, _23562_, _03583_);
  nor _74482_ (_23565_, _23544_, _03583_);
  or _74483_ (_23566_, _23565_, _23564_);
  and _74484_ (_23567_, _23566_, _03513_);
  and _74485_ (_23568_, _12914_, _05807_);
  nor _74486_ (_23569_, _23568_, _23555_);
  nor _74487_ (_23570_, _23569_, _03513_);
  or _74488_ (_23571_, _23570_, _03505_);
  or _74489_ (_23572_, _23571_, _23567_);
  nor _74490_ (_23573_, _23555_, _12949_);
  nor _74491_ (_23575_, _23573_, _23557_);
  or _74492_ (_23576_, _23575_, _03506_);
  and _74493_ (_23577_, _23576_, _03500_);
  and _74494_ (_23578_, _23577_, _23572_);
  nor _74495_ (_23579_, _12912_, _09570_);
  nor _74496_ (_23580_, _23579_, _23555_);
  nor _74497_ (_23581_, _23580_, _03500_);
  nor _74498_ (_23582_, _23581_, _07314_);
  not _74499_ (_23583_, _23582_);
  nor _74500_ (_23584_, _23583_, _23578_);
  nor _74501_ (_23585_, _23584_, _23542_);
  nor _74502_ (_23586_, _23585_, _03479_);
  and _74503_ (_23587_, _06721_, _05193_);
  nor _74504_ (_23588_, _23535_, _06044_);
  not _74505_ (_23589_, _23588_);
  nor _74506_ (_23590_, _23589_, _23587_);
  or _74507_ (_23591_, _23590_, _03221_);
  nor _74508_ (_23592_, _23591_, _23586_);
  nor _74509_ (_23593_, _13021_, _09531_);
  nor _74510_ (_23594_, _23593_, _23535_);
  nor _74511_ (_23596_, _23594_, _03474_);
  or _74512_ (_23597_, _23596_, _03437_);
  or _74513_ (_23598_, _23597_, _23592_);
  and _74514_ (_23599_, _06211_, _05193_);
  nor _74515_ (_23600_, _23599_, _23535_);
  nand _74516_ (_23601_, _23600_, _03437_);
  and _74517_ (_23602_, _23601_, _23598_);
  nor _74518_ (_23603_, _23602_, _03636_);
  and _74519_ (_23604_, _13036_, _05193_);
  or _74520_ (_23605_, _23535_, _04499_);
  nor _74521_ (_23607_, _23605_, _23604_);
  or _74522_ (_23608_, _23607_, _03769_);
  nor _74523_ (_23609_, _23608_, _23603_);
  nor _74524_ (_23610_, _23609_, _23538_);
  nor _74525_ (_23611_, _23610_, _04504_);
  not _74526_ (_23612_, _23535_);
  and _74527_ (_23613_, _23612_, _05471_);
  or _74528_ (_23614_, _23600_, _04505_);
  nor _74529_ (_23615_, _23614_, _23613_);
  nor _74530_ (_23616_, _23615_, _23611_);
  nor _74531_ (_23618_, _23616_, _03752_);
  or _74532_ (_23619_, _23613_, _03753_);
  nor _74533_ (_23620_, _23619_, _23544_);
  or _74534_ (_23621_, _23620_, _23618_);
  and _74535_ (_23622_, _23621_, _03759_);
  nor _74536_ (_23623_, _13035_, _09531_);
  nor _74537_ (_23624_, _23623_, _23535_);
  nor _74538_ (_23625_, _23624_, _03759_);
  or _74539_ (_23626_, _23625_, _23622_);
  and _74540_ (_23627_, _23626_, _04517_);
  nor _74541_ (_23629_, _13041_, _09531_);
  nor _74542_ (_23630_, _23629_, _23535_);
  nor _74543_ (_23631_, _23630_, _04517_);
  or _74544_ (_23632_, _23631_, _23627_);
  and _74545_ (_23633_, _23632_, _04192_);
  nor _74546_ (_23634_, _23550_, _04192_);
  or _74547_ (_23635_, _23634_, _23633_);
  and _74548_ (_23636_, _23635_, _03152_);
  nor _74549_ (_23637_, _23569_, _03152_);
  or _74550_ (_23638_, _23637_, _23636_);
  and _74551_ (_23640_, _23638_, _03521_);
  and _74552_ (_23641_, _13097_, _05193_);
  nor _74553_ (_23642_, _23641_, _23535_);
  nor _74554_ (_23643_, _23642_, _03521_);
  or _74555_ (_23644_, _23643_, _23640_);
  or _74556_ (_23645_, _23644_, _42967_);
  or _74557_ (_23646_, _42963_, \oc8051_golden_model_1.IE [5]);
  and _74558_ (_23647_, _23646_, _41755_);
  and _74559_ (_43296_, _23647_, _23645_);
  not _74560_ (_23648_, \oc8051_golden_model_1.IE [6]);
  nor _74561_ (_23650_, _05193_, _23648_);
  and _74562_ (_23651_, _13259_, _05193_);
  nor _74563_ (_23652_, _23651_, _23650_);
  nor _74564_ (_23653_, _23652_, _04501_);
  nor _74565_ (_23654_, _05327_, _09531_);
  nor _74566_ (_23655_, _23654_, _23650_);
  and _74567_ (_23656_, _23655_, _07314_);
  and _74568_ (_23657_, _05193_, \oc8051_golden_model_1.ACC [6]);
  nor _74569_ (_23658_, _23657_, _23650_);
  nor _74570_ (_23659_, _23658_, _04427_);
  nor _74571_ (_23661_, _04426_, _23648_);
  or _74572_ (_23662_, _23661_, _23659_);
  and _74573_ (_23663_, _23662_, _04444_);
  nor _74574_ (_23664_, _13122_, _09531_);
  nor _74575_ (_23665_, _23664_, _23650_);
  nor _74576_ (_23666_, _23665_, _04444_);
  or _74577_ (_23667_, _23666_, _23663_);
  and _74578_ (_23668_, _23667_, _03517_);
  nor _74579_ (_23669_, _05807_, _23648_);
  and _74580_ (_23670_, _13145_, _05807_);
  nor _74581_ (_23671_, _23670_, _23669_);
  nor _74582_ (_23672_, _23671_, _03517_);
  or _74583_ (_23673_, _23672_, _03568_);
  or _74584_ (_23674_, _23673_, _23668_);
  nand _74585_ (_23675_, _23655_, _03568_);
  and _74586_ (_23676_, _23675_, _23674_);
  and _74587_ (_23677_, _23676_, _03583_);
  nor _74588_ (_23678_, _23658_, _03583_);
  or _74589_ (_23679_, _23678_, _23677_);
  and _74590_ (_23680_, _23679_, _03513_);
  and _74591_ (_23682_, _13130_, _05807_);
  nor _74592_ (_23683_, _23682_, _23669_);
  nor _74593_ (_23684_, _23683_, _03513_);
  or _74594_ (_23685_, _23684_, _23680_);
  and _74595_ (_23686_, _23685_, _03506_);
  nor _74596_ (_23687_, _23669_, _13160_);
  nor _74597_ (_23688_, _23687_, _23671_);
  and _74598_ (_23689_, _23688_, _03505_);
  or _74599_ (_23690_, _23689_, _23686_);
  and _74600_ (_23691_, _23690_, _03500_);
  nor _74601_ (_23693_, _13178_, _09570_);
  nor _74602_ (_23694_, _23693_, _23669_);
  nor _74603_ (_23695_, _23694_, _03500_);
  nor _74604_ (_23696_, _23695_, _07314_);
  not _74605_ (_23697_, _23696_);
  nor _74606_ (_23698_, _23697_, _23691_);
  nor _74607_ (_23699_, _23698_, _23656_);
  nor _74608_ (_23700_, _23699_, _03479_);
  and _74609_ (_23701_, _06713_, _05193_);
  nor _74610_ (_23702_, _23650_, _06044_);
  not _74611_ (_23704_, _23702_);
  nor _74612_ (_23705_, _23704_, _23701_);
  or _74613_ (_23706_, _23705_, _03221_);
  nor _74614_ (_23707_, _23706_, _23700_);
  nor _74615_ (_23708_, _13237_, _09531_);
  nor _74616_ (_23709_, _23708_, _23650_);
  nor _74617_ (_23710_, _23709_, _03474_);
  or _74618_ (_23711_, _23710_, _03437_);
  or _74619_ (_23712_, _23711_, _23707_);
  and _74620_ (_23713_, _13244_, _05193_);
  nor _74621_ (_23715_, _23713_, _23650_);
  nand _74622_ (_23716_, _23715_, _03437_);
  and _74623_ (_23717_, _23716_, _23712_);
  nor _74624_ (_23718_, _23717_, _03636_);
  and _74625_ (_23719_, _13253_, _05193_);
  or _74626_ (_23720_, _23650_, _04499_);
  nor _74627_ (_23721_, _23720_, _23719_);
  or _74628_ (_23722_, _23721_, _03769_);
  nor _74629_ (_23723_, _23722_, _23718_);
  nor _74630_ (_23724_, _23723_, _23653_);
  nor _74631_ (_23726_, _23724_, _04504_);
  not _74632_ (_23727_, _23650_);
  and _74633_ (_23728_, _23727_, _05376_);
  or _74634_ (_23729_, _23715_, _04505_);
  nor _74635_ (_23730_, _23729_, _23728_);
  nor _74636_ (_23731_, _23730_, _23726_);
  nor _74637_ (_23732_, _23731_, _03752_);
  or _74638_ (_23733_, _23728_, _03753_);
  or _74639_ (_23734_, _23733_, _23658_);
  and _74640_ (_23735_, _23734_, _03759_);
  not _74641_ (_23736_, _23735_);
  nor _74642_ (_23737_, _23736_, _23732_);
  nor _74643_ (_23738_, _13251_, _09531_);
  or _74644_ (_23739_, _23650_, _03759_);
  nor _74645_ (_23740_, _23739_, _23738_);
  or _74646_ (_23741_, _23740_, _03760_);
  nor _74647_ (_23742_, _23741_, _23737_);
  nor _74648_ (_23743_, _13258_, _09531_);
  nor _74649_ (_23744_, _23743_, _23650_);
  nor _74650_ (_23745_, _23744_, _04517_);
  or _74651_ (_23747_, _23745_, _23742_);
  and _74652_ (_23748_, _23747_, _04192_);
  nor _74653_ (_23749_, _23665_, _04192_);
  or _74654_ (_23750_, _23749_, _23748_);
  and _74655_ (_23751_, _23750_, _03152_);
  nor _74656_ (_23752_, _23683_, _03152_);
  or _74657_ (_23753_, _23752_, _23751_);
  and _74658_ (_23754_, _23753_, _03521_);
  and _74659_ (_23755_, _13312_, _05193_);
  nor _74660_ (_23756_, _23755_, _23650_);
  nor _74661_ (_23758_, _23756_, _03521_);
  or _74662_ (_23759_, _23758_, _23754_);
  or _74663_ (_23760_, _23759_, _42967_);
  or _74664_ (_23761_, _42963_, \oc8051_golden_model_1.IE [6]);
  and _74665_ (_23762_, _23761_, _41755_);
  and _74666_ (_43297_, _23762_, _23760_);
  not _74667_ (_23763_, \oc8051_golden_model_1.IP [0]);
  nor _74668_ (_23764_, _05224_, _23763_);
  and _74669_ (_23765_, _11995_, _05224_);
  nor _74670_ (_23766_, _23765_, _23764_);
  nor _74671_ (_23768_, _23766_, _04501_);
  and _74672_ (_23769_, _05941_, _05224_);
  nor _74673_ (_23770_, _23769_, _23764_);
  nor _74674_ (_23771_, _23770_, _04444_);
  nor _74675_ (_23772_, _04426_, _23763_);
  and _74676_ (_23773_, _05224_, \oc8051_golden_model_1.ACC [0]);
  nor _74677_ (_23774_, _23773_, _23764_);
  nor _74678_ (_23775_, _23774_, _04427_);
  nor _74679_ (_23776_, _23775_, _23772_);
  nor _74680_ (_23777_, _23776_, _03570_);
  or _74681_ (_23779_, _23777_, _03516_);
  nor _74682_ (_23780_, _23779_, _23771_);
  and _74683_ (_23781_, _11887_, _05790_);
  nor _74684_ (_23782_, _05790_, _23763_);
  or _74685_ (_23783_, _23782_, _03517_);
  nor _74686_ (_23784_, _23783_, _23781_);
  or _74687_ (_23785_, _23784_, _03568_);
  nor _74688_ (_23786_, _23785_, _23780_);
  and _74689_ (_23787_, _05224_, _04419_);
  nor _74690_ (_23788_, _23787_, _23764_);
  nor _74691_ (_23790_, _23788_, _03983_);
  or _74692_ (_23791_, _23790_, _23786_);
  and _74693_ (_23792_, _23791_, _03583_);
  nor _74694_ (_23793_, _23774_, _03583_);
  or _74695_ (_23794_, _23793_, _23792_);
  and _74696_ (_23795_, _23794_, _03513_);
  and _74697_ (_23796_, _23764_, _03512_);
  or _74698_ (_23797_, _23796_, _23795_);
  and _74699_ (_23798_, _23797_, _03506_);
  nor _74700_ (_23799_, _23770_, _03506_);
  or _74701_ (_23801_, _23799_, _23798_);
  and _74702_ (_23802_, _23801_, _03500_);
  nor _74703_ (_23803_, _11916_, _09678_);
  nor _74704_ (_23804_, _23803_, _23782_);
  nor _74705_ (_23805_, _23804_, _03500_);
  or _74706_ (_23806_, _23805_, _07314_);
  nor _74707_ (_23807_, _23806_, _23802_);
  and _74708_ (_23808_, _23788_, _07314_);
  or _74709_ (_23809_, _23808_, _03479_);
  nor _74710_ (_23810_, _23809_, _23807_);
  and _74711_ (_23812_, _06715_, _05224_);
  or _74712_ (_23813_, _23812_, _23764_);
  and _74713_ (_23814_, _23813_, _03479_);
  or _74714_ (_23815_, _23814_, _03221_);
  or _74715_ (_23816_, _23815_, _23810_);
  nor _74716_ (_23817_, _11975_, _09641_);
  or _74717_ (_23818_, _23764_, _03474_);
  or _74718_ (_23819_, _23818_, _23817_);
  and _74719_ (_23820_, _23819_, _03438_);
  and _74720_ (_23821_, _23820_, _23816_);
  and _74721_ (_23823_, _05224_, _06202_);
  nor _74722_ (_23824_, _23823_, _23764_);
  nor _74723_ (_23825_, _23824_, _03438_);
  or _74724_ (_23826_, _23825_, _03636_);
  nor _74725_ (_23827_, _23826_, _23821_);
  and _74726_ (_23828_, _11990_, _05224_);
  or _74727_ (_23829_, _23764_, _04499_);
  nor _74728_ (_23830_, _23829_, _23828_);
  or _74729_ (_23831_, _23830_, _03769_);
  nor _74730_ (_23832_, _23831_, _23827_);
  nor _74731_ (_23834_, _23832_, _23768_);
  nor _74732_ (_23835_, _23834_, _04504_);
  or _74733_ (_23836_, _23824_, _04505_);
  nor _74734_ (_23837_, _23836_, _23769_);
  nor _74735_ (_23838_, _23837_, _23835_);
  nor _74736_ (_23839_, _23838_, _03752_);
  and _74737_ (_23840_, _11994_, _05224_);
  or _74738_ (_23841_, _23840_, _23764_);
  and _74739_ (_23842_, _23841_, _03752_);
  or _74740_ (_23843_, _23842_, _23839_);
  and _74741_ (_23845_, _23843_, _03759_);
  nor _74742_ (_23846_, _11988_, _09641_);
  nor _74743_ (_23847_, _23846_, _23764_);
  nor _74744_ (_23848_, _23847_, _03759_);
  or _74745_ (_23849_, _23848_, _23845_);
  and _74746_ (_23850_, _23849_, _04517_);
  nor _74747_ (_23851_, _11870_, _09641_);
  nor _74748_ (_23852_, _23851_, _23764_);
  nor _74749_ (_23853_, _23852_, _04517_);
  or _74750_ (_23854_, _23853_, _23850_);
  and _74751_ (_23856_, _23854_, _04192_);
  nor _74752_ (_23857_, _23770_, _04192_);
  or _74753_ (_23858_, _23857_, _23856_);
  and _74754_ (_23859_, _23858_, _03152_);
  and _74755_ (_23860_, _23764_, _03151_);
  nor _74756_ (_23861_, _23860_, _23859_);
  or _74757_ (_23862_, _23861_, _03520_);
  or _74758_ (_23863_, _23770_, _03521_);
  and _74759_ (_23864_, _23863_, _23862_);
  nand _74760_ (_23865_, _23864_, _42963_);
  or _74761_ (_23867_, _42963_, \oc8051_golden_model_1.IP [0]);
  and _74762_ (_23868_, _23867_, _41755_);
  and _74763_ (_43300_, _23868_, _23865_);
  not _74764_ (_23869_, \oc8051_golden_model_1.IP [1]);
  nor _74765_ (_23870_, _05224_, _23869_);
  and _74766_ (_23871_, _06714_, _05224_);
  or _74767_ (_23872_, _23871_, _23870_);
  and _74768_ (_23873_, _23872_, _03479_);
  nor _74769_ (_23874_, _05224_, \oc8051_golden_model_1.IP [1]);
  and _74770_ (_23875_, _05224_, _03233_);
  nor _74771_ (_23877_, _23875_, _23874_);
  and _74772_ (_23878_, _23877_, _04426_);
  nor _74773_ (_23879_, _04426_, _23869_);
  or _74774_ (_23880_, _23879_, _23878_);
  and _74775_ (_23881_, _23880_, _04444_);
  and _74776_ (_23882_, _12252_, _05224_);
  nor _74777_ (_23883_, _23882_, _23874_);
  and _74778_ (_23884_, _23883_, _03570_);
  or _74779_ (_23885_, _23884_, _23881_);
  and _74780_ (_23886_, _23885_, _03517_);
  and _74781_ (_23888_, _12083_, _05790_);
  nor _74782_ (_23889_, _05790_, _23869_);
  or _74783_ (_23890_, _23889_, _03568_);
  or _74784_ (_23891_, _23890_, _23888_);
  and _74785_ (_23892_, _23891_, _14165_);
  nor _74786_ (_23893_, _23892_, _23886_);
  nor _74787_ (_23894_, _09641_, _04603_);
  nor _74788_ (_23895_, _23894_, _23870_);
  and _74789_ (_23896_, _23895_, _03568_);
  nor _74790_ (_23897_, _23896_, _23893_);
  and _74791_ (_23899_, _23897_, _03583_);
  and _74792_ (_23900_, _23877_, _03575_);
  or _74793_ (_23901_, _23900_, _23899_);
  and _74794_ (_23902_, _23901_, _03513_);
  and _74795_ (_23903_, _12069_, _05790_);
  nor _74796_ (_23904_, _23903_, _23889_);
  nor _74797_ (_23905_, _23904_, _03513_);
  or _74798_ (_23906_, _23905_, _23902_);
  and _74799_ (_23907_, _23906_, _03506_);
  and _74800_ (_23908_, _23888_, _12098_);
  or _74801_ (_23910_, _23908_, _23889_);
  and _74802_ (_23911_, _23910_, _03505_);
  or _74803_ (_23912_, _23911_, _23907_);
  and _74804_ (_23913_, _23912_, _03500_);
  nor _74805_ (_23914_, _12116_, _09678_);
  nor _74806_ (_23915_, _23889_, _23914_);
  nor _74807_ (_23916_, _23915_, _03500_);
  or _74808_ (_23917_, _23916_, _07314_);
  nor _74809_ (_23918_, _23917_, _23913_);
  and _74810_ (_23919_, _23895_, _07314_);
  or _74811_ (_23921_, _23919_, _03479_);
  nor _74812_ (_23922_, _23921_, _23918_);
  or _74813_ (_23923_, _23922_, _23873_);
  and _74814_ (_23924_, _23923_, _03474_);
  nor _74815_ (_23925_, _12176_, _09641_);
  nor _74816_ (_23926_, _23925_, _23870_);
  nor _74817_ (_23927_, _23926_, _03474_);
  nor _74818_ (_23928_, _23927_, _23924_);
  nor _74819_ (_23929_, _23928_, _03437_);
  and _74820_ (_23930_, _05224_, _04317_);
  not _74821_ (_23932_, _23930_);
  nor _74822_ (_23933_, _23874_, _03438_);
  and _74823_ (_23934_, _23933_, _23932_);
  nor _74824_ (_23935_, _23934_, _23929_);
  nor _74825_ (_23936_, _23935_, _03636_);
  not _74826_ (_23937_, _23874_);
  nor _74827_ (_23938_, _12191_, _09641_);
  nor _74828_ (_23939_, _23938_, _04499_);
  and _74829_ (_23940_, _23939_, _23937_);
  nor _74830_ (_23941_, _23940_, _23936_);
  nor _74831_ (_23943_, _23941_, _03769_);
  nor _74832_ (_23944_, _12197_, _09641_);
  nor _74833_ (_23945_, _23944_, _04501_);
  and _74834_ (_23946_, _23945_, _23937_);
  nor _74835_ (_23947_, _23946_, _23943_);
  nor _74836_ (_23948_, _23947_, _04504_);
  nor _74837_ (_23949_, _12190_, _09641_);
  nor _74838_ (_23950_, _23949_, _05769_);
  and _74839_ (_23951_, _23950_, _23937_);
  nor _74840_ (_23952_, _23951_, _23948_);
  nor _74841_ (_23954_, _23952_, _03752_);
  nor _74842_ (_23955_, _23870_, _05569_);
  nor _74843_ (_23956_, _23955_, _03753_);
  and _74844_ (_23957_, _23956_, _23877_);
  nor _74845_ (_23958_, _23957_, _23954_);
  nor _74846_ (_23959_, _23958_, _03758_);
  and _74847_ (_23960_, _23930_, _05940_);
  nor _74848_ (_23961_, _23960_, _03759_);
  and _74849_ (_23962_, _23961_, _23937_);
  nor _74850_ (_23963_, _23962_, _23959_);
  nor _74851_ (_23965_, _23963_, _03760_);
  nand _74852_ (_23966_, _23875_, _05940_);
  nor _74853_ (_23967_, _23874_, _04517_);
  and _74854_ (_23968_, _23967_, _23966_);
  or _74855_ (_23969_, _23968_, _03790_);
  nor _74856_ (_23970_, _23969_, _23965_);
  nor _74857_ (_23971_, _23883_, _04192_);
  or _74858_ (_23972_, _23971_, _03151_);
  nor _74859_ (_23973_, _23972_, _23970_);
  nor _74860_ (_23974_, _23904_, _03152_);
  or _74861_ (_23976_, _23974_, _03520_);
  nor _74862_ (_23977_, _23976_, _23973_);
  or _74863_ (_23978_, _23870_, _03521_);
  nor _74864_ (_23979_, _23978_, _23882_);
  nor _74865_ (_23980_, _23979_, _23977_);
  or _74866_ (_23981_, _23980_, _42967_);
  or _74867_ (_23982_, _42963_, \oc8051_golden_model_1.IP [1]);
  and _74868_ (_23983_, _23982_, _41755_);
  and _74869_ (_43301_, _23983_, _23981_);
  not _74870_ (_23984_, \oc8051_golden_model_1.IP [2]);
  nor _74871_ (_23986_, _05224_, _23984_);
  and _74872_ (_23987_, _12401_, _05224_);
  nor _74873_ (_23988_, _23987_, _23986_);
  nor _74874_ (_23989_, _23988_, _04501_);
  nor _74875_ (_23990_, _09641_, _05026_);
  nor _74876_ (_23991_, _23990_, _23986_);
  and _74877_ (_23992_, _23991_, _07314_);
  and _74878_ (_23993_, _05224_, \oc8051_golden_model_1.ACC [2]);
  nor _74879_ (_23994_, _23993_, _23986_);
  nor _74880_ (_23995_, _23994_, _04427_);
  nor _74881_ (_23997_, _04426_, _23984_);
  or _74882_ (_23998_, _23997_, _23995_);
  and _74883_ (_23999_, _23998_, _04444_);
  nor _74884_ (_24000_, _12282_, _09641_);
  nor _74885_ (_24001_, _24000_, _23986_);
  nor _74886_ (_24002_, _24001_, _04444_);
  or _74887_ (_24003_, _24002_, _23999_);
  and _74888_ (_24004_, _24003_, _03517_);
  nor _74889_ (_24005_, _05790_, _23984_);
  and _74890_ (_24006_, _12278_, _05790_);
  nor _74891_ (_24008_, _24006_, _24005_);
  nor _74892_ (_24009_, _24008_, _03517_);
  or _74893_ (_24010_, _24009_, _24004_);
  and _74894_ (_24011_, _24010_, _03983_);
  nor _74895_ (_24012_, _23991_, _03983_);
  or _74896_ (_24013_, _24012_, _24011_);
  and _74897_ (_24014_, _24013_, _03583_);
  nor _74898_ (_24015_, _23994_, _03583_);
  or _74899_ (_24016_, _24015_, _24014_);
  and _74900_ (_24017_, _24016_, _03513_);
  and _74901_ (_24019_, _12276_, _05790_);
  nor _74902_ (_24020_, _24019_, _24005_);
  nor _74903_ (_24021_, _24020_, _03513_);
  or _74904_ (_24022_, _24021_, _03505_);
  or _74905_ (_24023_, _24022_, _24017_);
  and _74906_ (_24024_, _24006_, _12309_);
  or _74907_ (_24025_, _24005_, _03506_);
  or _74908_ (_24026_, _24025_, _24024_);
  and _74909_ (_24027_, _24026_, _03500_);
  and _74910_ (_24028_, _24027_, _24023_);
  nor _74911_ (_24030_, _12326_, _09678_);
  nor _74912_ (_24031_, _24030_, _24005_);
  nor _74913_ (_24032_, _24031_, _03500_);
  nor _74914_ (_24033_, _24032_, _07314_);
  not _74915_ (_24034_, _24033_);
  nor _74916_ (_24035_, _24034_, _24028_);
  nor _74917_ (_24036_, _24035_, _23992_);
  nor _74918_ (_24037_, _24036_, _03479_);
  and _74919_ (_24038_, _06718_, _05224_);
  nor _74920_ (_24039_, _23986_, _06044_);
  not _74921_ (_24041_, _24039_);
  nor _74922_ (_24042_, _24041_, _24038_);
  or _74923_ (_24043_, _24042_, _03221_);
  nor _74924_ (_24044_, _24043_, _24037_);
  nor _74925_ (_24045_, _12384_, _09641_);
  nor _74926_ (_24046_, _24045_, _23986_);
  nor _74927_ (_24047_, _24046_, _03474_);
  or _74928_ (_24048_, _24047_, _03437_);
  or _74929_ (_24049_, _24048_, _24044_);
  and _74930_ (_24050_, _05224_, _06261_);
  nor _74931_ (_24052_, _24050_, _23986_);
  nand _74932_ (_24053_, _24052_, _03437_);
  and _74933_ (_24054_, _24053_, _24049_);
  nor _74934_ (_24055_, _24054_, _03636_);
  and _74935_ (_24056_, _12273_, _05224_);
  or _74936_ (_24057_, _23986_, _04499_);
  nor _74937_ (_24058_, _24057_, _24056_);
  or _74938_ (_24059_, _24058_, _03769_);
  nor _74939_ (_24060_, _24059_, _24055_);
  nor _74940_ (_24061_, _24060_, _23989_);
  nor _74941_ (_24063_, _24061_, _04504_);
  not _74942_ (_24064_, _23986_);
  and _74943_ (_24065_, _24064_, _05664_);
  or _74944_ (_24066_, _24052_, _04505_);
  nor _74945_ (_24067_, _24066_, _24065_);
  nor _74946_ (_24068_, _24067_, _24063_);
  nor _74947_ (_24069_, _24068_, _03752_);
  or _74948_ (_24070_, _24065_, _03753_);
  or _74949_ (_24071_, _24070_, _23994_);
  and _74950_ (_24072_, _24071_, _03759_);
  not _74951_ (_24074_, _24072_);
  nor _74952_ (_24075_, _24074_, _24069_);
  nor _74953_ (_24076_, _12272_, _09641_);
  or _74954_ (_24077_, _23986_, _03759_);
  nor _74955_ (_24078_, _24077_, _24076_);
  or _74956_ (_24079_, _24078_, _03760_);
  nor _74957_ (_24080_, _24079_, _24075_);
  nor _74958_ (_24081_, _12400_, _09641_);
  nor _74959_ (_24082_, _24081_, _23986_);
  nor _74960_ (_24083_, _24082_, _04517_);
  or _74961_ (_24085_, _24083_, _24080_);
  and _74962_ (_24086_, _24085_, _04192_);
  nor _74963_ (_24087_, _24001_, _04192_);
  or _74964_ (_24088_, _24087_, _24086_);
  and _74965_ (_24089_, _24088_, _03152_);
  nor _74966_ (_24090_, _24020_, _03152_);
  or _74967_ (_24091_, _24090_, _24089_);
  and _74968_ (_24092_, _24091_, _03521_);
  and _74969_ (_24093_, _12456_, _05224_);
  nor _74970_ (_24094_, _24093_, _23986_);
  nor _74971_ (_24096_, _24094_, _03521_);
  or _74972_ (_24097_, _24096_, _24092_);
  or _74973_ (_24098_, _24097_, _42967_);
  or _74974_ (_24099_, _42963_, \oc8051_golden_model_1.IP [2]);
  and _74975_ (_24100_, _24099_, _41755_);
  and _74976_ (_43302_, _24100_, _24098_);
  not _74977_ (_24101_, \oc8051_golden_model_1.IP [3]);
  nor _74978_ (_24102_, _05224_, _24101_);
  and _74979_ (_24103_, _12604_, _05224_);
  nor _74980_ (_24104_, _24103_, _24102_);
  nor _74981_ (_24106_, _24104_, _04501_);
  nor _74982_ (_24107_, _09641_, _04843_);
  nor _74983_ (_24108_, _24107_, _24102_);
  and _74984_ (_24109_, _24108_, _07314_);
  and _74985_ (_24110_, _05224_, \oc8051_golden_model_1.ACC [3]);
  nor _74986_ (_24111_, _24110_, _24102_);
  nor _74987_ (_24112_, _24111_, _04427_);
  nor _74988_ (_24113_, _04426_, _24101_);
  or _74989_ (_24114_, _24113_, _24112_);
  and _74990_ (_24115_, _24114_, _04444_);
  nor _74991_ (_24117_, _12486_, _09641_);
  nor _74992_ (_24118_, _24117_, _24102_);
  nor _74993_ (_24119_, _24118_, _04444_);
  or _74994_ (_24120_, _24119_, _24115_);
  and _74995_ (_24121_, _24120_, _03517_);
  nor _74996_ (_24122_, _05790_, _24101_);
  and _74997_ (_24123_, _12490_, _05790_);
  nor _74998_ (_24124_, _24123_, _24122_);
  nor _74999_ (_24125_, _24124_, _03517_);
  or _75000_ (_24126_, _24125_, _03568_);
  or _75001_ (_24128_, _24126_, _24121_);
  nand _75002_ (_24129_, _24108_, _03568_);
  and _75003_ (_24130_, _24129_, _24128_);
  and _75004_ (_24131_, _24130_, _03583_);
  nor _75005_ (_24132_, _24111_, _03583_);
  or _75006_ (_24133_, _24132_, _24131_);
  and _75007_ (_24134_, _24133_, _03513_);
  and _75008_ (_24135_, _12500_, _05790_);
  nor _75009_ (_24136_, _24135_, _24122_);
  nor _75010_ (_24137_, _24136_, _03513_);
  or _75011_ (_24139_, _24137_, _24134_);
  and _75012_ (_24140_, _24139_, _03506_);
  nor _75013_ (_24141_, _24122_, _12507_);
  nor _75014_ (_24142_, _24141_, _24124_);
  and _75015_ (_24143_, _24142_, _03505_);
  or _75016_ (_24144_, _24143_, _24140_);
  and _75017_ (_24145_, _24144_, _03500_);
  nor _75018_ (_24146_, _12525_, _09678_);
  nor _75019_ (_24147_, _24146_, _24122_);
  nor _75020_ (_24148_, _24147_, _03500_);
  nor _75021_ (_24150_, _24148_, _07314_);
  not _75022_ (_24151_, _24150_);
  nor _75023_ (_24152_, _24151_, _24145_);
  nor _75024_ (_24153_, _24152_, _24109_);
  nor _75025_ (_24154_, _24153_, _03479_);
  and _75026_ (_24155_, _06717_, _05224_);
  nor _75027_ (_24156_, _24102_, _06044_);
  not _75028_ (_24157_, _24156_);
  nor _75029_ (_24158_, _24157_, _24155_);
  or _75030_ (_24159_, _24158_, _03221_);
  nor _75031_ (_24161_, _24159_, _24154_);
  nor _75032_ (_24162_, _12583_, _09641_);
  nor _75033_ (_24163_, _24162_, _24102_);
  nor _75034_ (_24164_, _24163_, _03474_);
  or _75035_ (_24165_, _24164_, _03437_);
  or _75036_ (_24166_, _24165_, _24161_);
  and _75037_ (_24167_, _05224_, _06217_);
  nor _75038_ (_24168_, _24167_, _24102_);
  nand _75039_ (_24169_, _24168_, _03437_);
  and _75040_ (_24170_, _24169_, _24166_);
  nor _75041_ (_24172_, _24170_, _03636_);
  and _75042_ (_24173_, _12598_, _05224_);
  or _75043_ (_24174_, _24102_, _04499_);
  nor _75044_ (_24175_, _24174_, _24173_);
  or _75045_ (_24176_, _24175_, _03769_);
  nor _75046_ (_24177_, _24176_, _24172_);
  nor _75047_ (_24178_, _24177_, _24106_);
  nor _75048_ (_24179_, _24178_, _04504_);
  not _75049_ (_24180_, _24102_);
  and _75050_ (_24181_, _24180_, _05520_);
  or _75051_ (_24184_, _24168_, _04505_);
  nor _75052_ (_24185_, _24184_, _24181_);
  nor _75053_ (_24186_, _24185_, _24179_);
  nor _75054_ (_24187_, _24186_, _03752_);
  or _75055_ (_24188_, _24181_, _03753_);
  or _75056_ (_24189_, _24188_, _24111_);
  and _75057_ (_24190_, _24189_, _03759_);
  not _75058_ (_24191_, _24190_);
  nor _75059_ (_24192_, _24191_, _24187_);
  nor _75060_ (_24193_, _12597_, _09641_);
  or _75061_ (_24196_, _24102_, _03759_);
  nor _75062_ (_24197_, _24196_, _24193_);
  or _75063_ (_24198_, _24197_, _03760_);
  nor _75064_ (_24199_, _24198_, _24192_);
  nor _75065_ (_24200_, _12603_, _09641_);
  nor _75066_ (_24201_, _24200_, _24102_);
  nor _75067_ (_24202_, _24201_, _04517_);
  or _75068_ (_24203_, _24202_, _24199_);
  and _75069_ (_24204_, _24203_, _04192_);
  nor _75070_ (_24205_, _24118_, _04192_);
  or _75071_ (_24208_, _24205_, _24204_);
  and _75072_ (_24209_, _24208_, _03152_);
  nor _75073_ (_24210_, _24136_, _03152_);
  or _75074_ (_24211_, _24210_, _24209_);
  and _75075_ (_24212_, _24211_, _03521_);
  and _75076_ (_24213_, _12658_, _05224_);
  nor _75077_ (_24214_, _24213_, _24102_);
  nor _75078_ (_24215_, _24214_, _03521_);
  or _75079_ (_24216_, _24215_, _24212_);
  or _75080_ (_24217_, _24216_, _42967_);
  or _75081_ (_24220_, _42963_, \oc8051_golden_model_1.IP [3]);
  and _75082_ (_24221_, _24220_, _41755_);
  and _75083_ (_43303_, _24221_, _24217_);
  not _75084_ (_24222_, \oc8051_golden_model_1.IP [4]);
  nor _75085_ (_24223_, _05224_, _24222_);
  and _75086_ (_24224_, _12844_, _05224_);
  nor _75087_ (_24225_, _24224_, _24223_);
  nor _75088_ (_24226_, _24225_, _04501_);
  nor _75089_ (_24227_, _05712_, _09641_);
  nor _75090_ (_24228_, _24227_, _24223_);
  and _75091_ (_24231_, _24228_, _07314_);
  and _75092_ (_24232_, _05224_, \oc8051_golden_model_1.ACC [4]);
  nor _75093_ (_24233_, _24232_, _24223_);
  nor _75094_ (_24234_, _24233_, _04427_);
  nor _75095_ (_24235_, _04426_, _24222_);
  or _75096_ (_24236_, _24235_, _24234_);
  and _75097_ (_24237_, _24236_, _04444_);
  nor _75098_ (_24238_, _12733_, _09641_);
  nor _75099_ (_24239_, _24238_, _24223_);
  nor _75100_ (_24240_, _24239_, _04444_);
  or _75101_ (_24243_, _24240_, _24237_);
  and _75102_ (_24244_, _24243_, _03517_);
  nor _75103_ (_24245_, _05790_, _24222_);
  and _75104_ (_24246_, _12737_, _05790_);
  nor _75105_ (_24247_, _24246_, _24245_);
  nor _75106_ (_24248_, _24247_, _03517_);
  or _75107_ (_24249_, _24248_, _03568_);
  or _75108_ (_24250_, _24249_, _24244_);
  nand _75109_ (_24251_, _24228_, _03568_);
  and _75110_ (_24252_, _24251_, _24250_);
  and _75111_ (_24255_, _24252_, _03583_);
  nor _75112_ (_24256_, _24233_, _03583_);
  or _75113_ (_24257_, _24256_, _24255_);
  and _75114_ (_24258_, _24257_, _03513_);
  and _75115_ (_24259_, _12718_, _05790_);
  nor _75116_ (_24260_, _24259_, _24245_);
  nor _75117_ (_24261_, _24260_, _03513_);
  or _75118_ (_24262_, _24261_, _24258_);
  and _75119_ (_24263_, _24262_, _03506_);
  nor _75120_ (_24264_, _24245_, _12752_);
  nor _75121_ (_24266_, _24264_, _24247_);
  and _75122_ (_24267_, _24266_, _03505_);
  or _75123_ (_24268_, _24267_, _24263_);
  and _75124_ (_24269_, _24268_, _03500_);
  nor _75125_ (_24270_, _12716_, _09678_);
  nor _75126_ (_24271_, _24270_, _24245_);
  nor _75127_ (_24272_, _24271_, _03500_);
  nor _75128_ (_24273_, _24272_, _07314_);
  not _75129_ (_24274_, _24273_);
  nor _75130_ (_24275_, _24274_, _24269_);
  nor _75131_ (_24277_, _24275_, _24231_);
  nor _75132_ (_24278_, _24277_, _03479_);
  and _75133_ (_24279_, _06722_, _05224_);
  nor _75134_ (_24280_, _24223_, _06044_);
  not _75135_ (_24281_, _24280_);
  nor _75136_ (_24282_, _24281_, _24279_);
  or _75137_ (_24283_, _24282_, _03221_);
  nor _75138_ (_24284_, _24283_, _24278_);
  nor _75139_ (_24285_, _12827_, _09641_);
  nor _75140_ (_24286_, _24285_, _24223_);
  nor _75141_ (_24288_, _24286_, _03474_);
  or _75142_ (_24289_, _24288_, _03437_);
  or _75143_ (_24290_, _24289_, _24284_);
  and _75144_ (_24291_, _06233_, _05224_);
  nor _75145_ (_24292_, _24291_, _24223_);
  nand _75146_ (_24293_, _24292_, _03437_);
  and _75147_ (_24294_, _24293_, _24290_);
  nor _75148_ (_24295_, _24294_, _03636_);
  and _75149_ (_24296_, _12711_, _05224_);
  or _75150_ (_24297_, _24223_, _04499_);
  nor _75151_ (_24299_, _24297_, _24296_);
  or _75152_ (_24300_, _24299_, _03769_);
  nor _75153_ (_24301_, _24300_, _24295_);
  nor _75154_ (_24302_, _24301_, _24226_);
  nor _75155_ (_24303_, _24302_, _04504_);
  not _75156_ (_24304_, _24223_);
  and _75157_ (_24305_, _24304_, _05760_);
  or _75158_ (_24306_, _24292_, _04505_);
  nor _75159_ (_24307_, _24306_, _24305_);
  nor _75160_ (_24308_, _24307_, _24303_);
  nor _75161_ (_24310_, _24308_, _03752_);
  or _75162_ (_24311_, _24305_, _03753_);
  nor _75163_ (_24312_, _24311_, _24233_);
  or _75164_ (_24313_, _24312_, _24310_);
  and _75165_ (_24314_, _24313_, _03759_);
  nor _75166_ (_24315_, _12710_, _09641_);
  nor _75167_ (_24316_, _24315_, _24223_);
  nor _75168_ (_24317_, _24316_, _03759_);
  or _75169_ (_24318_, _24317_, _24314_);
  and _75170_ (_24319_, _24318_, _04517_);
  nor _75171_ (_24321_, _12843_, _09641_);
  nor _75172_ (_24322_, _24321_, _24223_);
  nor _75173_ (_24323_, _24322_, _04517_);
  or _75174_ (_24324_, _24323_, _24319_);
  and _75175_ (_24325_, _24324_, _04192_);
  nor _75176_ (_24326_, _24239_, _04192_);
  or _75177_ (_24327_, _24326_, _24325_);
  and _75178_ (_24328_, _24327_, _03152_);
  nor _75179_ (_24329_, _24260_, _03152_);
  or _75180_ (_24330_, _24329_, _24328_);
  and _75181_ (_24332_, _24330_, _03521_);
  and _75182_ (_24333_, _12893_, _05224_);
  nor _75183_ (_24334_, _24333_, _24223_);
  nor _75184_ (_24335_, _24334_, _03521_);
  or _75185_ (_24336_, _24335_, _24332_);
  or _75186_ (_24337_, _24336_, _42967_);
  or _75187_ (_24338_, _42963_, \oc8051_golden_model_1.IP [4]);
  and _75188_ (_24339_, _24338_, _41755_);
  and _75189_ (_43304_, _24339_, _24337_);
  not _75190_ (_24340_, \oc8051_golden_model_1.IP [5]);
  nor _75191_ (_24342_, _05224_, _24340_);
  and _75192_ (_24343_, _13042_, _05224_);
  nor _75193_ (_24344_, _24343_, _24342_);
  nor _75194_ (_24345_, _24344_, _04501_);
  nor _75195_ (_24346_, _05422_, _09641_);
  nor _75196_ (_24347_, _24346_, _24342_);
  and _75197_ (_24348_, _24347_, _07314_);
  and _75198_ (_24349_, _05224_, \oc8051_golden_model_1.ACC [5]);
  nor _75199_ (_24350_, _24349_, _24342_);
  nor _75200_ (_24351_, _24350_, _04427_);
  nor _75201_ (_24353_, _04426_, _24340_);
  or _75202_ (_24354_, _24353_, _24351_);
  and _75203_ (_24355_, _24354_, _04444_);
  nor _75204_ (_24356_, _12930_, _09641_);
  nor _75205_ (_24357_, _24356_, _24342_);
  nor _75206_ (_24358_, _24357_, _04444_);
  or _75207_ (_24359_, _24358_, _24355_);
  and _75208_ (_24360_, _24359_, _03517_);
  nor _75209_ (_24361_, _05790_, _24340_);
  and _75210_ (_24362_, _12934_, _05790_);
  nor _75211_ (_24364_, _24362_, _24361_);
  nor _75212_ (_24365_, _24364_, _03517_);
  or _75213_ (_24366_, _24365_, _03568_);
  or _75214_ (_24367_, _24366_, _24360_);
  nand _75215_ (_24368_, _24347_, _03568_);
  and _75216_ (_24369_, _24368_, _24367_);
  and _75217_ (_24370_, _24369_, _03583_);
  nor _75218_ (_24371_, _24350_, _03583_);
  or _75219_ (_24372_, _24371_, _24370_);
  and _75220_ (_24373_, _24372_, _03513_);
  and _75221_ (_24375_, _12914_, _05790_);
  nor _75222_ (_24376_, _24375_, _24361_);
  nor _75223_ (_24377_, _24376_, _03513_);
  or _75224_ (_24378_, _24377_, _24373_);
  and _75225_ (_24379_, _24378_, _03506_);
  nor _75226_ (_24380_, _24361_, _12949_);
  nor _75227_ (_24381_, _24380_, _24364_);
  and _75228_ (_24382_, _24381_, _03505_);
  or _75229_ (_24383_, _24382_, _24379_);
  and _75230_ (_24384_, _24383_, _03500_);
  nor _75231_ (_24386_, _12912_, _09678_);
  nor _75232_ (_24387_, _24386_, _24361_);
  nor _75233_ (_24388_, _24387_, _03500_);
  nor _75234_ (_24389_, _24388_, _07314_);
  not _75235_ (_24390_, _24389_);
  nor _75236_ (_24391_, _24390_, _24384_);
  nor _75237_ (_24392_, _24391_, _24348_);
  nor _75238_ (_24393_, _24392_, _03479_);
  and _75239_ (_24394_, _06721_, _05224_);
  nor _75240_ (_24395_, _24342_, _06044_);
  not _75241_ (_24397_, _24395_);
  nor _75242_ (_24398_, _24397_, _24394_);
  or _75243_ (_24399_, _24398_, _03221_);
  nor _75244_ (_24400_, _24399_, _24393_);
  nor _75245_ (_24401_, _13021_, _09641_);
  nor _75246_ (_24402_, _24401_, _24342_);
  nor _75247_ (_24403_, _24402_, _03474_);
  or _75248_ (_24404_, _24403_, _03437_);
  or _75249_ (_24405_, _24404_, _24400_);
  and _75250_ (_24406_, _06211_, _05224_);
  nor _75251_ (_24408_, _24406_, _24342_);
  nand _75252_ (_24409_, _24408_, _03437_);
  and _75253_ (_24410_, _24409_, _24405_);
  nor _75254_ (_24411_, _24410_, _03636_);
  and _75255_ (_24412_, _13036_, _05224_);
  or _75256_ (_24413_, _24342_, _04499_);
  nor _75257_ (_24414_, _24413_, _24412_);
  or _75258_ (_24415_, _24414_, _03769_);
  nor _75259_ (_24416_, _24415_, _24411_);
  nor _75260_ (_24417_, _24416_, _24345_);
  nor _75261_ (_24419_, _24417_, _04504_);
  not _75262_ (_24420_, _24342_);
  and _75263_ (_24421_, _24420_, _05471_);
  or _75264_ (_24422_, _24408_, _04505_);
  nor _75265_ (_24423_, _24422_, _24421_);
  nor _75266_ (_24424_, _24423_, _24419_);
  nor _75267_ (_24425_, _24424_, _03752_);
  or _75268_ (_24426_, _24421_, _03753_);
  nor _75269_ (_24427_, _24426_, _24350_);
  or _75270_ (_24428_, _24427_, _24425_);
  and _75271_ (_24430_, _24428_, _03759_);
  nor _75272_ (_24431_, _13035_, _09641_);
  nor _75273_ (_24432_, _24431_, _24342_);
  nor _75274_ (_24433_, _24432_, _03759_);
  or _75275_ (_24434_, _24433_, _24430_);
  and _75276_ (_24435_, _24434_, _04517_);
  nor _75277_ (_24436_, _13041_, _09641_);
  nor _75278_ (_24437_, _24436_, _24342_);
  nor _75279_ (_24438_, _24437_, _04517_);
  or _75280_ (_24439_, _24438_, _24435_);
  and _75281_ (_24441_, _24439_, _04192_);
  nor _75282_ (_24442_, _24357_, _04192_);
  or _75283_ (_24443_, _24442_, _24441_);
  and _75284_ (_24444_, _24443_, _03152_);
  nor _75285_ (_24445_, _24376_, _03152_);
  or _75286_ (_24446_, _24445_, _24444_);
  and _75287_ (_24447_, _24446_, _03521_);
  and _75288_ (_24448_, _13097_, _05224_);
  nor _75289_ (_24449_, _24448_, _24342_);
  nor _75290_ (_24450_, _24449_, _03521_);
  or _75291_ (_24452_, _24450_, _24447_);
  or _75292_ (_24453_, _24452_, _42967_);
  or _75293_ (_24454_, _42963_, \oc8051_golden_model_1.IP [5]);
  and _75294_ (_24455_, _24454_, _41755_);
  and _75295_ (_43305_, _24455_, _24453_);
  not _75296_ (_24456_, \oc8051_golden_model_1.IP [6]);
  nor _75297_ (_24457_, _05224_, _24456_);
  and _75298_ (_24458_, _13259_, _05224_);
  nor _75299_ (_24459_, _24458_, _24457_);
  nor _75300_ (_24460_, _24459_, _04501_);
  nor _75301_ (_24462_, _05327_, _09641_);
  nor _75302_ (_24463_, _24462_, _24457_);
  and _75303_ (_24464_, _24463_, _07314_);
  and _75304_ (_24465_, _05224_, \oc8051_golden_model_1.ACC [6]);
  nor _75305_ (_24466_, _24465_, _24457_);
  nor _75306_ (_24467_, _24466_, _04427_);
  nor _75307_ (_24468_, _04426_, _24456_);
  or _75308_ (_24469_, _24468_, _24467_);
  and _75309_ (_24470_, _24469_, _04444_);
  nor _75310_ (_24471_, _13122_, _09641_);
  nor _75311_ (_24473_, _24471_, _24457_);
  nor _75312_ (_24474_, _24473_, _04444_);
  or _75313_ (_24475_, _24474_, _24470_);
  and _75314_ (_24476_, _24475_, _03517_);
  nor _75315_ (_24477_, _05790_, _24456_);
  and _75316_ (_24478_, _13145_, _05790_);
  nor _75317_ (_24479_, _24478_, _24477_);
  nor _75318_ (_24480_, _24479_, _03517_);
  or _75319_ (_24481_, _24480_, _03568_);
  or _75320_ (_24482_, _24481_, _24476_);
  nand _75321_ (_24484_, _24463_, _03568_);
  and _75322_ (_24485_, _24484_, _24482_);
  and _75323_ (_24486_, _24485_, _03583_);
  nor _75324_ (_24487_, _24466_, _03583_);
  or _75325_ (_24488_, _24487_, _24486_);
  and _75326_ (_24489_, _24488_, _03513_);
  and _75327_ (_24490_, _13130_, _05790_);
  nor _75328_ (_24491_, _24490_, _24477_);
  nor _75329_ (_24492_, _24491_, _03513_);
  or _75330_ (_24493_, _24492_, _03505_);
  or _75331_ (_24495_, _24493_, _24489_);
  nor _75332_ (_24496_, _24477_, _13160_);
  nor _75333_ (_24497_, _24496_, _24479_);
  or _75334_ (_24498_, _24497_, _03506_);
  and _75335_ (_24499_, _24498_, _03500_);
  and _75336_ (_24500_, _24499_, _24495_);
  nor _75337_ (_24501_, _13178_, _09678_);
  nor _75338_ (_24502_, _24501_, _24477_);
  nor _75339_ (_24503_, _24502_, _03500_);
  nor _75340_ (_24504_, _24503_, _07314_);
  not _75341_ (_24506_, _24504_);
  nor _75342_ (_24507_, _24506_, _24500_);
  nor _75343_ (_24508_, _24507_, _24464_);
  nor _75344_ (_24509_, _24508_, _03479_);
  and _75345_ (_24510_, _06713_, _05224_);
  nor _75346_ (_24511_, _24457_, _06044_);
  not _75347_ (_24512_, _24511_);
  nor _75348_ (_24513_, _24512_, _24510_);
  or _75349_ (_24514_, _24513_, _03221_);
  nor _75350_ (_24515_, _24514_, _24509_);
  nor _75351_ (_24517_, _13237_, _09641_);
  nor _75352_ (_24518_, _24517_, _24457_);
  nor _75353_ (_24519_, _24518_, _03474_);
  or _75354_ (_24520_, _24519_, _03437_);
  or _75355_ (_24521_, _24520_, _24515_);
  and _75356_ (_24522_, _13244_, _05224_);
  nor _75357_ (_24523_, _24522_, _24457_);
  nand _75358_ (_24524_, _24523_, _03437_);
  and _75359_ (_24525_, _24524_, _24521_);
  nor _75360_ (_24526_, _24525_, _03636_);
  and _75361_ (_24528_, _13253_, _05224_);
  or _75362_ (_24529_, _24457_, _04499_);
  nor _75363_ (_24530_, _24529_, _24528_);
  or _75364_ (_24531_, _24530_, _03769_);
  nor _75365_ (_24532_, _24531_, _24526_);
  nor _75366_ (_24533_, _24532_, _24460_);
  nor _75367_ (_24534_, _24533_, _04504_);
  not _75368_ (_24535_, _24457_);
  and _75369_ (_24536_, _24535_, _05376_);
  or _75370_ (_24537_, _24523_, _04505_);
  nor _75371_ (_24539_, _24537_, _24536_);
  nor _75372_ (_24540_, _24539_, _24534_);
  nor _75373_ (_24541_, _24540_, _03752_);
  or _75374_ (_24542_, _24536_, _03753_);
  nor _75375_ (_24543_, _24542_, _24466_);
  or _75376_ (_24544_, _24543_, _24541_);
  and _75377_ (_24545_, _24544_, _03759_);
  nor _75378_ (_24546_, _13251_, _09641_);
  nor _75379_ (_24547_, _24546_, _24457_);
  nor _75380_ (_24548_, _24547_, _03759_);
  or _75381_ (_24550_, _24548_, _24545_);
  and _75382_ (_24551_, _24550_, _04517_);
  nor _75383_ (_24552_, _13258_, _09641_);
  nor _75384_ (_24553_, _24552_, _24457_);
  nor _75385_ (_24554_, _24553_, _04517_);
  or _75386_ (_24555_, _24554_, _24551_);
  and _75387_ (_24556_, _24555_, _04192_);
  nor _75388_ (_24557_, _24473_, _04192_);
  or _75389_ (_24558_, _24557_, _24556_);
  and _75390_ (_24559_, _24558_, _03152_);
  nor _75391_ (_24561_, _24491_, _03152_);
  or _75392_ (_24562_, _24561_, _24559_);
  and _75393_ (_24563_, _24562_, _03521_);
  and _75394_ (_24564_, _13312_, _05224_);
  nor _75395_ (_24565_, _24564_, _24457_);
  nor _75396_ (_24566_, _24565_, _03521_);
  or _75397_ (_24567_, _24566_, _24563_);
  or _75398_ (_24568_, _24567_, _42967_);
  or _75399_ (_24569_, _42963_, \oc8051_golden_model_1.IP [6]);
  and _75400_ (_24570_, _24569_, _41755_);
  and _75401_ (_43306_, _24570_, _24568_);
  not _75402_ (_24572_, \oc8051_golden_model_1.DPL [0]);
  nor _75403_ (_24573_, _42963_, _24572_);
  nor _75404_ (_24574_, _05272_, _24572_);
  and _75405_ (_24575_, _05272_, _04419_);
  or _75406_ (_24576_, _24575_, _24574_);
  or _75407_ (_24577_, _24576_, _06039_);
  or _75408_ (_24578_, _24576_, _03983_);
  and _75409_ (_24579_, _05941_, _05272_);
  or _75410_ (_24580_, _24579_, _24574_);
  and _75411_ (_24582_, _24580_, _03570_);
  nor _75412_ (_24583_, _04426_, _24572_);
  and _75413_ (_24584_, _05272_, \oc8051_golden_model_1.ACC [0]);
  or _75414_ (_24585_, _24584_, _24574_);
  and _75415_ (_24586_, _24585_, _04426_);
  or _75416_ (_24587_, _24586_, _24583_);
  and _75417_ (_24588_, _24587_, _04444_);
  or _75418_ (_24589_, _24588_, _03568_);
  or _75419_ (_24590_, _24589_, _24582_);
  and _75420_ (_24591_, _24590_, _24578_);
  or _75421_ (_24593_, _24591_, _03575_);
  or _75422_ (_24594_, _24585_, _03583_);
  and _75423_ (_24595_, _24594_, _09771_);
  and _75424_ (_24596_, _24595_, _24593_);
  and _75425_ (_24597_, _09770_, _24572_);
  or _75426_ (_24598_, _24597_, _24596_);
  and _75427_ (_24599_, _24598_, _09755_);
  nor _75428_ (_24600_, _04109_, _09755_);
  or _75429_ (_24601_, _24600_, _07314_);
  or _75430_ (_24602_, _24601_, _24599_);
  and _75431_ (_24604_, _24602_, _24577_);
  or _75432_ (_24605_, _24604_, _03479_);
  and _75433_ (_24606_, _06715_, _05272_);
  or _75434_ (_24607_, _24574_, _06044_);
  or _75435_ (_24608_, _24607_, _24606_);
  and _75436_ (_24609_, _24608_, _24605_);
  or _75437_ (_24610_, _24609_, _03221_);
  nor _75438_ (_24611_, _11975_, _09751_);
  or _75439_ (_24612_, _24611_, _24574_);
  or _75440_ (_24613_, _24612_, _03474_);
  and _75441_ (_24616_, _24613_, _03438_);
  and _75442_ (_24617_, _24616_, _24610_);
  and _75443_ (_24618_, _05272_, _06202_);
  or _75444_ (_24619_, _24618_, _24574_);
  and _75445_ (_24620_, _24619_, _03437_);
  or _75446_ (_24621_, _24620_, _03636_);
  or _75447_ (_24622_, _24621_, _24617_);
  and _75448_ (_24623_, _11990_, _05272_);
  or _75449_ (_24624_, _24623_, _24574_);
  or _75450_ (_24625_, _24624_, _04499_);
  and _75451_ (_24627_, _24625_, _24622_);
  or _75452_ (_24628_, _24627_, _03769_);
  and _75453_ (_24629_, _11995_, _05272_);
  or _75454_ (_24630_, _24629_, _24574_);
  or _75455_ (_24631_, _24630_, _04501_);
  and _75456_ (_24632_, _24631_, _05769_);
  and _75457_ (_24633_, _24632_, _24628_);
  nand _75458_ (_24634_, _24619_, _04504_);
  nor _75459_ (_24635_, _24634_, _24579_);
  or _75460_ (_24636_, _24635_, _24633_);
  and _75461_ (_24638_, _24636_, _03753_);
  or _75462_ (_24639_, _24574_, _05617_);
  and _75463_ (_24640_, _24585_, _03752_);
  and _75464_ (_24641_, _24640_, _24639_);
  or _75465_ (_24642_, _24641_, _03758_);
  or _75466_ (_24643_, _24642_, _24638_);
  nor _75467_ (_24644_, _11988_, _09751_);
  or _75468_ (_24645_, _24574_, _03759_);
  or _75469_ (_24646_, _24645_, _24644_);
  and _75470_ (_24647_, _24646_, _04517_);
  and _75471_ (_24649_, _24647_, _24643_);
  nor _75472_ (_24650_, _11870_, _09751_);
  or _75473_ (_24651_, _24650_, _24574_);
  and _75474_ (_24652_, _24651_, _03760_);
  or _75475_ (_24653_, _24652_, _17076_);
  or _75476_ (_24654_, _24653_, _24649_);
  or _75477_ (_24655_, _24580_, _03882_);
  and _75478_ (_24656_, _24655_, _42963_);
  and _75479_ (_24657_, _24656_, _24654_);
  or _75480_ (_24658_, _24657_, _24573_);
  and _75481_ (_43307_, _24658_, _41755_);
  not _75482_ (_24660_, \oc8051_golden_model_1.DPL [1]);
  nor _75483_ (_24661_, _42963_, _24660_);
  or _75484_ (_24662_, _05272_, \oc8051_golden_model_1.DPL [1]);
  and _75485_ (_24663_, _12252_, _05272_);
  not _75486_ (_24664_, _24663_);
  and _75487_ (_24665_, _24664_, _24662_);
  or _75488_ (_24666_, _24665_, _04192_);
  nand _75489_ (_24667_, _05272_, _04603_);
  and _75490_ (_24668_, _24667_, _24662_);
  or _75491_ (_24670_, _24668_, _06039_);
  nor _75492_ (_24671_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor _75493_ (_24672_, _24671_, _09775_);
  and _75494_ (_24673_, _24672_, _09770_);
  or _75495_ (_24674_, _24665_, _04444_);
  nand _75496_ (_24675_, _05272_, _03233_);
  and _75497_ (_24676_, _24675_, _24662_);
  and _75498_ (_24677_, _24676_, _04426_);
  nor _75499_ (_24678_, _04426_, _24660_);
  or _75500_ (_24679_, _24678_, _03570_);
  or _75501_ (_24681_, _24679_, _24677_);
  and _75502_ (_24682_, _24681_, _03983_);
  and _75503_ (_24683_, _24682_, _24674_);
  and _75504_ (_24684_, _24668_, _03568_);
  or _75505_ (_24685_, _24684_, _03575_);
  or _75506_ (_24686_, _24685_, _24683_);
  or _75507_ (_24687_, _24676_, _03583_);
  and _75508_ (_24688_, _24687_, _09771_);
  and _75509_ (_24689_, _24688_, _24686_);
  or _75510_ (_24690_, _24689_, _24673_);
  and _75511_ (_24692_, _24690_, _09755_);
  nor _75512_ (_24693_, _04317_, _09755_);
  or _75513_ (_24694_, _24693_, _07314_);
  or _75514_ (_24695_, _24694_, _24692_);
  and _75515_ (_24696_, _24695_, _24670_);
  or _75516_ (_24697_, _24696_, _03479_);
  and _75517_ (_24698_, _24697_, _03474_);
  nor _75518_ (_24699_, _05272_, _24660_);
  and _75519_ (_24700_, _06714_, _05272_);
  or _75520_ (_24701_, _24700_, _24699_);
  or _75521_ (_24703_, _24701_, _06044_);
  and _75522_ (_24704_, _24703_, _24698_);
  nand _75523_ (_24705_, _12176_, _05272_);
  and _75524_ (_24706_, _24662_, _03221_);
  and _75525_ (_24707_, _24706_, _24705_);
  or _75526_ (_24708_, _24707_, _24704_);
  and _75527_ (_24709_, _24708_, _03438_);
  nand _75528_ (_24710_, _05272_, _04317_);
  and _75529_ (_24711_, _24662_, _03437_);
  and _75530_ (_24712_, _24711_, _24710_);
  or _75531_ (_24714_, _24712_, _24709_);
  and _75532_ (_24715_, _24714_, _04499_);
  or _75533_ (_24716_, _12191_, _09751_);
  and _75534_ (_24717_, _24662_, _03636_);
  and _75535_ (_24718_, _24717_, _24716_);
  or _75536_ (_24719_, _24718_, _24715_);
  and _75537_ (_24720_, _24719_, _04501_);
  or _75538_ (_24721_, _12197_, _09751_);
  and _75539_ (_24722_, _24662_, _03769_);
  and _75540_ (_24723_, _24722_, _24721_);
  or _75541_ (_24725_, _24723_, _24720_);
  and _75542_ (_24726_, _24725_, _05769_);
  or _75543_ (_24727_, _12190_, _09751_);
  and _75544_ (_24728_, _24727_, _03754_);
  and _75545_ (_24729_, _24728_, _24662_);
  or _75546_ (_24730_, _24729_, _24726_);
  and _75547_ (_24731_, _24730_, _03753_);
  or _75548_ (_24732_, _24699_, _05569_);
  and _75549_ (_24733_, _24676_, _03752_);
  and _75550_ (_24734_, _24733_, _24732_);
  or _75551_ (_24736_, _24734_, _24731_);
  and _75552_ (_24737_, _24736_, _03759_);
  or _75553_ (_24738_, _24710_, _05569_);
  and _75554_ (_24739_, _24662_, _03758_);
  and _75555_ (_24740_, _24739_, _24738_);
  or _75556_ (_24741_, _24740_, _24737_);
  and _75557_ (_24742_, _24741_, _04517_);
  or _75558_ (_24743_, _24675_, _05569_);
  and _75559_ (_24744_, _24662_, _03760_);
  and _75560_ (_24745_, _24744_, _24743_);
  or _75561_ (_24747_, _24745_, _03790_);
  or _75562_ (_24748_, _24747_, _24742_);
  and _75563_ (_24749_, _24748_, _24666_);
  or _75564_ (_24750_, _24749_, _03520_);
  or _75565_ (_24751_, _24699_, _03521_);
  or _75566_ (_24752_, _24751_, _24663_);
  and _75567_ (_24753_, _24752_, _42963_);
  and _75568_ (_24754_, _24753_, _24750_);
  or _75569_ (_24755_, _24754_, _24661_);
  and _75570_ (_43310_, _24755_, _41755_);
  not _75571_ (_24757_, \oc8051_golden_model_1.DPL [2]);
  nor _75572_ (_24758_, _42963_, _24757_);
  nor _75573_ (_24759_, _05272_, _24757_);
  nor _75574_ (_24760_, _12400_, _09751_);
  or _75575_ (_24761_, _24760_, _24759_);
  and _75576_ (_24762_, _24761_, _03760_);
  and _75577_ (_24763_, _12401_, _05272_);
  or _75578_ (_24764_, _24763_, _24759_);
  and _75579_ (_24765_, _24764_, _03769_);
  and _75580_ (_24766_, _06718_, _05272_);
  or _75581_ (_24768_, _24766_, _24759_);
  and _75582_ (_24769_, _24768_, _03479_);
  nor _75583_ (_24770_, _09775_, \oc8051_golden_model_1.DPL [2]);
  nor _75584_ (_24771_, _24770_, _09776_);
  and _75585_ (_24772_, _24771_, _09770_);
  nor _75586_ (_24773_, _12282_, _09751_);
  or _75587_ (_24774_, _24773_, _24759_);
  or _75588_ (_24775_, _24774_, _04444_);
  and _75589_ (_24776_, _05272_, \oc8051_golden_model_1.ACC [2]);
  or _75590_ (_24777_, _24776_, _24759_);
  and _75591_ (_24779_, _24777_, _04426_);
  nor _75592_ (_24780_, _04426_, _24757_);
  or _75593_ (_24781_, _24780_, _03570_);
  or _75594_ (_24782_, _24781_, _24779_);
  and _75595_ (_24783_, _24782_, _03983_);
  and _75596_ (_24784_, _24783_, _24775_);
  nor _75597_ (_24785_, _09751_, _05026_);
  or _75598_ (_24786_, _24785_, _24759_);
  and _75599_ (_24787_, _24786_, _03568_);
  or _75600_ (_24788_, _24787_, _03575_);
  or _75601_ (_24790_, _24788_, _24784_);
  or _75602_ (_24791_, _24777_, _03583_);
  and _75603_ (_24792_, _24791_, _09771_);
  and _75604_ (_24793_, _24792_, _24790_);
  or _75605_ (_24794_, _24793_, _24772_);
  and _75606_ (_24795_, _24794_, _09755_);
  nor _75607_ (_24796_, _03920_, _09755_);
  or _75608_ (_24797_, _24796_, _07314_);
  or _75609_ (_24798_, _24797_, _24795_);
  or _75610_ (_24799_, _24786_, _06039_);
  and _75611_ (_24801_, _24799_, _06044_);
  and _75612_ (_24802_, _24801_, _24798_);
  or _75613_ (_24803_, _24802_, _03221_);
  or _75614_ (_24804_, _24803_, _24769_);
  nor _75615_ (_24805_, _12384_, _09751_);
  or _75616_ (_24806_, _24759_, _03474_);
  or _75617_ (_24807_, _24806_, _24805_);
  and _75618_ (_24808_, _24807_, _03438_);
  and _75619_ (_24809_, _24808_, _24804_);
  and _75620_ (_24810_, _05272_, _06261_);
  or _75621_ (_24812_, _24810_, _24759_);
  and _75622_ (_24813_, _24812_, _03437_);
  or _75623_ (_24814_, _24813_, _03636_);
  or _75624_ (_24815_, _24814_, _24809_);
  and _75625_ (_24816_, _12273_, _05272_);
  or _75626_ (_24817_, _24816_, _24759_);
  or _75627_ (_24818_, _24817_, _04499_);
  and _75628_ (_24819_, _24818_, _04501_);
  and _75629_ (_24820_, _24819_, _24815_);
  or _75630_ (_24821_, _24820_, _24765_);
  and _75631_ (_24823_, _24821_, _05769_);
  or _75632_ (_24824_, _24759_, _05665_);
  and _75633_ (_24825_, _24824_, _03754_);
  and _75634_ (_24826_, _24825_, _24812_);
  or _75635_ (_24827_, _24826_, _24823_);
  and _75636_ (_24828_, _24827_, _03753_);
  and _75637_ (_24829_, _24777_, _03752_);
  and _75638_ (_24830_, _24829_, _24824_);
  or _75639_ (_24831_, _24830_, _03758_);
  or _75640_ (_24832_, _24831_, _24828_);
  nor _75641_ (_24834_, _12272_, _09751_);
  or _75642_ (_24835_, _24759_, _03759_);
  or _75643_ (_24836_, _24835_, _24834_);
  and _75644_ (_24837_, _24836_, _04517_);
  and _75645_ (_24838_, _24837_, _24832_);
  or _75646_ (_24839_, _24838_, _24762_);
  and _75647_ (_24840_, _24839_, _04192_);
  and _75648_ (_24841_, _24774_, _03790_);
  or _75649_ (_24842_, _24841_, _03520_);
  or _75650_ (_24843_, _24842_, _24840_);
  and _75651_ (_24845_, _12456_, _05272_);
  or _75652_ (_24846_, _24759_, _03521_);
  or _75653_ (_24847_, _24846_, _24845_);
  and _75654_ (_24848_, _24847_, _42963_);
  and _75655_ (_24849_, _24848_, _24843_);
  or _75656_ (_24850_, _24849_, _24758_);
  and _75657_ (_43311_, _24850_, _41755_);
  or _75658_ (_24851_, _42963_, \oc8051_golden_model_1.DPL [3]);
  and _75659_ (_24852_, _24851_, _41755_);
  and _75660_ (_24853_, _09751_, \oc8051_golden_model_1.DPL [3]);
  and _75661_ (_24855_, _12604_, _05272_);
  or _75662_ (_24856_, _24855_, _24853_);
  and _75663_ (_24857_, _24856_, _03769_);
  nor _75664_ (_24858_, _09751_, _04843_);
  or _75665_ (_24859_, _24858_, _24853_);
  or _75666_ (_24860_, _24859_, _06039_);
  nor _75667_ (_24861_, _09776_, \oc8051_golden_model_1.DPL [3]);
  nor _75668_ (_24862_, _24861_, _09777_);
  and _75669_ (_24863_, _24862_, _09770_);
  nor _75670_ (_24864_, _12486_, _09751_);
  or _75671_ (_24866_, _24864_, _24853_);
  or _75672_ (_24867_, _24866_, _04444_);
  and _75673_ (_24868_, _05272_, \oc8051_golden_model_1.ACC [3]);
  or _75674_ (_24869_, _24868_, _24853_);
  and _75675_ (_24870_, _24869_, _04426_);
  and _75676_ (_24871_, _04427_, \oc8051_golden_model_1.DPL [3]);
  or _75677_ (_24872_, _24871_, _03570_);
  or _75678_ (_24873_, _24872_, _24870_);
  and _75679_ (_24874_, _24873_, _03983_);
  and _75680_ (_24875_, _24874_, _24867_);
  and _75681_ (_24877_, _24859_, _03568_);
  or _75682_ (_24878_, _24877_, _03575_);
  or _75683_ (_24879_, _24878_, _24875_);
  or _75684_ (_24880_, _24869_, _03583_);
  and _75685_ (_24881_, _24880_, _09771_);
  and _75686_ (_24882_, _24881_, _24879_);
  or _75687_ (_24883_, _24882_, _24863_);
  and _75688_ (_24884_, _24883_, _09755_);
  nor _75689_ (_24885_, _03742_, _09755_);
  or _75690_ (_24886_, _24885_, _07314_);
  or _75691_ (_24888_, _24886_, _24884_);
  and _75692_ (_24889_, _24888_, _24860_);
  or _75693_ (_24890_, _24889_, _03479_);
  and _75694_ (_24891_, _06717_, _05272_);
  or _75695_ (_24892_, _24853_, _06044_);
  or _75696_ (_24893_, _24892_, _24891_);
  and _75697_ (_24894_, _24893_, _03474_);
  and _75698_ (_24895_, _24894_, _24890_);
  nor _75699_ (_24896_, _12583_, _09751_);
  or _75700_ (_24897_, _24896_, _24853_);
  and _75701_ (_24899_, _24897_, _03221_);
  or _75702_ (_24900_, _24899_, _03437_);
  or _75703_ (_24901_, _24900_, _24895_);
  and _75704_ (_24902_, _05272_, _06217_);
  or _75705_ (_24903_, _24902_, _24853_);
  or _75706_ (_24904_, _24903_, _03438_);
  and _75707_ (_24905_, _24904_, _24901_);
  or _75708_ (_24906_, _24905_, _03636_);
  and _75709_ (_24907_, _12598_, _05272_);
  or _75710_ (_24908_, _24907_, _24853_);
  or _75711_ (_24910_, _24908_, _04499_);
  and _75712_ (_24911_, _24910_, _04501_);
  and _75713_ (_24912_, _24911_, _24906_);
  or _75714_ (_24913_, _24912_, _24857_);
  and _75715_ (_24914_, _24913_, _05769_);
  or _75716_ (_24915_, _24853_, _05521_);
  and _75717_ (_24916_, _24915_, _03754_);
  and _75718_ (_24917_, _24916_, _24903_);
  or _75719_ (_24918_, _24917_, _24914_);
  and _75720_ (_24919_, _24918_, _03753_);
  and _75721_ (_24921_, _24869_, _03752_);
  and _75722_ (_24922_, _24921_, _24915_);
  or _75723_ (_24923_, _24922_, _03758_);
  or _75724_ (_24924_, _24923_, _24919_);
  nor _75725_ (_24925_, _12597_, _09751_);
  or _75726_ (_24926_, _24853_, _03759_);
  or _75727_ (_24927_, _24926_, _24925_);
  and _75728_ (_24928_, _24927_, _04517_);
  and _75729_ (_24929_, _24928_, _24924_);
  nor _75730_ (_24930_, _12603_, _09751_);
  or _75731_ (_24932_, _24930_, _24853_);
  and _75732_ (_24933_, _24932_, _03760_);
  or _75733_ (_24934_, _24933_, _03790_);
  or _75734_ (_24935_, _24934_, _24929_);
  or _75735_ (_24936_, _24866_, _04192_);
  and _75736_ (_24937_, _24936_, _03521_);
  and _75737_ (_24938_, _24937_, _24935_);
  and _75738_ (_24939_, _12658_, _05272_);
  or _75739_ (_24940_, _24939_, _24853_);
  and _75740_ (_24941_, _24940_, _03520_);
  or _75741_ (_24943_, _24941_, _42967_);
  or _75742_ (_24944_, _24943_, _24938_);
  and _75743_ (_43312_, _24944_, _24852_);
  or _75744_ (_24945_, _42963_, \oc8051_golden_model_1.DPL [4]);
  and _75745_ (_24946_, _24945_, _41755_);
  and _75746_ (_24947_, _09751_, \oc8051_golden_model_1.DPL [4]);
  and _75747_ (_24948_, _12844_, _05272_);
  or _75748_ (_24949_, _24948_, _24947_);
  and _75749_ (_24950_, _24949_, _03769_);
  nor _75750_ (_24951_, _05712_, _09751_);
  or _75751_ (_24953_, _24951_, _24947_);
  or _75752_ (_24954_, _24953_, _06039_);
  nor _75753_ (_24955_, _12733_, _09751_);
  or _75754_ (_24956_, _24955_, _24947_);
  or _75755_ (_24957_, _24956_, _04444_);
  and _75756_ (_24958_, _05272_, \oc8051_golden_model_1.ACC [4]);
  or _75757_ (_24959_, _24958_, _24947_);
  and _75758_ (_24960_, _24959_, _04426_);
  and _75759_ (_24961_, _04427_, \oc8051_golden_model_1.DPL [4]);
  or _75760_ (_24962_, _24961_, _03570_);
  or _75761_ (_24964_, _24962_, _24960_);
  and _75762_ (_24965_, _24964_, _03983_);
  and _75763_ (_24966_, _24965_, _24957_);
  and _75764_ (_24967_, _24953_, _03568_);
  or _75765_ (_24968_, _24967_, _03575_);
  or _75766_ (_24969_, _24968_, _24966_);
  or _75767_ (_24970_, _24959_, _03583_);
  and _75768_ (_24971_, _24970_, _09771_);
  and _75769_ (_24972_, _24971_, _24969_);
  nor _75770_ (_24973_, _09777_, \oc8051_golden_model_1.DPL [4]);
  nor _75771_ (_24975_, _24973_, _09778_);
  and _75772_ (_24976_, _24975_, _09770_);
  or _75773_ (_24977_, _24976_, _24972_);
  and _75774_ (_24978_, _24977_, _09755_);
  nor _75775_ (_24979_, _06195_, _09755_);
  or _75776_ (_24980_, _24979_, _07314_);
  or _75777_ (_24981_, _24980_, _24978_);
  and _75778_ (_24982_, _24981_, _24954_);
  or _75779_ (_24983_, _24982_, _03479_);
  and _75780_ (_24984_, _06722_, _05272_);
  or _75781_ (_24986_, _24947_, _06044_);
  or _75782_ (_24987_, _24986_, _24984_);
  and _75783_ (_24988_, _24987_, _03474_);
  and _75784_ (_24989_, _24988_, _24983_);
  nor _75785_ (_24990_, _12827_, _09751_);
  or _75786_ (_24991_, _24990_, _24947_);
  and _75787_ (_24992_, _24991_, _03221_);
  or _75788_ (_24993_, _24992_, _03437_);
  or _75789_ (_24994_, _24993_, _24989_);
  and _75790_ (_24995_, _06233_, _05272_);
  or _75791_ (_24997_, _24995_, _24947_);
  or _75792_ (_24998_, _24997_, _03438_);
  and _75793_ (_24999_, _24998_, _24994_);
  or _75794_ (_25000_, _24999_, _03636_);
  and _75795_ (_25001_, _12711_, _05272_);
  or _75796_ (_25002_, _25001_, _24947_);
  or _75797_ (_25003_, _25002_, _04499_);
  and _75798_ (_25004_, _25003_, _04501_);
  and _75799_ (_25005_, _25004_, _25000_);
  or _75800_ (_25006_, _25005_, _24950_);
  and _75801_ (_25008_, _25006_, _05769_);
  or _75802_ (_25009_, _24947_, _05761_);
  and _75803_ (_25010_, _25009_, _03754_);
  and _75804_ (_25011_, _25010_, _24997_);
  or _75805_ (_25012_, _25011_, _25008_);
  and _75806_ (_25013_, _25012_, _03753_);
  and _75807_ (_25014_, _24959_, _03752_);
  and _75808_ (_25015_, _25014_, _25009_);
  or _75809_ (_25016_, _25015_, _03758_);
  or _75810_ (_25017_, _25016_, _25013_);
  nor _75811_ (_25019_, _12710_, _09751_);
  or _75812_ (_25020_, _24947_, _03759_);
  or _75813_ (_25021_, _25020_, _25019_);
  and _75814_ (_25022_, _25021_, _04517_);
  and _75815_ (_25023_, _25022_, _25017_);
  nor _75816_ (_25024_, _12843_, _09751_);
  or _75817_ (_25025_, _25024_, _24947_);
  and _75818_ (_25026_, _25025_, _03760_);
  or _75819_ (_25027_, _25026_, _03790_);
  or _75820_ (_25028_, _25027_, _25023_);
  or _75821_ (_25030_, _24956_, _04192_);
  and _75822_ (_25031_, _25030_, _03521_);
  and _75823_ (_25032_, _25031_, _25028_);
  and _75824_ (_25033_, _12893_, _05272_);
  or _75825_ (_25034_, _25033_, _24947_);
  and _75826_ (_25035_, _25034_, _03520_);
  or _75827_ (_25036_, _25035_, _42967_);
  or _75828_ (_25037_, _25036_, _25032_);
  and _75829_ (_43313_, _25037_, _24946_);
  or _75830_ (_25038_, _42963_, \oc8051_golden_model_1.DPL [5]);
  and _75831_ (_25040_, _25038_, _41755_);
  and _75832_ (_25041_, _09751_, \oc8051_golden_model_1.DPL [5]);
  and _75833_ (_25042_, _13042_, _05272_);
  or _75834_ (_25043_, _25042_, _25041_);
  and _75835_ (_25044_, _25043_, _03769_);
  nor _75836_ (_25045_, _05422_, _09751_);
  or _75837_ (_25046_, _25045_, _25041_);
  or _75838_ (_25047_, _25046_, _06039_);
  nor _75839_ (_25048_, _12930_, _09751_);
  or _75840_ (_25049_, _25048_, _25041_);
  or _75841_ (_25051_, _25049_, _04444_);
  and _75842_ (_25052_, _05272_, \oc8051_golden_model_1.ACC [5]);
  or _75843_ (_25053_, _25052_, _25041_);
  and _75844_ (_25054_, _25053_, _04426_);
  and _75845_ (_25055_, _04427_, \oc8051_golden_model_1.DPL [5]);
  or _75846_ (_25056_, _25055_, _03570_);
  or _75847_ (_25057_, _25056_, _25054_);
  and _75848_ (_25058_, _25057_, _03983_);
  and _75849_ (_25059_, _25058_, _25051_);
  and _75850_ (_25060_, _25046_, _03568_);
  or _75851_ (_25062_, _25060_, _03575_);
  or _75852_ (_25063_, _25062_, _25059_);
  or _75853_ (_25064_, _25053_, _03583_);
  and _75854_ (_25065_, _25064_, _09771_);
  and _75855_ (_25066_, _25065_, _25063_);
  nor _75856_ (_25067_, _09778_, \oc8051_golden_model_1.DPL [5]);
  nor _75857_ (_25068_, _25067_, _09779_);
  and _75858_ (_25069_, _25068_, _09770_);
  or _75859_ (_25070_, _25069_, _25066_);
  and _75860_ (_25071_, _25070_, _09755_);
  nor _75861_ (_25073_, _06164_, _09755_);
  or _75862_ (_25074_, _25073_, _07314_);
  or _75863_ (_25075_, _25074_, _25071_);
  and _75864_ (_25076_, _25075_, _25047_);
  or _75865_ (_25077_, _25076_, _03479_);
  and _75866_ (_25078_, _06721_, _05272_);
  or _75867_ (_25079_, _25041_, _06044_);
  or _75868_ (_25080_, _25079_, _25078_);
  and _75869_ (_25081_, _25080_, _03474_);
  and _75870_ (_25082_, _25081_, _25077_);
  nor _75871_ (_25084_, _13021_, _09751_);
  or _75872_ (_25085_, _25084_, _25041_);
  and _75873_ (_25086_, _25085_, _03221_);
  or _75874_ (_25087_, _25086_, _03437_);
  or _75875_ (_25088_, _25087_, _25082_);
  and _75876_ (_25089_, _06211_, _05272_);
  or _75877_ (_25090_, _25089_, _25041_);
  or _75878_ (_25091_, _25090_, _03438_);
  and _75879_ (_25092_, _25091_, _25088_);
  or _75880_ (_25093_, _25092_, _03636_);
  and _75881_ (_25094_, _13036_, _05272_);
  or _75882_ (_25095_, _25094_, _25041_);
  or _75883_ (_25096_, _25095_, _04499_);
  and _75884_ (_25097_, _25096_, _04501_);
  and _75885_ (_25098_, _25097_, _25093_);
  or _75886_ (_25099_, _25098_, _25044_);
  and _75887_ (_25100_, _25099_, _05769_);
  or _75888_ (_25101_, _25041_, _05472_);
  and _75889_ (_25102_, _25101_, _03754_);
  and _75890_ (_25103_, _25102_, _25090_);
  or _75891_ (_25106_, _25103_, _25100_);
  and _75892_ (_25107_, _25106_, _03753_);
  and _75893_ (_25108_, _25053_, _03752_);
  and _75894_ (_25109_, _25108_, _25101_);
  or _75895_ (_25110_, _25109_, _03758_);
  or _75896_ (_25111_, _25110_, _25107_);
  nor _75897_ (_25112_, _13035_, _09751_);
  or _75898_ (_25113_, _25041_, _03759_);
  or _75899_ (_25114_, _25113_, _25112_);
  and _75900_ (_25115_, _25114_, _04517_);
  and _75901_ (_25117_, _25115_, _25111_);
  nor _75902_ (_25118_, _13041_, _09751_);
  or _75903_ (_25119_, _25118_, _25041_);
  and _75904_ (_25120_, _25119_, _03760_);
  or _75905_ (_25121_, _25120_, _03790_);
  or _75906_ (_25122_, _25121_, _25117_);
  or _75907_ (_25123_, _25049_, _04192_);
  and _75908_ (_25124_, _25123_, _03521_);
  and _75909_ (_25125_, _25124_, _25122_);
  and _75910_ (_25126_, _13097_, _05272_);
  or _75911_ (_25128_, _25126_, _25041_);
  and _75912_ (_25129_, _25128_, _03520_);
  or _75913_ (_25130_, _25129_, _42967_);
  or _75914_ (_25131_, _25130_, _25125_);
  and _75915_ (_43314_, _25131_, _25040_);
  or _75916_ (_25132_, _42963_, \oc8051_golden_model_1.DPL [6]);
  and _75917_ (_25133_, _25132_, _41755_);
  and _75918_ (_25134_, _09751_, \oc8051_golden_model_1.DPL [6]);
  and _75919_ (_25135_, _13259_, _05272_);
  or _75920_ (_25136_, _25135_, _25134_);
  and _75921_ (_25137_, _25136_, _03769_);
  nor _75922_ (_25138_, _05327_, _09751_);
  or _75923_ (_25139_, _25138_, _25134_);
  or _75924_ (_25140_, _25139_, _06039_);
  nor _75925_ (_25141_, _13122_, _09751_);
  or _75926_ (_25142_, _25141_, _25134_);
  or _75927_ (_25143_, _25142_, _04444_);
  and _75928_ (_25144_, _05272_, \oc8051_golden_model_1.ACC [6]);
  or _75929_ (_25145_, _25144_, _25134_);
  and _75930_ (_25146_, _25145_, _04426_);
  and _75931_ (_25149_, _04427_, \oc8051_golden_model_1.DPL [6]);
  or _75932_ (_25150_, _25149_, _03570_);
  or _75933_ (_25151_, _25150_, _25146_);
  and _75934_ (_25152_, _25151_, _03983_);
  and _75935_ (_25153_, _25152_, _25143_);
  and _75936_ (_25154_, _25139_, _03568_);
  or _75937_ (_25155_, _25154_, _03575_);
  or _75938_ (_25156_, _25155_, _25153_);
  or _75939_ (_25157_, _25145_, _03583_);
  and _75940_ (_25158_, _25157_, _09771_);
  and _75941_ (_25160_, _25158_, _25156_);
  nor _75942_ (_25161_, _09779_, \oc8051_golden_model_1.DPL [6]);
  nor _75943_ (_25162_, _25161_, _09780_);
  and _75944_ (_25163_, _25162_, _09770_);
  or _75945_ (_25164_, _25163_, _25160_);
  and _75946_ (_25165_, _25164_, _09755_);
  nor _75947_ (_25166_, _06132_, _09755_);
  or _75948_ (_25167_, _25166_, _07314_);
  or _75949_ (_25168_, _25167_, _25165_);
  and _75950_ (_25169_, _25168_, _25140_);
  or _75951_ (_25170_, _25169_, _03479_);
  and _75952_ (_25171_, _06713_, _05272_);
  or _75953_ (_25172_, _25134_, _06044_);
  or _75954_ (_25173_, _25172_, _25171_);
  and _75955_ (_25174_, _25173_, _03474_);
  and _75956_ (_25175_, _25174_, _25170_);
  nor _75957_ (_25176_, _13237_, _09751_);
  or _75958_ (_25177_, _25176_, _25134_);
  and _75959_ (_25178_, _25177_, _03221_);
  or _75960_ (_25179_, _25178_, _03437_);
  or _75961_ (_25182_, _25179_, _25175_);
  and _75962_ (_25183_, _13244_, _05272_);
  or _75963_ (_25184_, _25183_, _25134_);
  or _75964_ (_25185_, _25184_, _03438_);
  and _75965_ (_25186_, _25185_, _25182_);
  or _75966_ (_25187_, _25186_, _03636_);
  and _75967_ (_25188_, _13253_, _05272_);
  or _75968_ (_25189_, _25188_, _25134_);
  or _75969_ (_25190_, _25189_, _04499_);
  and _75970_ (_25191_, _25190_, _04501_);
  and _75971_ (_25193_, _25191_, _25187_);
  or _75972_ (_25194_, _25193_, _25137_);
  and _75973_ (_25195_, _25194_, _05769_);
  or _75974_ (_25196_, _25134_, _05377_);
  and _75975_ (_25197_, _25196_, _03754_);
  and _75976_ (_25198_, _25197_, _25184_);
  or _75977_ (_25199_, _25198_, _25195_);
  and _75978_ (_25200_, _25199_, _03753_);
  and _75979_ (_25201_, _25145_, _03752_);
  and _75980_ (_25202_, _25201_, _25196_);
  or _75981_ (_25204_, _25202_, _03758_);
  or _75982_ (_25205_, _25204_, _25200_);
  nor _75983_ (_25206_, _13251_, _09751_);
  or _75984_ (_25207_, _25134_, _03759_);
  or _75985_ (_25208_, _25207_, _25206_);
  and _75986_ (_25209_, _25208_, _04517_);
  and _75987_ (_25210_, _25209_, _25205_);
  nor _75988_ (_25211_, _13258_, _09751_);
  or _75989_ (_25212_, _25211_, _25134_);
  and _75990_ (_25213_, _25212_, _03760_);
  or _75991_ (_25215_, _25213_, _03790_);
  or _75992_ (_25216_, _25215_, _25210_);
  or _75993_ (_25217_, _25142_, _04192_);
  and _75994_ (_25218_, _25217_, _03521_);
  and _75995_ (_25219_, _25218_, _25216_);
  and _75996_ (_25220_, _13312_, _05272_);
  or _75997_ (_25221_, _25220_, _25134_);
  and _75998_ (_25222_, _25221_, _03520_);
  or _75999_ (_25223_, _25222_, _42967_);
  or _76000_ (_25224_, _25223_, _25219_);
  and _76001_ (_43315_, _25224_, _25133_);
  nor _76002_ (_25225_, _42963_, _10476_);
  nor _76003_ (_25226_, _05266_, _10476_);
  and _76004_ (_25227_, _05266_, _04419_);
  or _76005_ (_25228_, _25227_, _25226_);
  or _76006_ (_25229_, _25228_, _06039_);
  nor _76007_ (_25230_, _09782_, \oc8051_golden_model_1.DPH [0]);
  nor _76008_ (_25231_, _25230_, _09869_);
  and _76009_ (_25232_, _25231_, _09770_);
  or _76010_ (_25233_, _25228_, _03983_);
  and _76011_ (_25236_, _05941_, _05266_);
  or _76012_ (_25237_, _25236_, _25226_);
  and _76013_ (_25238_, _25237_, _03570_);
  nor _76014_ (_25239_, _04426_, _10476_);
  and _76015_ (_25240_, _05266_, \oc8051_golden_model_1.ACC [0]);
  or _76016_ (_25241_, _25240_, _25226_);
  and _76017_ (_25242_, _25241_, _04426_);
  or _76018_ (_25243_, _25242_, _25239_);
  and _76019_ (_25244_, _25243_, _04444_);
  or _76020_ (_25245_, _25244_, _03568_);
  or _76021_ (_25247_, _25245_, _25238_);
  and _76022_ (_25248_, _25247_, _25233_);
  or _76023_ (_25249_, _25248_, _03575_);
  or _76024_ (_25250_, _25241_, _03583_);
  and _76025_ (_25251_, _25250_, _09771_);
  and _76026_ (_25252_, _25251_, _25249_);
  or _76027_ (_25253_, _25252_, _25232_);
  and _76028_ (_25254_, _25253_, _09755_);
  nor _76029_ (_25255_, _09755_, _03471_);
  or _76030_ (_25256_, _25255_, _07314_);
  or _76031_ (_25258_, _25256_, _25254_);
  and _76032_ (_25259_, _25258_, _25229_);
  or _76033_ (_25260_, _25259_, _03479_);
  and _76034_ (_25261_, _06715_, _05266_);
  or _76035_ (_25262_, _25226_, _06044_);
  or _76036_ (_25263_, _25262_, _25261_);
  and _76037_ (_25264_, _25263_, _25260_);
  or _76038_ (_25265_, _25264_, _03221_);
  nor _76039_ (_25266_, _11975_, _09848_);
  or _76040_ (_25267_, _25266_, _25226_);
  or _76041_ (_25269_, _25267_, _03474_);
  and _76042_ (_25270_, _25269_, _03438_);
  and _76043_ (_25271_, _25270_, _25265_);
  and _76044_ (_25272_, _05266_, _06202_);
  or _76045_ (_25273_, _25272_, _25226_);
  and _76046_ (_25274_, _25273_, _03437_);
  or _76047_ (_25275_, _25274_, _03636_);
  or _76048_ (_25276_, _25275_, _25271_);
  and _76049_ (_25277_, _11990_, _05266_);
  or _76050_ (_25278_, _25277_, _25226_);
  or _76051_ (_25280_, _25278_, _04499_);
  and _76052_ (_25281_, _25280_, _25276_);
  or _76053_ (_25282_, _25281_, _03769_);
  and _76054_ (_25283_, _11995_, _05266_);
  or _76055_ (_25284_, _25283_, _25226_);
  or _76056_ (_25285_, _25284_, _04501_);
  and _76057_ (_25286_, _25285_, _05769_);
  and _76058_ (_25287_, _25286_, _25282_);
  nand _76059_ (_25288_, _25273_, _04504_);
  nor _76060_ (_25289_, _25288_, _25236_);
  or _76061_ (_25291_, _25289_, _25287_);
  and _76062_ (_25292_, _25291_, _03753_);
  or _76063_ (_25293_, _25226_, _05617_);
  and _76064_ (_25294_, _25241_, _03752_);
  and _76065_ (_25295_, _25294_, _25293_);
  or _76066_ (_25296_, _25295_, _03758_);
  or _76067_ (_25297_, _25296_, _25292_);
  nor _76068_ (_25298_, _11988_, _09848_);
  or _76069_ (_25299_, _25226_, _03759_);
  or _76070_ (_25300_, _25299_, _25298_);
  and _76071_ (_25302_, _25300_, _04517_);
  and _76072_ (_25303_, _25302_, _25297_);
  nor _76073_ (_25304_, _11870_, _09848_);
  or _76074_ (_25305_, _25304_, _25226_);
  and _76075_ (_25306_, _25305_, _03760_);
  or _76076_ (_25307_, _25306_, _17076_);
  or _76077_ (_25308_, _25307_, _25303_);
  or _76078_ (_25309_, _25237_, _03882_);
  and _76079_ (_25310_, _25309_, _42963_);
  and _76080_ (_25311_, _25310_, _25308_);
  or _76081_ (_25313_, _25311_, _25225_);
  and _76082_ (_43318_, _25313_, _41755_);
  not _76083_ (_25314_, \oc8051_golden_model_1.DPH [1]);
  nor _76084_ (_25315_, _42963_, _25314_);
  and _76085_ (_25316_, _12252_, _05266_);
  not _76086_ (_25317_, _25316_);
  or _76087_ (_25318_, _05266_, \oc8051_golden_model_1.DPH [1]);
  and _76088_ (_25319_, _25318_, _25317_);
  or _76089_ (_25320_, _25319_, _04192_);
  nor _76090_ (_25321_, _05266_, _25314_);
  nor _76091_ (_25323_, _09848_, _04603_);
  or _76092_ (_25324_, _25323_, _25321_);
  or _76093_ (_25325_, _25324_, _03983_);
  and _76094_ (_25326_, _25319_, _03570_);
  nand _76095_ (_25327_, _05266_, _03233_);
  and _76096_ (_25328_, _25327_, _25318_);
  and _76097_ (_25329_, _25328_, _04426_);
  nor _76098_ (_25330_, _04426_, _25314_);
  or _76099_ (_25331_, _25330_, _25329_);
  and _76100_ (_25332_, _25331_, _04444_);
  or _76101_ (_25334_, _25332_, _03568_);
  or _76102_ (_25335_, _25334_, _25326_);
  and _76103_ (_25336_, _25335_, _25325_);
  or _76104_ (_25337_, _25336_, _03575_);
  or _76105_ (_25338_, _25328_, _03583_);
  and _76106_ (_25339_, _25338_, _09771_);
  and _76107_ (_25340_, _25339_, _25337_);
  nor _76108_ (_25341_, _09869_, \oc8051_golden_model_1.DPH [1]);
  nor _76109_ (_25342_, _25341_, _09870_);
  and _76110_ (_25343_, _25342_, _09770_);
  or _76111_ (_25345_, _25343_, _25340_);
  and _76112_ (_25346_, _25345_, _09755_);
  nor _76113_ (_25347_, _04284_, _09755_);
  or _76114_ (_25348_, _25347_, _07314_);
  or _76115_ (_25349_, _25348_, _25346_);
  or _76116_ (_25350_, _25324_, _06039_);
  and _76117_ (_25351_, _25350_, _25349_);
  or _76118_ (_25352_, _25351_, _03479_);
  and _76119_ (_25353_, _06714_, _05266_);
  or _76120_ (_25354_, _25321_, _06044_);
  or _76121_ (_25355_, _25354_, _25353_);
  and _76122_ (_25356_, _25355_, _03474_);
  and _76123_ (_25357_, _25356_, _25352_);
  nand _76124_ (_25358_, _12176_, _05266_);
  and _76125_ (_25359_, _25318_, _03221_);
  and _76126_ (_25360_, _25359_, _25358_);
  or _76127_ (_25361_, _25360_, _25357_);
  and _76128_ (_25362_, _25361_, _03438_);
  nand _76129_ (_25363_, _05266_, _04317_);
  and _76130_ (_25364_, _25318_, _03437_);
  and _76131_ (_25367_, _25364_, _25363_);
  or _76132_ (_25368_, _25367_, _25362_);
  and _76133_ (_25369_, _25368_, _04499_);
  or _76134_ (_25370_, _12191_, _09848_);
  and _76135_ (_25371_, _25318_, _03636_);
  and _76136_ (_25372_, _25371_, _25370_);
  or _76137_ (_25373_, _25372_, _25369_);
  and _76138_ (_25374_, _25373_, _04501_);
  or _76139_ (_25375_, _12197_, _09848_);
  and _76140_ (_25376_, _25318_, _03769_);
  and _76141_ (_25378_, _25376_, _25375_);
  or _76142_ (_25379_, _25378_, _25374_);
  and _76143_ (_25380_, _25379_, _05769_);
  or _76144_ (_25381_, _12190_, _09848_);
  and _76145_ (_25382_, _25381_, _03754_);
  and _76146_ (_25383_, _25382_, _25318_);
  or _76147_ (_25384_, _25383_, _25380_);
  and _76148_ (_25385_, _25384_, _03753_);
  or _76149_ (_25386_, _25321_, _05569_);
  and _76150_ (_25387_, _25328_, _03752_);
  and _76151_ (_25389_, _25387_, _25386_);
  or _76152_ (_25390_, _25389_, _25385_);
  and _76153_ (_25391_, _25390_, _03759_);
  or _76154_ (_25392_, _25363_, _05569_);
  and _76155_ (_25393_, _25318_, _03758_);
  and _76156_ (_25394_, _25393_, _25392_);
  or _76157_ (_25395_, _25394_, _25391_);
  and _76158_ (_25396_, _25395_, _04517_);
  nand _76159_ (_25397_, _12196_, _05266_);
  and _76160_ (_25398_, _25397_, _03760_);
  and _76161_ (_25400_, _25398_, _25318_);
  or _76162_ (_25401_, _25400_, _03790_);
  or _76163_ (_25402_, _25401_, _25396_);
  and _76164_ (_25403_, _25402_, _25320_);
  or _76165_ (_25404_, _25403_, _03520_);
  or _76166_ (_25405_, _25321_, _03521_);
  or _76167_ (_25406_, _25405_, _25316_);
  and _76168_ (_25407_, _25406_, _42963_);
  and _76169_ (_25408_, _25407_, _25404_);
  or _76170_ (_25409_, _25408_, _25315_);
  and _76171_ (_43319_, _25409_, _41755_);
  not _76172_ (_25411_, \oc8051_golden_model_1.DPH [2]);
  nor _76173_ (_25412_, _42963_, _25411_);
  nor _76174_ (_25413_, _05266_, _25411_);
  nor _76175_ (_25414_, _12400_, _09848_);
  or _76176_ (_25415_, _25414_, _25413_);
  and _76177_ (_25416_, _25415_, _03760_);
  and _76178_ (_25417_, _12401_, _05266_);
  or _76179_ (_25418_, _25417_, _25413_);
  and _76180_ (_25419_, _25418_, _03769_);
  and _76181_ (_25421_, _06718_, _05266_);
  or _76182_ (_25422_, _25421_, _25413_);
  and _76183_ (_25423_, _25422_, _03479_);
  nor _76184_ (_25424_, _12282_, _09848_);
  or _76185_ (_25425_, _25424_, _25413_);
  or _76186_ (_25426_, _25425_, _04444_);
  and _76187_ (_25427_, _05266_, \oc8051_golden_model_1.ACC [2]);
  or _76188_ (_25428_, _25427_, _25413_);
  and _76189_ (_25429_, _25428_, _04426_);
  nor _76190_ (_25430_, _04426_, _25411_);
  or _76191_ (_25432_, _25430_, _03570_);
  or _76192_ (_25433_, _25432_, _25429_);
  and _76193_ (_25434_, _25433_, _03983_);
  and _76194_ (_25435_, _25434_, _25426_);
  nor _76195_ (_25436_, _09848_, _05026_);
  or _76196_ (_25437_, _25436_, _25413_);
  and _76197_ (_25438_, _25437_, _03568_);
  or _76198_ (_25439_, _25438_, _03575_);
  or _76199_ (_25440_, _25439_, _25435_);
  or _76200_ (_25441_, _25428_, _03583_);
  and _76201_ (_25443_, _25441_, _09771_);
  and _76202_ (_25444_, _25443_, _25440_);
  or _76203_ (_25445_, _09870_, \oc8051_golden_model_1.DPH [2]);
  nor _76204_ (_25446_, _09871_, _09771_);
  and _76205_ (_25447_, _25446_, _25445_);
  or _76206_ (_25448_, _25447_, _25444_);
  and _76207_ (_25449_, _25448_, _09755_);
  nor _76208_ (_25450_, _03877_, _09755_);
  or _76209_ (_25451_, _25450_, _07314_);
  or _76210_ (_25452_, _25451_, _25449_);
  or _76211_ (_25454_, _25437_, _06039_);
  and _76212_ (_25455_, _25454_, _06044_);
  and _76213_ (_25456_, _25455_, _25452_);
  or _76214_ (_25457_, _25456_, _03221_);
  or _76215_ (_25458_, _25457_, _25423_);
  nor _76216_ (_25459_, _12384_, _09848_);
  or _76217_ (_25460_, _25413_, _03474_);
  or _76218_ (_25461_, _25460_, _25459_);
  and _76219_ (_25462_, _25461_, _03438_);
  and _76220_ (_25463_, _25462_, _25458_);
  and _76221_ (_25465_, _05266_, _06261_);
  or _76222_ (_25466_, _25465_, _25413_);
  and _76223_ (_25467_, _25466_, _03437_);
  or _76224_ (_25468_, _25467_, _03636_);
  or _76225_ (_25469_, _25468_, _25463_);
  and _76226_ (_25470_, _12273_, _05266_);
  or _76227_ (_25471_, _25470_, _25413_);
  or _76228_ (_25472_, _25471_, _04499_);
  and _76229_ (_25473_, _25472_, _04501_);
  and _76230_ (_25474_, _25473_, _25469_);
  or _76231_ (_25476_, _25474_, _25419_);
  and _76232_ (_25477_, _25476_, _05769_);
  or _76233_ (_25478_, _25413_, _05665_);
  and _76234_ (_25479_, _25478_, _03754_);
  and _76235_ (_25480_, _25479_, _25466_);
  or _76236_ (_25481_, _25480_, _25477_);
  and _76237_ (_25482_, _25481_, _03753_);
  and _76238_ (_25483_, _25428_, _03752_);
  and _76239_ (_25484_, _25483_, _25478_);
  or _76240_ (_25485_, _25484_, _03758_);
  or _76241_ (_25487_, _25485_, _25482_);
  nor _76242_ (_25488_, _12272_, _09848_);
  or _76243_ (_25489_, _25413_, _03759_);
  or _76244_ (_25490_, _25489_, _25488_);
  and _76245_ (_25491_, _25490_, _04517_);
  and _76246_ (_25492_, _25491_, _25487_);
  or _76247_ (_25493_, _25492_, _25416_);
  and _76248_ (_25494_, _25493_, _04192_);
  and _76249_ (_25495_, _25425_, _03790_);
  or _76250_ (_25496_, _25495_, _03520_);
  or _76251_ (_25498_, _25496_, _25494_);
  and _76252_ (_25499_, _12456_, _05266_);
  or _76253_ (_25500_, _25413_, _03521_);
  or _76254_ (_25501_, _25500_, _25499_);
  and _76255_ (_25502_, _25501_, _42963_);
  and _76256_ (_25503_, _25502_, _25498_);
  or _76257_ (_25504_, _25503_, _25412_);
  and _76258_ (_43320_, _25504_, _41755_);
  or _76259_ (_25505_, _42963_, \oc8051_golden_model_1.DPH [3]);
  and _76260_ (_25506_, _25505_, _41755_);
  and _76261_ (_25508_, _09848_, \oc8051_golden_model_1.DPH [3]);
  and _76262_ (_25509_, _12604_, _05266_);
  or _76263_ (_25510_, _25509_, _25508_);
  and _76264_ (_25511_, _25510_, _03769_);
  nor _76265_ (_25512_, _09848_, _04843_);
  or _76266_ (_25513_, _25512_, _25508_);
  or _76267_ (_25514_, _25513_, _06039_);
  nor _76268_ (_25515_, _12486_, _09848_);
  or _76269_ (_25516_, _25515_, _25508_);
  or _76270_ (_25517_, _25516_, _04444_);
  and _76271_ (_25519_, _05266_, \oc8051_golden_model_1.ACC [3]);
  or _76272_ (_25520_, _25519_, _25508_);
  and _76273_ (_25521_, _25520_, _04426_);
  and _76274_ (_25522_, _04427_, \oc8051_golden_model_1.DPH [3]);
  or _76275_ (_25523_, _25522_, _03570_);
  or _76276_ (_25524_, _25523_, _25521_);
  and _76277_ (_25525_, _25524_, _03983_);
  and _76278_ (_25526_, _25525_, _25517_);
  and _76279_ (_25527_, _25513_, _03568_);
  or _76280_ (_25528_, _25527_, _03575_);
  or _76281_ (_25529_, _25528_, _25526_);
  or _76282_ (_25530_, _25520_, _03583_);
  and _76283_ (_25531_, _25530_, _09771_);
  and _76284_ (_25532_, _25531_, _25529_);
  or _76285_ (_25533_, _09871_, \oc8051_golden_model_1.DPH [3]);
  nor _76286_ (_25534_, _09872_, _09771_);
  and _76287_ (_25535_, _25534_, _25533_);
  or _76288_ (_25536_, _25535_, _25532_);
  and _76289_ (_25537_, _25536_, _09755_);
  nor _76290_ (_25538_, _09755_, _03432_);
  or _76291_ (_25541_, _25538_, _07314_);
  or _76292_ (_25542_, _25541_, _25537_);
  and _76293_ (_25543_, _25542_, _25514_);
  or _76294_ (_25544_, _25543_, _03479_);
  and _76295_ (_25545_, _06717_, _05266_);
  or _76296_ (_25546_, _25508_, _06044_);
  or _76297_ (_25547_, _25546_, _25545_);
  and _76298_ (_25548_, _25547_, _03474_);
  and _76299_ (_25549_, _25548_, _25544_);
  nor _76300_ (_25550_, _12583_, _09848_);
  or _76301_ (_25552_, _25550_, _25508_);
  and _76302_ (_25553_, _25552_, _03221_);
  or _76303_ (_25554_, _25553_, _03437_);
  or _76304_ (_25555_, _25554_, _25549_);
  and _76305_ (_25556_, _05266_, _06217_);
  or _76306_ (_25557_, _25556_, _25508_);
  or _76307_ (_25558_, _25557_, _03438_);
  and _76308_ (_25559_, _25558_, _25555_);
  or _76309_ (_25560_, _25559_, _03636_);
  and _76310_ (_25561_, _12598_, _05266_);
  or _76311_ (_25563_, _25561_, _25508_);
  or _76312_ (_25564_, _25563_, _04499_);
  and _76313_ (_25565_, _25564_, _04501_);
  and _76314_ (_25566_, _25565_, _25560_);
  or _76315_ (_25567_, _25566_, _25511_);
  and _76316_ (_25568_, _25567_, _05769_);
  or _76317_ (_25569_, _25508_, _05521_);
  and _76318_ (_25570_, _25569_, _03754_);
  and _76319_ (_25571_, _25570_, _25557_);
  or _76320_ (_25572_, _25571_, _25568_);
  and _76321_ (_25574_, _25572_, _03753_);
  and _76322_ (_25575_, _25520_, _03752_);
  and _76323_ (_25576_, _25575_, _25569_);
  or _76324_ (_25577_, _25576_, _03758_);
  or _76325_ (_25578_, _25577_, _25574_);
  nor _76326_ (_25579_, _12597_, _09848_);
  or _76327_ (_25580_, _25508_, _03759_);
  or _76328_ (_25581_, _25580_, _25579_);
  and _76329_ (_25582_, _25581_, _04517_);
  and _76330_ (_25583_, _25582_, _25578_);
  nor _76331_ (_25585_, _12603_, _09848_);
  or _76332_ (_25586_, _25585_, _25508_);
  and _76333_ (_25587_, _25586_, _03760_);
  or _76334_ (_25588_, _25587_, _03790_);
  or _76335_ (_25589_, _25588_, _25583_);
  or _76336_ (_25590_, _25516_, _04192_);
  and _76337_ (_25591_, _25590_, _03521_);
  and _76338_ (_25592_, _25591_, _25589_);
  and _76339_ (_25593_, _12658_, _05266_);
  or _76340_ (_25594_, _25593_, _25508_);
  and _76341_ (_25596_, _25594_, _03520_);
  or _76342_ (_25597_, _25596_, _42967_);
  or _76343_ (_25598_, _25597_, _25592_);
  and _76344_ (_43321_, _25598_, _25506_);
  or _76345_ (_25599_, _42963_, \oc8051_golden_model_1.DPH [4]);
  and _76346_ (_25600_, _25599_, _41755_);
  not _76347_ (_25601_, \oc8051_golden_model_1.DPH [4]);
  nor _76348_ (_25602_, _05266_, _25601_);
  and _76349_ (_25603_, _12844_, _05266_);
  or _76350_ (_25604_, _25603_, _25602_);
  and _76351_ (_25606_, _25604_, _03769_);
  nor _76352_ (_25607_, _05712_, _09848_);
  or _76353_ (_25608_, _25607_, _25602_);
  or _76354_ (_25609_, _25608_, _06039_);
  nor _76355_ (_25610_, _12733_, _09848_);
  or _76356_ (_25611_, _25610_, _25602_);
  or _76357_ (_25612_, _25611_, _04444_);
  and _76358_ (_25613_, _05266_, \oc8051_golden_model_1.ACC [4]);
  or _76359_ (_25614_, _25613_, _25602_);
  and _76360_ (_25615_, _25614_, _04426_);
  nor _76361_ (_25617_, _04426_, _25601_);
  or _76362_ (_25618_, _25617_, _03570_);
  or _76363_ (_25619_, _25618_, _25615_);
  and _76364_ (_25620_, _25619_, _03983_);
  and _76365_ (_25621_, _25620_, _25612_);
  and _76366_ (_25622_, _25608_, _03568_);
  or _76367_ (_25623_, _25622_, _03575_);
  or _76368_ (_25624_, _25623_, _25621_);
  or _76369_ (_25625_, _25614_, _03583_);
  and _76370_ (_25626_, _25625_, _09771_);
  and _76371_ (_25628_, _25626_, _25624_);
  or _76372_ (_25629_, _09872_, \oc8051_golden_model_1.DPH [4]);
  nor _76373_ (_25630_, _09873_, _09771_);
  and _76374_ (_25631_, _25630_, _25629_);
  or _76375_ (_25632_, _25631_, _25628_);
  and _76376_ (_25633_, _25632_, _09755_);
  nor _76377_ (_25634_, _04249_, _09755_);
  or _76378_ (_25635_, _25634_, _07314_);
  or _76379_ (_25636_, _25635_, _25633_);
  and _76380_ (_25637_, _25636_, _25609_);
  or _76381_ (_25639_, _25637_, _03479_);
  and _76382_ (_25640_, _06722_, _05266_);
  or _76383_ (_25641_, _25602_, _06044_);
  or _76384_ (_25642_, _25641_, _25640_);
  and _76385_ (_25643_, _25642_, _03474_);
  and _76386_ (_25644_, _25643_, _25639_);
  nor _76387_ (_25645_, _12827_, _09848_);
  or _76388_ (_25646_, _25645_, _25602_);
  and _76389_ (_25647_, _25646_, _03221_);
  or _76390_ (_25648_, _25647_, _03437_);
  or _76391_ (_25650_, _25648_, _25644_);
  and _76392_ (_25651_, _06233_, _05266_);
  or _76393_ (_25652_, _25651_, _25602_);
  or _76394_ (_25653_, _25652_, _03438_);
  and _76395_ (_25654_, _25653_, _25650_);
  or _76396_ (_25655_, _25654_, _03636_);
  and _76397_ (_25656_, _12711_, _05266_);
  or _76398_ (_25657_, _25656_, _25602_);
  or _76399_ (_25658_, _25657_, _04499_);
  and _76400_ (_25659_, _25658_, _04501_);
  and _76401_ (_25661_, _25659_, _25655_);
  or _76402_ (_25662_, _25661_, _25606_);
  and _76403_ (_25663_, _25662_, _05769_);
  or _76404_ (_25664_, _25602_, _05761_);
  and _76405_ (_25665_, _25664_, _03754_);
  and _76406_ (_25666_, _25665_, _25652_);
  or _76407_ (_25667_, _25666_, _25663_);
  and _76408_ (_25668_, _25667_, _03753_);
  and _76409_ (_25669_, _25614_, _03752_);
  and _76410_ (_25670_, _25669_, _25664_);
  or _76411_ (_25672_, _25670_, _03758_);
  or _76412_ (_25673_, _25672_, _25668_);
  nor _76413_ (_25674_, _12710_, _09848_);
  or _76414_ (_25675_, _25602_, _03759_);
  or _76415_ (_25676_, _25675_, _25674_);
  and _76416_ (_25677_, _25676_, _04517_);
  and _76417_ (_25678_, _25677_, _25673_);
  nor _76418_ (_25679_, _12843_, _09848_);
  or _76419_ (_25680_, _25679_, _25602_);
  and _76420_ (_25681_, _25680_, _03760_);
  or _76421_ (_25683_, _25681_, _03790_);
  or _76422_ (_25684_, _25683_, _25678_);
  or _76423_ (_25685_, _25611_, _04192_);
  and _76424_ (_25686_, _25685_, _03521_);
  and _76425_ (_25687_, _25686_, _25684_);
  and _76426_ (_25688_, _12893_, _05266_);
  or _76427_ (_25689_, _25688_, _25602_);
  and _76428_ (_25690_, _25689_, _03520_);
  or _76429_ (_25691_, _25690_, _42967_);
  or _76430_ (_25692_, _25691_, _25687_);
  and _76431_ (_43322_, _25692_, _25600_);
  or _76432_ (_25694_, _42963_, \oc8051_golden_model_1.DPH [5]);
  and _76433_ (_25695_, _25694_, _41755_);
  and _76434_ (_25696_, _09848_, \oc8051_golden_model_1.DPH [5]);
  and _76435_ (_25697_, _13042_, _05266_);
  or _76436_ (_25698_, _25697_, _25696_);
  and _76437_ (_25699_, _25698_, _03769_);
  nor _76438_ (_25700_, _05422_, _09848_);
  or _76439_ (_25701_, _25700_, _25696_);
  or _76440_ (_25702_, _25701_, _06039_);
  nor _76441_ (_25704_, _12930_, _09848_);
  or _76442_ (_25705_, _25704_, _25696_);
  or _76443_ (_25706_, _25705_, _04444_);
  and _76444_ (_25707_, _05266_, \oc8051_golden_model_1.ACC [5]);
  or _76445_ (_25708_, _25707_, _25696_);
  and _76446_ (_25709_, _25708_, _04426_);
  and _76447_ (_25710_, _04427_, \oc8051_golden_model_1.DPH [5]);
  or _76448_ (_25711_, _25710_, _03570_);
  or _76449_ (_25712_, _25711_, _25709_);
  and _76450_ (_25713_, _25712_, _03983_);
  and _76451_ (_25715_, _25713_, _25706_);
  and _76452_ (_25716_, _25701_, _03568_);
  or _76453_ (_25717_, _25716_, _03575_);
  or _76454_ (_25718_, _25717_, _25715_);
  or _76455_ (_25719_, _25708_, _03583_);
  and _76456_ (_25720_, _25719_, _09771_);
  and _76457_ (_25721_, _25720_, _25718_);
  or _76458_ (_25722_, _09873_, \oc8051_golden_model_1.DPH [5]);
  nor _76459_ (_25723_, _09874_, _09771_);
  and _76460_ (_25724_, _25723_, _25722_);
  or _76461_ (_25725_, _25724_, _25721_);
  and _76462_ (_25726_, _25725_, _09755_);
  nor _76463_ (_25727_, _03834_, _09755_);
  or _76464_ (_25728_, _25727_, _07314_);
  or _76465_ (_25729_, _25728_, _25726_);
  and _76466_ (_25730_, _25729_, _25702_);
  or _76467_ (_25731_, _25730_, _03479_);
  and _76468_ (_25732_, _06721_, _05266_);
  or _76469_ (_25733_, _25696_, _06044_);
  or _76470_ (_25734_, _25733_, _25732_);
  and _76471_ (_25737_, _25734_, _03474_);
  and _76472_ (_25738_, _25737_, _25731_);
  nor _76473_ (_25739_, _13021_, _09848_);
  or _76474_ (_25740_, _25739_, _25696_);
  and _76475_ (_25741_, _25740_, _03221_);
  or _76476_ (_25742_, _25741_, _03437_);
  or _76477_ (_25743_, _25742_, _25738_);
  and _76478_ (_25744_, _06211_, _05266_);
  or _76479_ (_25745_, _25744_, _25696_);
  or _76480_ (_25746_, _25745_, _03438_);
  and _76481_ (_25748_, _25746_, _25743_);
  or _76482_ (_25749_, _25748_, _03636_);
  and _76483_ (_25750_, _13036_, _05266_);
  or _76484_ (_25751_, _25750_, _25696_);
  or _76485_ (_25752_, _25751_, _04499_);
  and _76486_ (_25753_, _25752_, _04501_);
  and _76487_ (_25754_, _25753_, _25749_);
  or _76488_ (_25755_, _25754_, _25699_);
  and _76489_ (_25756_, _25755_, _05769_);
  or _76490_ (_25757_, _25696_, _05472_);
  and _76491_ (_25759_, _25757_, _03754_);
  and _76492_ (_25760_, _25759_, _25745_);
  or _76493_ (_25761_, _25760_, _25756_);
  and _76494_ (_25762_, _25761_, _03753_);
  and _76495_ (_25763_, _25708_, _03752_);
  and _76496_ (_25764_, _25763_, _25757_);
  or _76497_ (_25765_, _25764_, _03758_);
  or _76498_ (_25766_, _25765_, _25762_);
  nor _76499_ (_25767_, _13035_, _09848_);
  or _76500_ (_25768_, _25696_, _03759_);
  or _76501_ (_25770_, _25768_, _25767_);
  and _76502_ (_25771_, _25770_, _04517_);
  and _76503_ (_25772_, _25771_, _25766_);
  nor _76504_ (_25773_, _13041_, _09848_);
  or _76505_ (_25774_, _25773_, _25696_);
  and _76506_ (_25775_, _25774_, _03760_);
  or _76507_ (_25776_, _25775_, _03790_);
  or _76508_ (_25777_, _25776_, _25772_);
  or _76509_ (_25778_, _25705_, _04192_);
  and _76510_ (_25779_, _25778_, _03521_);
  and _76511_ (_25781_, _25779_, _25777_);
  and _76512_ (_25782_, _13097_, _05266_);
  or _76513_ (_25783_, _25782_, _25696_);
  and _76514_ (_25784_, _25783_, _03520_);
  or _76515_ (_25785_, _25784_, _42967_);
  or _76516_ (_25786_, _25785_, _25781_);
  and _76517_ (_43323_, _25786_, _25695_);
  or _76518_ (_25787_, _42963_, \oc8051_golden_model_1.DPH [6]);
  and _76519_ (_25788_, _25787_, _41755_);
  not _76520_ (_25789_, \oc8051_golden_model_1.DPH [6]);
  nor _76521_ (_25791_, _05266_, _25789_);
  and _76522_ (_25792_, _13259_, _05266_);
  or _76523_ (_25793_, _25792_, _25791_);
  and _76524_ (_25794_, _25793_, _03769_);
  nor _76525_ (_25795_, _05327_, _09848_);
  or _76526_ (_25796_, _25795_, _25791_);
  or _76527_ (_25797_, _25796_, _06039_);
  nor _76528_ (_25798_, _13122_, _09848_);
  or _76529_ (_25799_, _25798_, _25791_);
  or _76530_ (_25800_, _25799_, _04444_);
  and _76531_ (_25802_, _05266_, \oc8051_golden_model_1.ACC [6]);
  or _76532_ (_25803_, _25802_, _25791_);
  and _76533_ (_25804_, _25803_, _04426_);
  nor _76534_ (_25805_, _04426_, _25789_);
  or _76535_ (_25806_, _25805_, _03570_);
  or _76536_ (_25807_, _25806_, _25804_);
  and _76537_ (_25808_, _25807_, _03983_);
  and _76538_ (_25809_, _25808_, _25800_);
  and _76539_ (_25810_, _25796_, _03568_);
  or _76540_ (_25811_, _25810_, _03575_);
  or _76541_ (_25813_, _25811_, _25809_);
  or _76542_ (_25814_, _25803_, _03583_);
  and _76543_ (_25815_, _25814_, _09771_);
  and _76544_ (_25816_, _25815_, _25813_);
  or _76545_ (_25817_, _09874_, \oc8051_golden_model_1.DPH [6]);
  and _76546_ (_25818_, _09875_, _09770_);
  and _76547_ (_25819_, _25818_, _25817_);
  or _76548_ (_25820_, _25819_, _25816_);
  and _76549_ (_25821_, _25820_, _09755_);
  nor _76550_ (_25822_, _09755_, _03561_);
  or _76551_ (_25824_, _25822_, _07314_);
  or _76552_ (_25825_, _25824_, _25821_);
  and _76553_ (_25826_, _25825_, _25797_);
  or _76554_ (_25827_, _25826_, _03479_);
  and _76555_ (_25828_, _06713_, _05266_);
  or _76556_ (_25829_, _25791_, _06044_);
  or _76557_ (_25830_, _25829_, _25828_);
  and _76558_ (_25831_, _25830_, _03474_);
  and _76559_ (_25832_, _25831_, _25827_);
  nor _76560_ (_25833_, _13237_, _09848_);
  or _76561_ (_25835_, _25833_, _25791_);
  and _76562_ (_25836_, _25835_, _03221_);
  or _76563_ (_25837_, _25836_, _03437_);
  or _76564_ (_25838_, _25837_, _25832_);
  and _76565_ (_25839_, _13244_, _05266_);
  or _76566_ (_25840_, _25839_, _25791_);
  or _76567_ (_25841_, _25840_, _03438_);
  and _76568_ (_25842_, _25841_, _25838_);
  or _76569_ (_25843_, _25842_, _03636_);
  and _76570_ (_25844_, _13253_, _05266_);
  or _76571_ (_25846_, _25844_, _25791_);
  or _76572_ (_25847_, _25846_, _04499_);
  and _76573_ (_25848_, _25847_, _04501_);
  and _76574_ (_25849_, _25848_, _25843_);
  or _76575_ (_25850_, _25849_, _25794_);
  and _76576_ (_25851_, _25850_, _05769_);
  or _76577_ (_25852_, _25791_, _05377_);
  and _76578_ (_25853_, _25852_, _03754_);
  and _76579_ (_25854_, _25853_, _25840_);
  or _76580_ (_25855_, _25854_, _25851_);
  and _76581_ (_25857_, _25855_, _03753_);
  and _76582_ (_25858_, _25803_, _03752_);
  and _76583_ (_25859_, _25858_, _25852_);
  or _76584_ (_25860_, _25859_, _03758_);
  or _76585_ (_25861_, _25860_, _25857_);
  nor _76586_ (_25862_, _13251_, _09848_);
  or _76587_ (_25863_, _25791_, _03759_);
  or _76588_ (_25864_, _25863_, _25862_);
  and _76589_ (_25865_, _25864_, _04517_);
  and _76590_ (_25866_, _25865_, _25861_);
  nor _76591_ (_25868_, _13258_, _09848_);
  or _76592_ (_25869_, _25868_, _25791_);
  and _76593_ (_25870_, _25869_, _03760_);
  or _76594_ (_25871_, _25870_, _03790_);
  or _76595_ (_25872_, _25871_, _25866_);
  or _76596_ (_25873_, _25799_, _04192_);
  and _76597_ (_25874_, _25873_, _03521_);
  and _76598_ (_25875_, _25874_, _25872_);
  and _76599_ (_25876_, _13312_, _05266_);
  or _76600_ (_25877_, _25876_, _25791_);
  and _76601_ (_25879_, _25877_, _03520_);
  or _76602_ (_25880_, _25879_, _42967_);
  or _76603_ (_25881_, _25880_, _25875_);
  and _76604_ (_43324_, _25881_, _25788_);
  nor _76605_ (_25882_, _03645_, _03166_);
  not _76606_ (_25883_, _25882_);
  and _76607_ (_25884_, _25883_, _04109_);
  and _76608_ (_25885_, _10821_, _10828_);
  nor _76609_ (_25886_, _25885_, _02887_);
  not _76610_ (_25887_, _03172_);
  and _76611_ (_25889_, _09949_, _10803_);
  nor _76612_ (_25890_, _25889_, _02887_);
  not _76613_ (_25891_, _03192_);
  nor _76614_ (_25892_, _10545_, _04504_);
  nor _76615_ (_25893_, _25892_, _02887_);
  not _76616_ (_25894_, _03194_);
  and _76617_ (_25895_, _10520_, _04499_);
  nor _76618_ (_25896_, _25895_, _02887_);
  not _76619_ (_25897_, _10472_);
  and _76620_ (_25898_, _03437_, _02887_);
  nor _76621_ (_25900_, _04109_, _03213_);
  and _76622_ (_25901_, _10316_, _10307_);
  nor _76623_ (_25902_, _25901_, _02887_);
  and _76624_ (_25903_, _04109_, _03923_);
  nor _76625_ (_25904_, _10290_, _02887_);
  and _76626_ (_25905_, _10278_, _10275_);
  nor _76627_ (_25906_, _25905_, _02887_);
  and _76628_ (_25907_, _25905_, _02887_);
  nor _76629_ (_25908_, _25907_, _25906_);
  and _76630_ (_25909_, _10290_, _04762_);
  not _76631_ (_25911_, _25909_);
  nor _76632_ (_25912_, _25911_, _25908_);
  nor _76633_ (_25913_, _25912_, _25904_);
  not _76634_ (_25914_, _25913_);
  nor _76635_ (_25915_, _25914_, _25903_);
  nor _76636_ (_25916_, _25915_, _05833_);
  and _76637_ (_25917_, _10269_, \oc8051_golden_model_1.PC [0]);
  and _76638_ (_25918_, _03471_, _02887_);
  nor _76639_ (_25919_, _25918_, _10022_);
  and _76640_ (_25920_, _25919_, _10271_);
  or _76641_ (_25922_, _25920_, _25917_);
  nor _76642_ (_25923_, _25922_, _05831_);
  nor _76643_ (_25924_, _25923_, _25916_);
  nor _76644_ (_25925_, _25924_, _04438_);
  and _76645_ (_25926_, _04438_, \oc8051_golden_model_1.PC [0]);
  nor _76646_ (_25927_, _25926_, _25925_);
  and _76647_ (_25928_, _25927_, _04444_);
  not _76648_ (_25929_, _25928_);
  and _76649_ (_25930_, _04109_, \oc8051_golden_model_1.PC [0]);
  nor _76650_ (_25931_, _25930_, _10192_);
  nor _76651_ (_25933_, _25931_, _10261_);
  and _76652_ (_25934_, _05664_, _05940_);
  and _76653_ (_25935_, _05617_, _05520_);
  and _76654_ (_25936_, _25935_, _10260_);
  nand _76655_ (_25937_, _25936_, _25934_);
  nor _76656_ (_25938_, _25937_, _02887_);
  or _76657_ (_25939_, _25938_, _04444_);
  or _76658_ (_25940_, _25939_, _25933_);
  and _76659_ (_25941_, _25940_, _10255_);
  and _76660_ (_25942_, _25941_, _25929_);
  nor _76661_ (_25944_, _10255_, _02887_);
  nor _76662_ (_25945_, _25944_, _04746_);
  not _76663_ (_25946_, _25945_);
  nor _76664_ (_25947_, _25946_, _25942_);
  nor _76665_ (_25948_, _04109_, _03203_);
  not _76666_ (_25949_, _25901_);
  nor _76667_ (_25950_, _25949_, _25948_);
  not _76668_ (_25951_, _25950_);
  nor _76669_ (_25952_, _25951_, _25947_);
  or _76670_ (_25953_, _25952_, _10249_);
  nor _76671_ (_25955_, _25953_, _25902_);
  nor _76672_ (_25956_, _04109_, _03206_);
  nor _76673_ (_25957_, _25956_, _10326_);
  not _76674_ (_25958_, _25957_);
  nor _76675_ (_25959_, _25958_, _25955_);
  and _76676_ (_25960_, _10360_, _02887_);
  not _76677_ (_25961_, _25931_);
  nor _76678_ (_25962_, _25961_, _10360_);
  or _76679_ (_25963_, _25962_, _25960_);
  nor _76680_ (_25964_, _25963_, _10325_);
  or _76681_ (_25966_, _25964_, _03657_);
  nor _76682_ (_25967_, _25966_, _25959_);
  nand _76683_ (_25968_, _10116_, \oc8051_golden_model_1.PC [0]);
  or _76684_ (_25969_, _25931_, _10116_);
  and _76685_ (_25970_, _25969_, _03657_);
  and _76686_ (_25971_, _25970_, _25968_);
  or _76687_ (_25972_, _25971_, _25967_);
  and _76688_ (_25973_, _25972_, _03998_);
  and _76689_ (_25974_, _10382_, _02887_);
  nor _76690_ (_25975_, _25961_, _10382_);
  nor _76691_ (_25977_, _25975_, _25974_);
  nor _76692_ (_25978_, _25977_, _03998_);
  nor _76693_ (_25979_, _25978_, _25973_);
  nor _76694_ (_25980_, _25979_, _03638_);
  and _76695_ (_25981_, _10398_, _02887_);
  nor _76696_ (_25982_, _25961_, _10398_);
  or _76697_ (_25983_, _25982_, _25981_);
  and _76698_ (_25984_, _25983_, _03638_);
  or _76699_ (_25985_, _25984_, _25980_);
  and _76700_ (_25986_, _25985_, _10084_);
  and _76701_ (_25988_, _10083_, _02887_);
  or _76702_ (_25989_, _25988_, _25986_);
  and _76703_ (_25990_, _25989_, _03200_);
  not _76704_ (_25991_, _10415_);
  nor _76705_ (_25992_, _04109_, _03200_);
  nor _76706_ (_25993_, _25992_, _25991_);
  not _76707_ (_25994_, _25993_);
  nor _76708_ (_25995_, _25994_, _25990_);
  nor _76709_ (_25996_, _10415_, _02887_);
  nor _76710_ (_25997_, _25996_, _10420_);
  not _76711_ (_25999_, _25997_);
  nor _76712_ (_26000_, _25999_, _25995_);
  and _76713_ (_26001_, _10426_, _03254_);
  not _76714_ (_26002_, _26001_);
  or _76715_ (_26003_, _26002_, _26000_);
  nor _76716_ (_26004_, _26003_, _25900_);
  nor _76717_ (_26005_, _26001_, _02887_);
  nor _76718_ (_26006_, _26005_, _03223_);
  not _76719_ (_26007_, _26006_);
  nor _76720_ (_26008_, _26007_, _26004_);
  nor _76721_ (_26010_, _04109_, _04853_);
  nor _76722_ (_26011_, _03632_, _03221_);
  and _76723_ (_26012_, _26011_, _10081_);
  not _76724_ (_26013_, _26012_);
  nor _76725_ (_26014_, _26013_, _26010_);
  not _76726_ (_26015_, _26014_);
  nor _76727_ (_26016_, _26015_, _26008_);
  nor _76728_ (_26017_, _26012_, _02887_);
  nor _76729_ (_26018_, _26017_, _03187_);
  not _76730_ (_26019_, _26018_);
  nor _76731_ (_26021_, _26019_, _26016_);
  not _76732_ (_26022_, _03187_);
  nor _76733_ (_26023_, _04109_, _26022_);
  or _76734_ (_26024_, _26023_, _10458_);
  nor _76735_ (_26025_, _26024_, _26021_);
  nor _76736_ (_26026_, _25919_, _10459_);
  nor _76737_ (_26027_, _26026_, _26025_);
  and _76738_ (_26028_, _26027_, _03438_);
  or _76739_ (_26029_, _26028_, _25898_);
  and _76740_ (_26030_, _26029_, _25897_);
  and _76741_ (_26032_, _10472_, _03313_);
  or _76742_ (_26033_, _26032_, _26030_);
  and _76743_ (_26034_, _26033_, _11376_);
  nor _76744_ (_26035_, _04109_, _11376_);
  or _76745_ (_26036_, _26035_, _26034_);
  and _76746_ (_26037_, _26036_, _10515_);
  not _76747_ (_26038_, _25895_);
  and _76748_ (_26039_, _08698_, \oc8051_golden_model_1.PC [0]);
  and _76749_ (_26040_, _25919_, _10077_);
  or _76750_ (_26041_, _26040_, _26039_);
  and _76751_ (_26043_, _26041_, _10076_);
  nor _76752_ (_26044_, _26043_, _26038_);
  not _76753_ (_26045_, _26044_);
  nor _76754_ (_26046_, _26045_, _26037_);
  nor _76755_ (_26047_, _26046_, _25896_);
  and _76756_ (_26048_, _26047_, _25894_);
  nor _76757_ (_26049_, _04109_, _25894_);
  or _76758_ (_26050_, _26049_, _26048_);
  and _76759_ (_26051_, _26050_, _10535_);
  not _76760_ (_26052_, _25892_);
  nor _76761_ (_26054_, _25919_, _10077_);
  nor _76762_ (_26055_, _08698_, \oc8051_golden_model_1.PC [0]);
  nor _76763_ (_26056_, _26055_, _10535_);
  not _76764_ (_26057_, _26056_);
  nor _76765_ (_26058_, _26057_, _26054_);
  nor _76766_ (_26059_, _26058_, _26052_);
  not _76767_ (_26060_, _26059_);
  nor _76768_ (_26061_, _26060_, _26051_);
  nor _76769_ (_26062_, _26061_, _25893_);
  and _76770_ (_26063_, _26062_, _25891_);
  nor _76771_ (_26065_, _04109_, _25891_);
  or _76772_ (_26066_, _26065_, _26063_);
  and _76773_ (_26067_, _26066_, _09959_);
  and _76774_ (_26068_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and _76775_ (_26069_, _25919_, _07888_);
  or _76776_ (_26070_, _26069_, _26068_);
  and _76777_ (_26071_, _26070_, _09958_);
  and _76778_ (_26072_, _09956_, _03759_);
  not _76779_ (_26073_, _26072_);
  nor _76780_ (_26074_, _26073_, _26071_);
  not _76781_ (_26075_, _26074_);
  nor _76782_ (_26076_, _26075_, _26067_);
  nor _76783_ (_26077_, _10576_, _03183_);
  not _76784_ (_26078_, _26077_);
  nor _76785_ (_26079_, _26072_, _02887_);
  or _76786_ (_26080_, _26079_, _26078_);
  nor _76787_ (_26081_, _26080_, _26076_);
  not _76788_ (_26082_, _03183_);
  nor _76789_ (_26083_, _04109_, _26082_);
  nor _76790_ (_26084_, _08328_, _02887_);
  and _76791_ (_26087_, _08328_, _02887_);
  nor _76792_ (_26088_, _26087_, _26084_);
  nor _76793_ (_26089_, _26088_, _10577_);
  and _76794_ (_26090_, _09951_, _08556_);
  not _76795_ (_26091_, _26090_);
  or _76796_ (_26092_, _26091_, _26089_);
  nor _76797_ (_26093_, _26092_, _26083_);
  not _76798_ (_26094_, _26093_);
  nor _76799_ (_26095_, _26094_, _26081_);
  nor _76800_ (_26096_, _26090_, _02887_);
  nor _76801_ (_26098_, _26096_, _03775_);
  not _76802_ (_26099_, _26098_);
  nor _76803_ (_26100_, _26099_, _26095_);
  and _76804_ (_26101_, _06715_, _03775_);
  or _76805_ (_26102_, _26101_, _26100_);
  and _76806_ (_26103_, _26102_, _06328_);
  nor _76807_ (_26104_, _04109_, _06328_);
  or _76808_ (_26105_, _26104_, _26103_);
  and _76809_ (_26106_, _26105_, _10599_);
  and _76810_ (_26107_, _25961_, _10794_);
  nor _76811_ (_26109_, _10794_, _02887_);
  or _76812_ (_26110_, _26109_, _10599_);
  or _76813_ (_26111_, _26110_, _26107_);
  and _76814_ (_26112_, _26111_, _25889_);
  not _76815_ (_26113_, _26112_);
  nor _76816_ (_26114_, _26113_, _26106_);
  nor _76817_ (_26115_, _26114_, _25890_);
  and _76818_ (_26116_, _26115_, _03523_);
  and _76819_ (_26117_, _06715_, _03522_);
  or _76820_ (_26118_, _26117_, _26116_);
  and _76821_ (_26120_, _26118_, _25887_);
  nor _76822_ (_26121_, _04109_, _25887_);
  nor _76823_ (_26122_, _26121_, _26120_);
  nor _76824_ (_26123_, _26122_, _03628_);
  not _76825_ (_26124_, _25885_);
  and _76826_ (_26125_, _10794_, \oc8051_golden_model_1.PC [0]);
  nor _76827_ (_26126_, _25931_, _10794_);
  nor _76828_ (_26127_, _26126_, _26125_);
  and _76829_ (_26128_, _26127_, _03628_);
  nor _76830_ (_26129_, _26128_, _26124_);
  not _76831_ (_26131_, _26129_);
  nor _76832_ (_26132_, _26131_, _26123_);
  nor _76833_ (_26133_, _26132_, _25886_);
  nor _76834_ (_26134_, _26133_, _04947_);
  and _76835_ (_26135_, _04947_, _04109_);
  nor _76836_ (_26136_, _26135_, _03151_);
  not _76837_ (_26137_, _26136_);
  nor _76838_ (_26138_, _26137_, _26134_);
  and _76839_ (_26139_, _26127_, _03151_);
  and _76840_ (_26140_, _10844_, _10851_);
  not _76841_ (_26142_, _26140_);
  nor _76842_ (_26143_, _26142_, _26139_);
  not _76843_ (_26144_, _26143_);
  nor _76844_ (_26145_, _26144_, _26138_);
  nor _76845_ (_26146_, _26140_, _02887_);
  nor _76846_ (_26147_, _26146_, _26145_);
  nor _76847_ (_26148_, _26147_, _25883_);
  or _76848_ (_26149_, _26148_, _10862_);
  nor _76849_ (_26150_, _26149_, _25884_);
  and _76850_ (_26151_, _10862_, _02887_);
  nor _76851_ (_26153_, _26151_, _26150_);
  nand _76852_ (_26154_, _26153_, _42963_);
  or _76853_ (_26155_, _42963_, \oc8051_golden_model_1.PC [0]);
  and _76854_ (_26156_, _26155_, _41755_);
  and _76855_ (_43327_, _26156_, _26154_);
  and _76856_ (_26157_, _25883_, _04317_);
  and _76857_ (_26158_, _03520_, _02860_);
  and _76858_ (_26159_, _03661_, _03165_);
  nor _76859_ (_26160_, _26159_, _04766_);
  and _76860_ (_26161_, _03790_, _02860_);
  and _76861_ (_26163_, _13062_, _03234_);
  nor _76862_ (_26164_, _09949_, _10190_);
  nor _76863_ (_26165_, _09953_, _10190_);
  and _76864_ (_26166_, _03752_, \oc8051_golden_model_1.PC [1]);
  nor _76865_ (_26167_, _10520_, _10190_);
  nor _76866_ (_26168_, _10426_, _10190_);
  nor _76867_ (_26169_, _04317_, _03203_);
  nor _76868_ (_26170_, _10194_, _10192_);
  nor _76869_ (_26171_, _26170_, _10195_);
  or _76870_ (_26172_, _26171_, _10261_);
  and _76871_ (_26174_, _26172_, _03570_);
  nand _76872_ (_26175_, _10261_, _10190_);
  and _76873_ (_26176_, _26175_, _26174_);
  nand _76874_ (_26177_, _04317_, _03923_);
  nor _76875_ (_26178_, _04426_, \oc8051_golden_model_1.PC [0]);
  not _76876_ (_26179_, _03922_);
  and _76877_ (_26180_, _10278_, _26179_);
  nor _76878_ (_26181_, _26180_, _26178_);
  and _76879_ (_26182_, _26181_, \oc8051_golden_model_1.PC [1]);
  nor _76880_ (_26183_, _26181_, \oc8051_golden_model_1.PC [1]);
  nor _76881_ (_26184_, _26183_, _26182_);
  or _76882_ (_26185_, _26184_, _25911_);
  nor _76883_ (_26186_, _10290_, _10190_);
  nor _76884_ (_26187_, _26186_, _05833_);
  and _76885_ (_26188_, _26187_, _26185_);
  and _76886_ (_26189_, _26188_, _26177_);
  not _76887_ (_26190_, _26189_);
  nor _76888_ (_26191_, _10024_, _10022_);
  nor _76889_ (_26192_, _26191_, _10025_);
  nand _76890_ (_26193_, _26192_, _10271_);
  or _76891_ (_26196_, _10271_, \oc8051_golden_model_1.PC [1]);
  nand _76892_ (_26197_, _26196_, _26193_);
  nand _76893_ (_26198_, _26197_, _05833_);
  and _76894_ (_26199_, _26198_, _26190_);
  nor _76895_ (_26200_, _26199_, _10297_);
  or _76896_ (_26201_, _26200_, _26176_);
  and _76897_ (_26202_, _26201_, _10255_);
  nor _76898_ (_26203_, _10303_, _03234_);
  or _76899_ (_26204_, _26203_, _03516_);
  or _76900_ (_26205_, _26204_, _26202_);
  and _76901_ (_26207_, _03516_, \oc8051_golden_model_1.PC [1]);
  nor _76902_ (_26208_, _26207_, _04746_);
  and _76903_ (_26209_, _26208_, _26205_);
  or _76904_ (_26210_, _26209_, _26169_);
  nand _76905_ (_26211_, _26210_, _03983_);
  not _76906_ (_26212_, _10307_);
  and _76907_ (_26213_, _03568_, _02860_);
  nor _76908_ (_26214_, _26213_, _26212_);
  nand _76909_ (_26215_, _26214_, _26211_);
  nor _76910_ (_26216_, _10307_, _10190_);
  nor _76911_ (_26218_, _26216_, _03575_);
  nand _76912_ (_26219_, _26218_, _26215_);
  not _76913_ (_26220_, _10316_);
  and _76914_ (_26221_, _03575_, _02860_);
  nor _76915_ (_26222_, _26221_, _26220_);
  nand _76916_ (_26223_, _26222_, _26219_);
  nor _76917_ (_26224_, _10316_, _10190_);
  nor _76918_ (_26225_, _26224_, _03512_);
  nand _76919_ (_26226_, _26225_, _26223_);
  and _76920_ (_26227_, _03512_, _02860_);
  nor _76921_ (_26229_, _26227_, _10249_);
  nand _76922_ (_26230_, _26229_, _26226_);
  and _76923_ (_26231_, _04317_, _10249_);
  nor _76924_ (_26232_, _26231_, _03511_);
  nand _76925_ (_26233_, _26232_, _26230_);
  and _76926_ (_26234_, _03511_, _02860_);
  nor _76927_ (_26235_, _26234_, _10326_);
  nand _76928_ (_26236_, _26235_, _26233_);
  and _76929_ (_26237_, _10360_, _03234_);
  not _76930_ (_26238_, _26171_);
  nor _76931_ (_26240_, _26238_, _10360_);
  or _76932_ (_26241_, _26240_, _26237_);
  nor _76933_ (_26242_, _26241_, _10325_);
  nor _76934_ (_26243_, _26242_, _03657_);
  nand _76935_ (_26244_, _26243_, _26236_);
  or _76936_ (_26245_, _26238_, _10116_);
  nand _76937_ (_26246_, _10116_, _03234_);
  and _76938_ (_26247_, _26246_, _26245_);
  or _76939_ (_26248_, _26247_, _10328_);
  and _76940_ (_26249_, _26248_, _03998_);
  and _76941_ (_26251_, _26249_, _26244_);
  nor _76942_ (_26252_, _26238_, _10382_);
  and _76943_ (_26253_, _10382_, _03234_);
  or _76944_ (_26254_, _26253_, _03998_);
  nor _76945_ (_26255_, _26254_, _26252_);
  or _76946_ (_26256_, _26255_, _03638_);
  or _76947_ (_26257_, _26256_, _26251_);
  nor _76948_ (_26258_, _26171_, _10398_);
  and _76949_ (_26259_, _10398_, _10190_);
  or _76950_ (_26260_, _26259_, _10085_);
  or _76951_ (_26262_, _26260_, _26258_);
  and _76952_ (_26263_, _26262_, _10084_);
  and _76953_ (_26264_, _26263_, _26257_);
  and _76954_ (_26265_, _10083_, _03234_);
  or _76955_ (_26266_, _26265_, _26264_);
  nand _76956_ (_26267_, _26266_, _03506_);
  and _76957_ (_26268_, _03505_, \oc8051_golden_model_1.PC [1]);
  nor _76958_ (_26269_, _26268_, _04743_);
  nand _76959_ (_26270_, _26269_, _26267_);
  nor _76960_ (_26271_, _04317_, _03200_);
  and _76961_ (_26273_, _03483_, _03596_);
  not _76962_ (_26274_, _26273_);
  and _76963_ (_26275_, _03601_, _26274_);
  and _76964_ (_26276_, _03633_, _03596_);
  nor _76965_ (_26277_, _26276_, _03592_);
  and _76966_ (_26278_, _03655_, _03596_);
  nor _76967_ (_26279_, _04478_, _26278_);
  and _76968_ (_26280_, _26279_, _26277_);
  and _76969_ (_26281_, _26280_, _26275_);
  not _76970_ (_26282_, _26281_);
  nor _76971_ (_26284_, _26282_, _26271_);
  nand _76972_ (_26285_, _26284_, _26270_);
  nor _76973_ (_26286_, _26281_, _02860_);
  nor _76974_ (_26287_, _26286_, _10412_);
  nand _76975_ (_26288_, _26287_, _26285_);
  and _76976_ (_26289_, _10414_, _03234_);
  or _76977_ (_26290_, _26289_, _10415_);
  nand _76978_ (_26291_, _26290_, _26288_);
  nor _76979_ (_26292_, _10414_, _10190_);
  nor _76980_ (_26293_, _26292_, _03607_);
  nand _76981_ (_26295_, _26293_, _26291_);
  and _76982_ (_26296_, _03607_, _02860_);
  nor _76983_ (_26297_, _26296_, _10420_);
  nand _76984_ (_26298_, _26297_, _26295_);
  and _76985_ (_26299_, _04317_, _10420_);
  nor _76986_ (_26300_, _26299_, _03606_);
  nand _76987_ (_26301_, _26300_, _26298_);
  not _76988_ (_26302_, _10426_);
  and _76989_ (_26303_, _03606_, _02860_);
  nor _76990_ (_26304_, _26303_, _26302_);
  and _76991_ (_26306_, _26304_, _26301_);
  or _76992_ (_26307_, _26306_, _26168_);
  nand _76993_ (_26308_, _26307_, _10430_);
  nor _76994_ (_26309_, _10430_, _02860_);
  nor _76995_ (_26310_, _26309_, _03311_);
  and _76996_ (_26311_, _26310_, _26308_);
  nor _76997_ (_26312_, _03254_, _03234_);
  or _76998_ (_26313_, _26312_, _03499_);
  nor _76999_ (_26314_, _26313_, _26311_);
  and _77000_ (_26315_, _03499_, \oc8051_golden_model_1.PC [1]);
  or _77001_ (_26317_, _26315_, _26314_);
  nand _77002_ (_26318_, _26317_, _04853_);
  and _77003_ (_26319_, _04317_, _03223_);
  nor _77004_ (_26320_, _26319_, _03632_);
  nand _77005_ (_26321_, _26320_, _26318_);
  not _77006_ (_26322_, _03493_);
  and _77007_ (_26323_, _03632_, _03234_);
  nor _77008_ (_26324_, _26323_, _26322_);
  nand _77009_ (_26325_, _26324_, _26321_);
  nor _77010_ (_26326_, _03493_, _02860_);
  nor _77011_ (_26328_, _26326_, _03221_);
  nand _77012_ (_26329_, _26328_, _26325_);
  not _77013_ (_26330_, _10081_);
  and _77014_ (_26331_, _03234_, _03221_);
  nor _77015_ (_26332_, _26331_, _26330_);
  nand _77016_ (_26333_, _26332_, _26329_);
  nor _77017_ (_26334_, _10081_, _10190_);
  nor _77018_ (_26335_, _26334_, _03745_);
  nand _77019_ (_26336_, _26335_, _26333_);
  and _77020_ (_26337_, _03745_, _02860_);
  nor _77021_ (_26339_, _26337_, _03187_);
  nand _77022_ (_26340_, _26339_, _26336_);
  and _77023_ (_26341_, _04317_, _03187_);
  nor _77024_ (_26342_, _26341_, _10458_);
  nand _77025_ (_26343_, _26342_, _26340_);
  and _77026_ (_26344_, _26192_, _10458_);
  nor _77027_ (_26345_, _26344_, _06055_);
  nand _77028_ (_26346_, _26345_, _26343_);
  nor _77029_ (_26347_, _05775_, _02860_);
  nor _77030_ (_26348_, _26347_, _03437_);
  nand _77031_ (_26350_, _26348_, _26346_);
  and _77032_ (_26351_, _03437_, _03234_);
  nor _77033_ (_26352_, _26351_, _08385_);
  and _77034_ (_26353_, _26352_, _26350_);
  and _77035_ (_26354_, _08385_, \oc8051_golden_model_1.PC [1]);
  or _77036_ (_26355_, _26354_, _26353_);
  nand _77037_ (_26356_, _26355_, _25897_);
  nor _77038_ (_26357_, _25897_, _03332_);
  nor _77039_ (_26358_, _26357_, _03744_);
  nand _77040_ (_26359_, _26358_, _26356_);
  and _77041_ (_26361_, _03744_, _02860_);
  nor _77042_ (_26362_, _26361_, _03189_);
  nand _77043_ (_26363_, _26362_, _26359_);
  and _77044_ (_26364_, _04317_, _03189_);
  nor _77045_ (_26365_, _26364_, _10076_);
  nand _77046_ (_26366_, _26365_, _26363_);
  nor _77047_ (_26367_, _26192_, _08698_);
  nand _77048_ (_26368_, _08698_, \oc8051_golden_model_1.PC [1]);
  nand _77049_ (_26369_, _26368_, _10076_);
  or _77050_ (_26370_, _26369_, _26367_);
  and _77051_ (_26372_, _26370_, _10520_);
  and _77052_ (_26373_, _26372_, _26366_);
  or _77053_ (_26374_, _26373_, _26167_);
  nand _77054_ (_26375_, _26374_, _10523_);
  nor _77055_ (_26376_, _10523_, _02860_);
  nor _77056_ (_26377_, _26376_, _03636_);
  and _77057_ (_26378_, _26377_, _26375_);
  and _77058_ (_26379_, _03636_, _03234_);
  or _77059_ (_26380_, _26379_, _03769_);
  nor _77060_ (_26381_, _26380_, _26378_);
  and _77061_ (_26383_, _03769_, \oc8051_golden_model_1.PC [1]);
  or _77062_ (_26384_, _26383_, _26381_);
  nand _77063_ (_26385_, _26384_, _25894_);
  and _77064_ (_26386_, _04317_, _03194_);
  nor _77065_ (_26387_, _26386_, _10534_);
  nand _77066_ (_26388_, _26387_, _26385_);
  nor _77067_ (_26389_, _08698_, _02860_);
  nor _77068_ (_26390_, _26192_, _10077_);
  or _77069_ (_26391_, _26390_, _10535_);
  or _77070_ (_26392_, _26391_, _26389_);
  nand _77071_ (_26394_, _26392_, _26388_);
  nand _77072_ (_26395_, _26394_, _08435_);
  and _77073_ (_26396_, _11572_, _03191_);
  nor _77074_ (_26397_, _26396_, _04135_);
  not _77075_ (_26398_, _26397_);
  nor _77076_ (_26399_, _08435_, _03234_);
  nor _77077_ (_26400_, _26399_, _26398_);
  nand _77078_ (_26401_, _26400_, _26395_);
  nor _77079_ (_26402_, _26397_, _10190_);
  nor _77080_ (_26403_, _26402_, _04138_);
  nand _77081_ (_26405_, _26403_, _26401_);
  and _77082_ (_26406_, _04138_, _10190_);
  nor _77083_ (_26407_, _26406_, _10549_);
  nand _77084_ (_26408_, _26407_, _26405_);
  nor _77085_ (_26409_, _10548_, _02860_);
  nor _77086_ (_26410_, _26409_, _04504_);
  nand _77087_ (_26411_, _26410_, _26408_);
  and _77088_ (_26412_, _03754_, _03234_);
  nor _77089_ (_26413_, _26412_, _03752_);
  and _77090_ (_26414_, _26413_, _26411_);
  or _77091_ (_26416_, _26414_, _26166_);
  nand _77092_ (_26417_, _26416_, _25891_);
  and _77093_ (_26418_, _04317_, _03192_);
  nor _77094_ (_26419_, _26418_, _09958_);
  nand _77095_ (_26420_, _26419_, _26417_);
  and _77096_ (_26421_, \oc8051_golden_model_1.PSW [7], _02860_);
  and _77097_ (_26422_, _26192_, _07888_);
  or _77098_ (_26423_, _26422_, _26421_);
  and _77099_ (_26424_, _26423_, _09958_);
  nor _77100_ (_26425_, _26424_, _15622_);
  and _77101_ (_26427_, _26425_, _26420_);
  or _77102_ (_26428_, _26427_, _26165_);
  and _77103_ (_26429_, _08469_, _04032_);
  nor _77104_ (_26430_, _26429_, _09954_);
  nand _77105_ (_26431_, _26430_, _26428_);
  nor _77106_ (_26432_, _26430_, _10190_);
  nor _77107_ (_26433_, _26432_, _04165_);
  nand _77108_ (_26434_, _26433_, _26431_);
  and _77109_ (_26435_, _04165_, _10190_);
  nor _77110_ (_26436_, _26435_, _08479_);
  nand _77111_ (_26438_, _26436_, _26434_);
  nor _77112_ (_26439_, _08478_, _02860_);
  nor _77113_ (_26440_, _26439_, _03758_);
  nand _77114_ (_26441_, _26440_, _26438_);
  and _77115_ (_26442_, _03758_, _03234_);
  nor _77116_ (_26443_, _26442_, _03760_);
  and _77117_ (_26444_, _26443_, _26441_);
  and _77118_ (_26445_, _03760_, \oc8051_golden_model_1.PC [1]);
  nor _77119_ (_26446_, _26445_, _26444_);
  nand _77120_ (_26447_, _26446_, _26077_);
  nor _77121_ (_26449_, _04317_, _26082_);
  nor _77122_ (_26450_, _26192_, _07888_);
  and _77123_ (_26451_, _07888_, \oc8051_golden_model_1.PC [1]);
  nor _77124_ (_26452_, _26451_, _10577_);
  not _77125_ (_26453_, _26452_);
  nor _77126_ (_26454_, _26453_, _26450_);
  nor _77127_ (_26455_, _26454_, _26449_);
  nand _77128_ (_26456_, _26455_, _26447_);
  nand _77129_ (_26457_, _26456_, _09951_);
  nor _77130_ (_26458_, _09951_, _03234_);
  nor _77131_ (_26460_, _26458_, _08525_);
  nand _77132_ (_26461_, _26460_, _26457_);
  nor _77133_ (_26462_, _08524_, _02860_);
  nor _77134_ (_26463_, _26462_, _08555_);
  and _77135_ (_26464_, _26463_, _26461_);
  and _77136_ (_26465_, _08555_, _10190_);
  or _77137_ (_26466_, _26465_, _03775_);
  nor _77138_ (_26467_, _26466_, _26464_);
  and _77139_ (_26468_, _06433_, _03775_);
  or _77140_ (_26469_, _26468_, _26467_);
  nand _77141_ (_26471_, _26469_, _06328_);
  and _77142_ (_26472_, _04317_, _03179_);
  nor _77143_ (_26473_, _26472_, _03627_);
  nand _77144_ (_26474_, _26473_, _26471_);
  and _77145_ (_26475_, _26238_, _10794_);
  nor _77146_ (_26476_, _10794_, _03234_);
  or _77147_ (_26477_, _26476_, _10599_);
  nor _77148_ (_26478_, _26477_, _26475_);
  nor _77149_ (_26479_, _26478_, _10603_);
  and _77150_ (_26480_, _26479_, _26474_);
  or _77151_ (_26482_, _26480_, _26164_);
  nand _77152_ (_26483_, _26482_, _09936_);
  nor _77153_ (_26484_, _09936_, _02860_);
  nor _77154_ (_26485_, _26484_, _07729_);
  and _77155_ (_26486_, _26485_, _26483_);
  and _77156_ (_26487_, _07729_, _10190_);
  or _77157_ (_26488_, _26487_, _03522_);
  nor _77158_ (_26489_, _26488_, _26486_);
  and _77159_ (_26490_, _06433_, _03522_);
  or _77160_ (_26491_, _26490_, _26489_);
  nand _77161_ (_26493_, _26491_, _25887_);
  and _77162_ (_26494_, _04317_, _03172_);
  nor _77163_ (_26495_, _26494_, _03628_);
  nand _77164_ (_26496_, _26495_, _26493_);
  nor _77165_ (_26497_, _26171_, _10794_);
  and _77166_ (_26498_, _10794_, _10190_);
  nor _77167_ (_26499_, _26498_, _26497_);
  and _77168_ (_26500_, _26499_, _03628_);
  nor _77169_ (_26501_, _26500_, _13062_);
  and _77170_ (_26502_, _26501_, _26496_);
  nor _77171_ (_26504_, _26502_, _26163_);
  and _77172_ (_26505_, _07930_, _03010_);
  or _77173_ (_26506_, _26505_, _26504_);
  and _77174_ (_26507_, _26505_, _03234_);
  nor _77175_ (_26508_, _26507_, _03790_);
  and _77176_ (_26509_, _26508_, _26506_);
  or _77177_ (_26510_, _26509_, _26161_);
  nand _77178_ (_26511_, _26510_, _10828_);
  nor _77179_ (_26512_, _10828_, _03234_);
  nor _77180_ (_26513_, _26512_, _04947_);
  nand _77181_ (_26515_, _26513_, _26511_);
  and _77182_ (_26516_, _04947_, _04317_);
  nor _77183_ (_26517_, _26516_, _03151_);
  and _77184_ (_26518_, _26517_, _26515_);
  and _77185_ (_26519_, _26499_, _03151_);
  nor _77186_ (_26520_, _26519_, _26518_);
  nand _77187_ (_26521_, _26520_, _26160_);
  and _77188_ (_26522_, _12643_, _03228_);
  nor _77189_ (_26523_, _26160_, _10190_);
  nor _77190_ (_26524_, _26523_, _26522_);
  nand _77191_ (_26526_, _26524_, _26521_);
  and _77192_ (_26527_, _26522_, _10190_);
  nor _77193_ (_26528_, _26527_, _04722_);
  nand _77194_ (_26529_, _26528_, _26526_);
  nor _77195_ (_26530_, _04721_, _10190_);
  nor _77196_ (_26531_, _26530_, _03520_);
  and _77197_ (_26532_, _26531_, _26529_);
  or _77198_ (_26533_, _26532_, _26158_);
  nand _77199_ (_26534_, _26533_, _10851_);
  nor _77200_ (_26535_, _10851_, _03234_);
  nor _77201_ (_26537_, _26535_, _25883_);
  and _77202_ (_26538_, _26537_, _26534_);
  or _77203_ (_26539_, _26538_, _26157_);
  and _77204_ (_26540_, _26539_, _10863_);
  and _77205_ (_26541_, _10862_, _03234_);
  nor _77206_ (_26542_, _26541_, _26540_);
  or _77207_ (_26543_, _26542_, _42967_);
  or _77208_ (_26544_, _42963_, \oc8051_golden_model_1.PC [1]);
  and _77209_ (_26545_, _26544_, _41755_);
  and _77210_ (_43328_, _26545_, _26543_);
  and _77211_ (_26547_, _10862_, _03243_);
  and _77212_ (_26548_, _03520_, _03155_);
  and _77213_ (_26549_, _03790_, _03155_);
  nor _77214_ (_26550_, _09949_, _03243_);
  and _77215_ (_26551_, _06569_, _03775_);
  nor _77216_ (_26552_, _09951_, _03243_);
  nor _77217_ (_26553_, _09956_, _03243_);
  and _77218_ (_26554_, _10545_, _03270_);
  nor _77219_ (_26555_, _10520_, _03243_);
  nor _77220_ (_26556_, _03492_, _03155_);
  and _77221_ (_26558_, _03499_, _03626_);
  nor _77222_ (_26559_, _26281_, _03155_);
  and _77223_ (_26560_, _10083_, _03270_);
  and _77224_ (_26561_, _10199_, _10196_);
  nor _77225_ (_26562_, _26561_, _10200_);
  nor _77226_ (_26563_, _26562_, _10261_);
  and _77227_ (_26564_, _10261_, _10188_);
  nor _77228_ (_26565_, _26564_, _26563_);
  or _77229_ (_26566_, _26565_, _04444_);
  and _77230_ (_26567_, _10269_, _03155_);
  and _77231_ (_26569_, _10029_, _10026_);
  nor _77232_ (_26570_, _26569_, _10030_);
  and _77233_ (_26571_, _26570_, _10271_);
  or _77234_ (_26572_, _26571_, _26567_);
  nor _77235_ (_26573_, _26572_, _05831_);
  and _77236_ (_26574_, _03923_, _03920_);
  nor _77237_ (_26575_, _10290_, _03243_);
  nand _77238_ (_26576_, _03922_, _03626_);
  and _77239_ (_26577_, _03922_, _03043_);
  not _77240_ (_26578_, _26577_);
  and _77241_ (_26580_, _10278_, \oc8051_golden_model_1.PC [2]);
  or _77242_ (_26581_, _26580_, _04426_);
  and _77243_ (_26582_, _26581_, _26578_);
  nor _77244_ (_26583_, _10278_, _03270_);
  or _77245_ (_26584_, _26583_, _26582_);
  and _77246_ (_26585_, _26584_, _26576_);
  nand _77247_ (_26586_, _26577_, _03243_);
  nand _77248_ (_26587_, _26586_, _25909_);
  nor _77249_ (_26588_, _26587_, _26585_);
  or _77250_ (_26589_, _26588_, _26575_);
  nor _77251_ (_26591_, _26589_, _26574_);
  nor _77252_ (_26592_, _26591_, _05833_);
  or _77253_ (_26593_, _26592_, _04438_);
  nor _77254_ (_26594_, _26593_, _26573_);
  and _77255_ (_26595_, _04438_, _03243_);
  or _77256_ (_26596_, _26595_, _03570_);
  or _77257_ (_26597_, _26596_, _26594_);
  and _77258_ (_26598_, _26597_, _26566_);
  nor _77259_ (_26599_, _26598_, _10256_);
  nor _77260_ (_26600_, _10255_, _03243_);
  nor _77261_ (_26602_, _26600_, _03516_);
  not _77262_ (_26603_, _26602_);
  nor _77263_ (_26604_, _26603_, _26599_);
  and _77264_ (_26605_, _03516_, _03155_);
  nor _77265_ (_26606_, _26605_, _26604_);
  or _77266_ (_26607_, _26606_, _04746_);
  or _77267_ (_26608_, _03920_, _03203_);
  and _77268_ (_26609_, _26608_, _26607_);
  or _77269_ (_26610_, _26609_, _03568_);
  and _77270_ (_26611_, _03568_, _03155_);
  nor _77271_ (_26613_, _26611_, _26212_);
  nand _77272_ (_26614_, _26613_, _26610_);
  nor _77273_ (_26615_, _10307_, _03243_);
  nor _77274_ (_26616_, _26615_, _03575_);
  nand _77275_ (_26617_, _26616_, _26614_);
  and _77276_ (_26618_, _03575_, _03155_);
  nor _77277_ (_26619_, _26618_, _26220_);
  nand _77278_ (_26620_, _26619_, _26617_);
  nor _77279_ (_26621_, _10316_, _03243_);
  nor _77280_ (_26622_, _26621_, _03512_);
  nand _77281_ (_26624_, _26622_, _26620_);
  and _77282_ (_26625_, _03512_, _03155_);
  nor _77283_ (_26626_, _26625_, _10249_);
  nand _77284_ (_26627_, _26626_, _26624_);
  and _77285_ (_26628_, _03920_, _10249_);
  nor _77286_ (_26629_, _26628_, _03511_);
  nand _77287_ (_26630_, _26629_, _26627_);
  and _77288_ (_26631_, _03511_, _03155_);
  nor _77289_ (_26632_, _26631_, _10326_);
  nand _77290_ (_26633_, _26632_, _26630_);
  and _77291_ (_26634_, _10360_, _10187_);
  not _77292_ (_26635_, _26562_);
  nor _77293_ (_26636_, _26635_, _10360_);
  or _77294_ (_26637_, _26636_, _26634_);
  nor _77295_ (_26638_, _26637_, _10325_);
  nor _77296_ (_26639_, _26638_, _03657_);
  nand _77297_ (_26640_, _26639_, _26633_);
  nor _77298_ (_26641_, _26635_, _10116_);
  and _77299_ (_26642_, _10187_, _10116_);
  nor _77300_ (_26643_, _26642_, _26641_);
  nor _77301_ (_26646_, _26643_, _10328_);
  nor _77302_ (_26647_, _26646_, _03527_);
  nand _77303_ (_26648_, _26647_, _26640_);
  and _77304_ (_26649_, _10382_, _10187_);
  not _77305_ (_26650_, _26649_);
  nor _77306_ (_26651_, _26635_, _10382_);
  nor _77307_ (_26652_, _26651_, _03998_);
  and _77308_ (_26653_, _26652_, _26650_);
  nor _77309_ (_26654_, _26653_, _03638_);
  nand _77310_ (_26655_, _26654_, _26648_);
  and _77311_ (_26657_, _10398_, _10188_);
  nor _77312_ (_26658_, _26562_, _10398_);
  or _77313_ (_26659_, _26658_, _10085_);
  nor _77314_ (_26660_, _26659_, _26657_);
  nor _77315_ (_26661_, _26660_, _10083_);
  and _77316_ (_26662_, _26661_, _26655_);
  or _77317_ (_26663_, _26662_, _26560_);
  nand _77318_ (_26664_, _26663_, _03506_);
  and _77319_ (_26665_, _03505_, _03626_);
  nor _77320_ (_26666_, _26665_, _04743_);
  nand _77321_ (_26668_, _26666_, _26664_);
  nor _77322_ (_26669_, _03920_, _03200_);
  nor _77323_ (_26670_, _26669_, _26282_);
  and _77324_ (_26671_, _26670_, _26668_);
  or _77325_ (_26672_, _26671_, _26559_);
  nand _77326_ (_26673_, _26672_, _10415_);
  nor _77327_ (_26674_, _10415_, _03243_);
  nor _77328_ (_26675_, _26674_, _03607_);
  nand _77329_ (_26676_, _26675_, _26673_);
  and _77330_ (_26677_, _03607_, _03155_);
  nor _77331_ (_26679_, _26677_, _10420_);
  nand _77332_ (_26680_, _26679_, _26676_);
  and _77333_ (_26681_, _03920_, _10420_);
  nor _77334_ (_26682_, _26681_, _03606_);
  nand _77335_ (_26683_, _26682_, _26680_);
  and _77336_ (_26684_, _03606_, _03155_);
  nor _77337_ (_26685_, _26684_, _26302_);
  and _77338_ (_26686_, _26685_, _26683_);
  nor _77339_ (_26687_, _10426_, _03243_);
  or _77340_ (_26688_, _26687_, _26686_);
  nand _77341_ (_26690_, _26688_, _10430_);
  nor _77342_ (_26691_, _10430_, _03155_);
  nor _77343_ (_26692_, _26691_, _03311_);
  nand _77344_ (_26693_, _26692_, _26690_);
  nor _77345_ (_26694_, _03254_, _03270_);
  nor _77346_ (_26695_, _26694_, _03499_);
  and _77347_ (_26696_, _26695_, _26693_);
  or _77348_ (_26697_, _26696_, _26558_);
  nand _77349_ (_26698_, _26697_, _04853_);
  and _77350_ (_26699_, _03920_, _03223_);
  nor _77351_ (_26701_, _26699_, _03632_);
  nand _77352_ (_26702_, _26701_, _26698_);
  and _77353_ (_26703_, _10187_, _03632_);
  not _77354_ (_26704_, _26703_);
  and _77355_ (_26705_, _26704_, _03492_);
  and _77356_ (_26706_, _26705_, _26702_);
  or _77357_ (_26707_, _26706_, _26556_);
  nand _77358_ (_26708_, _26707_, _03480_);
  nor _77359_ (_26709_, _03480_, _03155_);
  nor _77360_ (_26710_, _26709_, _03221_);
  nand _77361_ (_26712_, _26710_, _26708_);
  and _77362_ (_26713_, _10187_, _03221_);
  nor _77363_ (_26714_, _26713_, _26330_);
  nand _77364_ (_26715_, _26714_, _26712_);
  nor _77365_ (_26716_, _10081_, _03243_);
  nor _77366_ (_26717_, _26716_, _03745_);
  and _77367_ (_26718_, _26717_, _26715_);
  and _77368_ (_26719_, _03745_, _03155_);
  or _77369_ (_26720_, _26719_, _03187_);
  nor _77370_ (_26721_, _26720_, _26718_);
  and _77371_ (_26723_, _03920_, _03187_);
  or _77372_ (_26724_, _26723_, _26721_);
  nand _77373_ (_26725_, _26724_, _10459_);
  not _77374_ (_26726_, _05773_);
  nor _77375_ (_26727_, _26570_, _10459_);
  nor _77376_ (_26728_, _26727_, _26726_);
  nand _77377_ (_26729_, _26728_, _26725_);
  not _77378_ (_26730_, _05774_);
  nor _77379_ (_26731_, _05773_, _03626_);
  nor _77380_ (_26732_, _26731_, _26730_);
  nand _77381_ (_26734_, _26732_, _26729_);
  nor _77382_ (_26735_, _05774_, _03155_);
  nor _77383_ (_26736_, _26735_, _03437_);
  and _77384_ (_26737_, _26736_, _26734_);
  and _77385_ (_26738_, _10187_, _03437_);
  or _77386_ (_26739_, _26738_, _08385_);
  nor _77387_ (_26740_, _26739_, _26737_);
  and _77388_ (_26741_, _08385_, _03626_);
  or _77389_ (_26742_, _26741_, _26740_);
  nand _77390_ (_26743_, _26742_, _25897_);
  nor _77391_ (_26745_, _25897_, _03267_);
  nor _77392_ (_26746_, _26745_, _03744_);
  nand _77393_ (_26747_, _26746_, _26743_);
  and _77394_ (_26748_, _03744_, _03155_);
  nor _77395_ (_26749_, _26748_, _03189_);
  nand _77396_ (_26750_, _26749_, _26747_);
  and _77397_ (_26751_, _03920_, _03189_);
  nor _77398_ (_26752_, _26751_, _10076_);
  nand _77399_ (_26753_, _26752_, _26750_);
  not _77400_ (_26754_, _10520_);
  and _77401_ (_26756_, _08698_, _03155_);
  and _77402_ (_26757_, _26570_, _10077_);
  or _77403_ (_26758_, _26757_, _26756_);
  and _77404_ (_26759_, _26758_, _10076_);
  nor _77405_ (_26760_, _26759_, _26754_);
  and _77406_ (_26761_, _26760_, _26753_);
  or _77407_ (_26762_, _26761_, _26555_);
  nand _77408_ (_26763_, _26762_, _10523_);
  nor _77409_ (_26764_, _10523_, _03155_);
  nor _77410_ (_26765_, _26764_, _03636_);
  and _77411_ (_26767_, _26765_, _26763_);
  and _77412_ (_26768_, _10187_, _03636_);
  or _77413_ (_26769_, _26768_, _03769_);
  nor _77414_ (_26770_, _26769_, _26767_);
  and _77415_ (_26771_, _03769_, _03626_);
  or _77416_ (_26772_, _26771_, _26770_);
  nand _77417_ (_26773_, _26772_, _25894_);
  and _77418_ (_26774_, _03920_, _03194_);
  nor _77419_ (_26775_, _26774_, _10534_);
  nand _77420_ (_26776_, _26775_, _26773_);
  nor _77421_ (_26778_, _26570_, _10077_);
  nor _77422_ (_26779_, _08698_, _03155_);
  nor _77423_ (_26780_, _26779_, _10535_);
  not _77424_ (_26781_, _26780_);
  nor _77425_ (_26782_, _26781_, _26778_);
  nor _77426_ (_26783_, _26782_, _10545_);
  and _77427_ (_26784_, _26783_, _26776_);
  or _77428_ (_26785_, _26784_, _26554_);
  nand _77429_ (_26786_, _26785_, _10548_);
  nor _77430_ (_26787_, _10548_, _03155_);
  nor _77431_ (_26789_, _26787_, _03754_);
  nand _77432_ (_26790_, _26789_, _26786_);
  and _77433_ (_26791_, _10187_, _03754_);
  nor _77434_ (_26792_, _26791_, _03752_);
  and _77435_ (_26793_, _26792_, _26790_);
  and _77436_ (_26794_, _03752_, _03626_);
  or _77437_ (_26795_, _26794_, _26793_);
  nand _77438_ (_26796_, _26795_, _25891_);
  and _77439_ (_26797_, _03920_, _03192_);
  nor _77440_ (_26798_, _26797_, _09958_);
  nand _77441_ (_26800_, _26798_, _26796_);
  and _77442_ (_26801_, _03155_, \oc8051_golden_model_1.PSW [7]);
  and _77443_ (_26802_, _26570_, _07888_);
  or _77444_ (_26803_, _26802_, _26801_);
  and _77445_ (_26804_, _26803_, _09958_);
  nor _77446_ (_26805_, _26804_, _10560_);
  and _77447_ (_26806_, _26805_, _26800_);
  or _77448_ (_26807_, _26806_, _26553_);
  nand _77449_ (_26808_, _26807_, _08478_);
  nor _77450_ (_26809_, _08478_, _03155_);
  nor _77451_ (_26811_, _26809_, _03758_);
  and _77452_ (_26812_, _26811_, _26808_);
  and _77453_ (_26813_, _10187_, _03758_);
  or _77454_ (_26814_, _26813_, _03760_);
  nor _77455_ (_26815_, _26814_, _26812_);
  and _77456_ (_26816_, _03760_, _03626_);
  or _77457_ (_26817_, _26816_, _26815_);
  nand _77458_ (_26818_, _26817_, _26082_);
  and _77459_ (_26819_, _03920_, _03183_);
  nor _77460_ (_26820_, _26819_, _10576_);
  nand _77461_ (_26822_, _26820_, _26818_);
  nor _77462_ (_26823_, _26570_, _07888_);
  nor _77463_ (_26824_, _03155_, \oc8051_golden_model_1.PSW [7]);
  nor _77464_ (_26825_, _26824_, _10577_);
  not _77465_ (_26826_, _26825_);
  nor _77466_ (_26827_, _26826_, _26823_);
  nor _77467_ (_26828_, _26827_, _10581_);
  and _77468_ (_26829_, _26828_, _26822_);
  or _77469_ (_26830_, _26829_, _26552_);
  nand _77470_ (_26831_, _26830_, _08524_);
  nor _77471_ (_26833_, _08524_, _03155_);
  nor _77472_ (_26834_, _26833_, _08555_);
  nand _77473_ (_26835_, _26834_, _26831_);
  and _77474_ (_26836_, _08555_, _03243_);
  nor _77475_ (_26837_, _26836_, _03775_);
  and _77476_ (_26838_, _26837_, _26835_);
  or _77477_ (_26839_, _26838_, _26551_);
  nand _77478_ (_26840_, _26839_, _06328_);
  and _77479_ (_26841_, _03920_, _03179_);
  nor _77480_ (_26842_, _26841_, _03627_);
  nand _77481_ (_26844_, _26842_, _26840_);
  nor _77482_ (_26845_, _10794_, _10187_);
  and _77483_ (_26846_, _26635_, _10794_);
  or _77484_ (_26847_, _26846_, _10599_);
  nor _77485_ (_26848_, _26847_, _26845_);
  nor _77486_ (_26849_, _26848_, _10603_);
  and _77487_ (_26850_, _26849_, _26844_);
  or _77488_ (_26851_, _26850_, _26550_);
  nand _77489_ (_26852_, _26851_, _09936_);
  nor _77490_ (_26853_, _09936_, _03155_);
  nor _77491_ (_26855_, _26853_, _07729_);
  and _77492_ (_26856_, _26855_, _26852_);
  and _77493_ (_26857_, _07729_, _03243_);
  or _77494_ (_26858_, _26857_, _03522_);
  nor _77495_ (_26859_, _26858_, _26856_);
  and _77496_ (_26860_, _06569_, _03522_);
  or _77497_ (_26861_, _26860_, _26859_);
  nand _77498_ (_26862_, _26861_, _25887_);
  and _77499_ (_26863_, _03920_, _03172_);
  nor _77500_ (_26864_, _26863_, _03628_);
  nand _77501_ (_26866_, _26864_, _26862_);
  nor _77502_ (_26867_, _26562_, _10794_);
  and _77503_ (_26868_, _10794_, _10188_);
  nor _77504_ (_26869_, _26868_, _26867_);
  and _77505_ (_26870_, _26869_, _03628_);
  nor _77506_ (_26871_, _26870_, _10822_);
  nand _77507_ (_26872_, _26871_, _26866_);
  nor _77508_ (_26873_, _10821_, _03243_);
  nor _77509_ (_26874_, _26873_, _03790_);
  and _77510_ (_26875_, _26874_, _26872_);
  or _77511_ (_26877_, _26875_, _26549_);
  nand _77512_ (_26878_, _26877_, _10828_);
  nor _77513_ (_26879_, _10828_, _03270_);
  nor _77514_ (_26880_, _26879_, _04947_);
  nand _77515_ (_26881_, _26880_, _26878_);
  and _77516_ (_26882_, _04947_, _03920_);
  nor _77517_ (_26883_, _26882_, _03151_);
  nand _77518_ (_26884_, _26883_, _26881_);
  and _77519_ (_26885_, _26869_, _03151_);
  nor _77520_ (_26886_, _26885_, _10845_);
  nand _77521_ (_26888_, _26886_, _26884_);
  nor _77522_ (_26889_, _10844_, _03243_);
  nor _77523_ (_26890_, _26889_, _03520_);
  and _77524_ (_26891_, _26890_, _26888_);
  or _77525_ (_26892_, _26891_, _26548_);
  nand _77526_ (_26893_, _26892_, _10851_);
  nor _77527_ (_26894_, _10851_, _03270_);
  nor _77528_ (_26895_, _26894_, _25883_);
  nand _77529_ (_26896_, _26895_, _26893_);
  and _77530_ (_26897_, _25883_, _03920_);
  nor _77531_ (_26899_, _26897_, _10862_);
  and _77532_ (_26900_, _26899_, _26896_);
  or _77533_ (_26901_, _26900_, _26547_);
  or _77534_ (_26902_, _26901_, _42967_);
  or _77535_ (_26903_, _42963_, \oc8051_golden_model_1.PC [2]);
  and _77536_ (_26904_, _26903_, _41755_);
  and _77537_ (_43329_, _26904_, _26902_);
  and _77538_ (_26905_, _10862_, _03677_);
  and _77539_ (_26906_, _03520_, _03280_);
  nor _77540_ (_26907_, _10828_, _03677_);
  nor _77541_ (_26909_, _09949_, _03677_);
  nor _77542_ (_26910_, _09951_, _03677_);
  nor _77543_ (_26911_, _09956_, _03677_);
  and _77544_ (_26912_, _10545_, _03293_);
  nor _77545_ (_26913_, _10520_, _03677_);
  nor _77546_ (_26914_, _03493_, _03280_);
  or _77547_ (_26915_, _26914_, _03221_);
  and _77548_ (_26916_, _03499_, _03675_);
  nor _77549_ (_26917_, _03742_, _03200_);
  and _77550_ (_26918_, _10083_, _03293_);
  and _77551_ (_26920_, _10261_, _10183_);
  or _77552_ (_26921_, _10185_, _10184_);
  and _77553_ (_26922_, _26921_, _10201_);
  nor _77554_ (_26923_, _26921_, _10201_);
  nor _77555_ (_26924_, _26923_, _26922_);
  nor _77556_ (_26925_, _26924_, _10261_);
  nor _77557_ (_26926_, _26925_, _26920_);
  or _77558_ (_26927_, _26926_, _04444_);
  and _77559_ (_26928_, _10269_, _03280_);
  or _77560_ (_26929_, _10019_, _10018_);
  and _77561_ (_26930_, _26929_, _10031_);
  nor _77562_ (_26931_, _26929_, _10031_);
  nor _77563_ (_26932_, _26931_, _26930_);
  and _77564_ (_26933_, _26932_, _10271_);
  or _77565_ (_26934_, _26933_, _26928_);
  nor _77566_ (_26935_, _26934_, _05831_);
  nor _77567_ (_26936_, _04762_, _03742_);
  nand _77568_ (_26937_, _03922_, _03675_);
  and _77569_ (_26938_, _10278_, \oc8051_golden_model_1.PC [3]);
  or _77570_ (_26939_, _26938_, _04426_);
  and _77571_ (_26942_, _26939_, _26578_);
  nor _77572_ (_26943_, _10278_, _03293_);
  or _77573_ (_26944_, _26943_, _26942_);
  and _77574_ (_26945_, _26944_, _26937_);
  nand _77575_ (_26946_, _26577_, _03677_);
  nand _77576_ (_26947_, _26946_, _10290_);
  or _77577_ (_26948_, _26947_, _26945_);
  and _77578_ (_26949_, _26948_, _04762_);
  nor _77579_ (_26950_, _26949_, _26936_);
  nor _77580_ (_26951_, _10290_, _03677_);
  nor _77581_ (_26953_, _26951_, _26950_);
  nor _77582_ (_26954_, _26953_, _05833_);
  or _77583_ (_26955_, _26954_, _04438_);
  nor _77584_ (_26956_, _26955_, _26935_);
  and _77585_ (_26957_, _04438_, _03677_);
  or _77586_ (_26958_, _26957_, _03570_);
  or _77587_ (_26959_, _26958_, _26956_);
  and _77588_ (_26960_, _26959_, _26927_);
  nor _77589_ (_26961_, _26960_, _10256_);
  nor _77590_ (_26962_, _10255_, _03677_);
  nor _77591_ (_26964_, _26962_, _03516_);
  not _77592_ (_26965_, _26964_);
  nor _77593_ (_26966_, _26965_, _26961_);
  and _77594_ (_26967_, _03516_, _03280_);
  nor _77595_ (_26968_, _26967_, _26966_);
  or _77596_ (_26969_, _26968_, _04746_);
  or _77597_ (_26970_, _03742_, _03203_);
  and _77598_ (_26971_, _26970_, _26969_);
  or _77599_ (_26972_, _26971_, _03568_);
  and _77600_ (_26973_, _03568_, _03280_);
  nor _77601_ (_26975_, _26973_, _26212_);
  nand _77602_ (_26976_, _26975_, _26972_);
  nor _77603_ (_26977_, _10307_, _03677_);
  nor _77604_ (_26978_, _26977_, _03575_);
  nand _77605_ (_26979_, _26978_, _26976_);
  and _77606_ (_26980_, _03575_, _03280_);
  nor _77607_ (_26981_, _26980_, _26220_);
  nand _77608_ (_26982_, _26981_, _26979_);
  nor _77609_ (_26983_, _10316_, _03677_);
  nor _77610_ (_26984_, _26983_, _03512_);
  nand _77611_ (_26986_, _26984_, _26982_);
  and _77612_ (_26987_, _03512_, _03280_);
  nor _77613_ (_26988_, _26987_, _10249_);
  nand _77614_ (_26989_, _26988_, _26986_);
  and _77615_ (_26990_, _03742_, _10249_);
  nor _77616_ (_26991_, _26990_, _03511_);
  nand _77617_ (_26992_, _26991_, _26989_);
  and _77618_ (_26993_, _03511_, _03280_);
  nor _77619_ (_26994_, _26993_, _10326_);
  nand _77620_ (_26995_, _26994_, _26992_);
  and _77621_ (_26997_, _10360_, _10182_);
  not _77622_ (_26998_, _26924_);
  nor _77623_ (_26999_, _26998_, _10360_);
  or _77624_ (_27000_, _26999_, _10325_);
  nor _77625_ (_27001_, _27000_, _26997_);
  nor _77626_ (_27002_, _27001_, _03657_);
  nand _77627_ (_27003_, _27002_, _26995_);
  nor _77628_ (_27004_, _26998_, _10116_);
  and _77629_ (_27005_, _10182_, _10116_);
  nor _77630_ (_27006_, _27005_, _27004_);
  nor _77631_ (_27008_, _27006_, _10328_);
  nor _77632_ (_27009_, _27008_, _03527_);
  nand _77633_ (_27010_, _27009_, _27003_);
  nor _77634_ (_27011_, _26998_, _10382_);
  not _77635_ (_27012_, _27011_);
  and _77636_ (_27013_, _10382_, _10182_);
  nor _77637_ (_27014_, _27013_, _03998_);
  and _77638_ (_27015_, _27014_, _27012_);
  nor _77639_ (_27016_, _27015_, _03638_);
  nand _77640_ (_27017_, _27016_, _27010_);
  and _77641_ (_27019_, _10398_, _10182_);
  and _77642_ (_27020_, _26924_, _10399_);
  or _77643_ (_27021_, _27020_, _27019_);
  and _77644_ (_27022_, _27021_, _03638_);
  nor _77645_ (_27023_, _27022_, _10083_);
  and _77646_ (_27024_, _27023_, _27017_);
  or _77647_ (_27025_, _27024_, _26918_);
  nand _77648_ (_27026_, _27025_, _03506_);
  and _77649_ (_27027_, _03505_, _03675_);
  nor _77650_ (_27028_, _27027_, _04743_);
  and _77651_ (_27030_, _27028_, _27026_);
  or _77652_ (_27031_, _27030_, _26917_);
  nand _77653_ (_27032_, _27031_, _26281_);
  nor _77654_ (_27033_, _26281_, _03675_);
  nor _77655_ (_27034_, _27033_, _25991_);
  nand _77656_ (_27035_, _27034_, _27032_);
  nor _77657_ (_27036_, _10415_, _03677_);
  nor _77658_ (_27037_, _27036_, _03607_);
  nand _77659_ (_27038_, _27037_, _27035_);
  and _77660_ (_27039_, _03607_, _03280_);
  nor _77661_ (_27040_, _27039_, _10420_);
  nand _77662_ (_27041_, _27040_, _27038_);
  and _77663_ (_27042_, _03742_, _10420_);
  nor _77664_ (_27043_, _27042_, _03606_);
  nand _77665_ (_27044_, _27043_, _27041_);
  and _77666_ (_27045_, _03606_, _03280_);
  nor _77667_ (_27046_, _27045_, _26302_);
  and _77668_ (_27047_, _27046_, _27044_);
  nor _77669_ (_27048_, _10426_, _03677_);
  or _77670_ (_27049_, _27048_, _27047_);
  nand _77671_ (_27052_, _27049_, _10430_);
  nor _77672_ (_27053_, _10430_, _03280_);
  nor _77673_ (_27054_, _27053_, _03311_);
  nand _77674_ (_27055_, _27054_, _27052_);
  nor _77675_ (_27056_, _03254_, _03293_);
  nor _77676_ (_27057_, _27056_, _03499_);
  and _77677_ (_27058_, _27057_, _27055_);
  or _77678_ (_27059_, _27058_, _26916_);
  nand _77679_ (_27060_, _27059_, _04853_);
  and _77680_ (_27061_, _03742_, _03223_);
  nor _77681_ (_27063_, _27061_, _03632_);
  nand _77682_ (_27064_, _27063_, _27060_);
  and _77683_ (_27065_, _10182_, _03632_);
  nor _77684_ (_27066_, _27065_, _26322_);
  and _77685_ (_27067_, _27066_, _27064_);
  or _77686_ (_27068_, _27067_, _26915_);
  and _77687_ (_27069_, _10182_, _03221_);
  nor _77688_ (_27070_, _27069_, _26330_);
  nand _77689_ (_27071_, _27070_, _27068_);
  nor _77690_ (_27072_, _10081_, _03677_);
  nor _77691_ (_27074_, _27072_, _03745_);
  and _77692_ (_27075_, _27074_, _27071_);
  and _77693_ (_27076_, _03745_, _03280_);
  or _77694_ (_27077_, _27076_, _03187_);
  or _77695_ (_27078_, _27077_, _27075_);
  and _77696_ (_27079_, _03742_, _03187_);
  nor _77697_ (_27080_, _27079_, _10458_);
  nand _77698_ (_27081_, _27080_, _27078_);
  and _77699_ (_27082_, _26932_, _10458_);
  nor _77700_ (_27083_, _27082_, _06055_);
  nand _77701_ (_27085_, _27083_, _27081_);
  nor _77702_ (_27086_, _05775_, _03280_);
  nor _77703_ (_27087_, _27086_, _03437_);
  nand _77704_ (_27088_, _27087_, _27085_);
  and _77705_ (_27089_, _10182_, _03437_);
  nor _77706_ (_27090_, _27089_, _08385_);
  and _77707_ (_27091_, _27090_, _27088_);
  and _77708_ (_27092_, _08385_, _03675_);
  or _77709_ (_27093_, _27092_, _27091_);
  nand _77710_ (_27094_, _27093_, _25897_);
  nor _77711_ (_27096_, _25897_, _03289_);
  nor _77712_ (_27097_, _27096_, _03744_);
  nand _77713_ (_27098_, _27097_, _27094_);
  and _77714_ (_27099_, _03744_, _03280_);
  nor _77715_ (_27100_, _27099_, _03189_);
  nand _77716_ (_27101_, _27100_, _27098_);
  and _77717_ (_27102_, _03742_, _03189_);
  nor _77718_ (_27103_, _27102_, _10076_);
  nand _77719_ (_27104_, _27103_, _27101_);
  and _77720_ (_27105_, _08698_, _03280_);
  and _77721_ (_27107_, _26932_, _10077_);
  or _77722_ (_27108_, _27107_, _27105_);
  and _77723_ (_27109_, _27108_, _10076_);
  nor _77724_ (_27110_, _27109_, _26754_);
  and _77725_ (_27111_, _27110_, _27104_);
  or _77726_ (_27112_, _27111_, _26913_);
  nand _77727_ (_27113_, _27112_, _10523_);
  nor _77728_ (_27114_, _10523_, _03280_);
  nor _77729_ (_27115_, _27114_, _03636_);
  and _77730_ (_27116_, _27115_, _27113_);
  and _77731_ (_27118_, _10182_, _03636_);
  or _77732_ (_27119_, _27118_, _03769_);
  nor _77733_ (_27120_, _27119_, _27116_);
  and _77734_ (_27121_, _03769_, _03675_);
  or _77735_ (_27122_, _27121_, _27120_);
  nand _77736_ (_27123_, _27122_, _25894_);
  and _77737_ (_27124_, _03742_, _03194_);
  nor _77738_ (_27125_, _27124_, _10534_);
  nand _77739_ (_27126_, _27125_, _27123_);
  nor _77740_ (_27127_, _26932_, _10077_);
  nor _77741_ (_27129_, _08698_, _03280_);
  nor _77742_ (_27130_, _27129_, _10535_);
  not _77743_ (_27131_, _27130_);
  nor _77744_ (_27132_, _27131_, _27127_);
  nor _77745_ (_27133_, _27132_, _10545_);
  and _77746_ (_27134_, _27133_, _27126_);
  or _77747_ (_27135_, _27134_, _26912_);
  nand _77748_ (_27136_, _27135_, _10548_);
  nor _77749_ (_27137_, _10548_, _03280_);
  nor _77750_ (_27138_, _27137_, _04504_);
  nand _77751_ (_27140_, _27138_, _27136_);
  and _77752_ (_27141_, _10182_, _03754_);
  nor _77753_ (_27142_, _27141_, _03752_);
  and _77754_ (_27143_, _27142_, _27140_);
  and _77755_ (_27144_, _03752_, _03675_);
  or _77756_ (_27145_, _27144_, _27143_);
  nand _77757_ (_27146_, _27145_, _25891_);
  and _77758_ (_27147_, _03742_, _03192_);
  nor _77759_ (_27148_, _27147_, _09958_);
  nand _77760_ (_27149_, _27148_, _27146_);
  and _77761_ (_27151_, _03280_, \oc8051_golden_model_1.PSW [7]);
  and _77762_ (_27152_, _26932_, _07888_);
  or _77763_ (_27153_, _27152_, _27151_);
  and _77764_ (_27154_, _27153_, _09958_);
  nor _77765_ (_27155_, _27154_, _10560_);
  and _77766_ (_27156_, _27155_, _27149_);
  or _77767_ (_27157_, _27156_, _26911_);
  nand _77768_ (_27158_, _27157_, _08478_);
  nor _77769_ (_27159_, _08478_, _03280_);
  nor _77770_ (_27160_, _27159_, _03758_);
  and _77771_ (_27162_, _27160_, _27158_);
  and _77772_ (_27163_, _10182_, _03758_);
  or _77773_ (_27164_, _27163_, _03760_);
  nor _77774_ (_27165_, _27164_, _27162_);
  and _77775_ (_27166_, _03760_, _03675_);
  or _77776_ (_27167_, _27166_, _27165_);
  nand _77777_ (_27168_, _27167_, _26082_);
  and _77778_ (_27169_, _03742_, _03183_);
  nor _77779_ (_27170_, _27169_, _10576_);
  nand _77780_ (_27171_, _27170_, _27168_);
  nor _77781_ (_27173_, _26932_, _07888_);
  nor _77782_ (_27174_, _03280_, \oc8051_golden_model_1.PSW [7]);
  nor _77783_ (_27175_, _27174_, _10577_);
  not _77784_ (_27176_, _27175_);
  nor _77785_ (_27177_, _27176_, _27173_);
  nor _77786_ (_27178_, _27177_, _10581_);
  and _77787_ (_27179_, _27178_, _27171_);
  or _77788_ (_27180_, _27179_, _26910_);
  nand _77789_ (_27181_, _27180_, _08524_);
  nor _77790_ (_27182_, _08524_, _03280_);
  nor _77791_ (_27184_, _27182_, _08555_);
  and _77792_ (_27185_, _27184_, _27181_);
  and _77793_ (_27186_, _08555_, _03677_);
  or _77794_ (_27187_, _27186_, _03775_);
  nor _77795_ (_27188_, _27187_, _27185_);
  and _77796_ (_27189_, _06524_, _03775_);
  or _77797_ (_27190_, _27189_, _27188_);
  nand _77798_ (_27191_, _27190_, _06328_);
  and _77799_ (_27192_, _03742_, _03179_);
  nor _77800_ (_27193_, _27192_, _03627_);
  nand _77801_ (_27195_, _27193_, _27191_);
  and _77802_ (_27196_, _26998_, _10794_);
  nor _77803_ (_27197_, _10794_, _10182_);
  or _77804_ (_27198_, _27197_, _10599_);
  or _77805_ (_27199_, _27198_, _27196_);
  and _77806_ (_27200_, _27199_, _09949_);
  and _77807_ (_27201_, _27200_, _27195_);
  or _77808_ (_27202_, _27201_, _26909_);
  nand _77809_ (_27203_, _27202_, _09936_);
  nor _77810_ (_27204_, _09936_, _03280_);
  nor _77811_ (_27206_, _27204_, _07729_);
  and _77812_ (_27207_, _27206_, _27203_);
  and _77813_ (_27208_, _07729_, _03677_);
  or _77814_ (_27209_, _27208_, _03522_);
  nor _77815_ (_27210_, _27209_, _27207_);
  and _77816_ (_27211_, _06524_, _03522_);
  or _77817_ (_27212_, _27211_, _27210_);
  nand _77818_ (_27213_, _27212_, _25887_);
  and _77819_ (_27214_, _03742_, _03172_);
  nor _77820_ (_27215_, _27214_, _03628_);
  nand _77821_ (_27217_, _27215_, _27213_);
  nor _77822_ (_27218_, _26924_, _10794_);
  and _77823_ (_27219_, _10794_, _10183_);
  nor _77824_ (_27220_, _27219_, _27218_);
  and _77825_ (_27221_, _27220_, _03628_);
  nor _77826_ (_27222_, _27221_, _10822_);
  nand _77827_ (_27223_, _27222_, _27217_);
  nor _77828_ (_27224_, _10821_, _03677_);
  nor _77829_ (_27225_, _27224_, _03790_);
  nand _77830_ (_27226_, _27225_, _27223_);
  not _77831_ (_27228_, _10828_);
  and _77832_ (_27229_, _03790_, _03280_);
  nor _77833_ (_27230_, _27229_, _27228_);
  and _77834_ (_27231_, _27230_, _27226_);
  or _77835_ (_27232_, _27231_, _26907_);
  nand _77836_ (_27233_, _27232_, _04533_);
  and _77837_ (_27234_, _04947_, _03742_);
  nor _77838_ (_27235_, _27234_, _03151_);
  nand _77839_ (_27236_, _27235_, _27233_);
  and _77840_ (_27237_, _27220_, _03151_);
  nor _77841_ (_27239_, _27237_, _10845_);
  nand _77842_ (_27240_, _27239_, _27236_);
  nor _77843_ (_27241_, _10844_, _03677_);
  nor _77844_ (_27242_, _27241_, _03520_);
  and _77845_ (_27243_, _27242_, _27240_);
  or _77846_ (_27244_, _27243_, _26906_);
  nand _77847_ (_27245_, _27244_, _10851_);
  nor _77848_ (_27246_, _10851_, _03293_);
  nor _77849_ (_27247_, _27246_, _25883_);
  nand _77850_ (_27248_, _27247_, _27245_);
  and _77851_ (_27250_, _25883_, _03742_);
  nor _77852_ (_27251_, _27250_, _10862_);
  and _77853_ (_27252_, _27251_, _27248_);
  or _77854_ (_27253_, _27252_, _26905_);
  or _77855_ (_27254_, _27253_, _42967_);
  or _77856_ (_27255_, _42963_, \oc8051_golden_model_1.PC [3]);
  and _77857_ (_27256_, _27255_, _41755_);
  and _77858_ (_43330_, _27256_, _27254_);
  nand _77859_ (_27257_, _06195_, _04947_);
  nor _77860_ (_27258_, _10036_, _10034_);
  nor _77861_ (_27259_, _27258_, _10037_);
  or _77862_ (_27260_, _27259_, \oc8051_golden_model_1.PSW [7]);
  or _77863_ (_27261_, _10015_, _07888_);
  and _77864_ (_27262_, _27261_, _09958_);
  and _77865_ (_27263_, _27262_, _27260_);
  or _77866_ (_27264_, _26281_, _10015_);
  and _77867_ (_27265_, _09938_, \oc8051_golden_model_1.PC [4]);
  nor _77868_ (_27266_, _09938_, \oc8051_golden_model_1.PC [4]);
  nor _77869_ (_27267_, _27266_, _27265_);
  not _77870_ (_27268_, _27267_);
  nand _77871_ (_27271_, _27268_, _10083_);
  not _77872_ (_27272_, _11574_);
  nand _77873_ (_27273_, _10016_, _03512_);
  or _77874_ (_27274_, _27267_, _10307_);
  and _77875_ (_27275_, _27259_, _10271_);
  and _77876_ (_27276_, _10269_, _10015_);
  or _77877_ (_27277_, _27276_, _05831_);
  or _77878_ (_27278_, _27277_, _27275_);
  nand _77879_ (_27279_, _06195_, _03923_);
  or _77880_ (_27280_, _27267_, _10278_);
  not _77881_ (_27282_, _10278_);
  or _77882_ (_27283_, _27282_, \oc8051_golden_model_1.PC [4]);
  and _77883_ (_27284_, _27283_, _27280_);
  or _77884_ (_27285_, _27284_, _04426_);
  nand _77885_ (_27286_, _10016_, _04426_);
  and _77886_ (_27287_, _27286_, _10275_);
  and _77887_ (_27288_, _27287_, _27285_);
  and _77888_ (_27289_, _27267_, _26577_);
  or _77889_ (_27290_, _27289_, _03923_);
  or _77890_ (_27291_, _27290_, _27288_);
  and _77891_ (_27293_, _27291_, _10290_);
  and _77892_ (_27294_, _27293_, _27279_);
  nor _77893_ (_27295_, _27268_, _10290_);
  or _77894_ (_27296_, _27295_, _05833_);
  or _77895_ (_27297_, _27296_, _27294_);
  and _77896_ (_27298_, _27297_, _27278_);
  or _77897_ (_27299_, _27298_, _04438_);
  nand _77898_ (_27300_, _27268_, _04438_);
  and _77899_ (_27301_, _27300_, _04444_);
  and _77900_ (_27302_, _27301_, _27299_);
  and _77901_ (_27304_, _10206_, _10203_);
  nor _77902_ (_27305_, _27304_, _10207_);
  or _77903_ (_27306_, _27305_, _10261_);
  and _77904_ (_27307_, _27306_, _03570_);
  nand _77905_ (_27308_, _10261_, _10179_);
  and _77906_ (_27309_, _27308_, _27307_);
  or _77907_ (_27310_, _27309_, _27302_);
  and _77908_ (_27311_, _27310_, _10255_);
  nor _77909_ (_27312_, _27268_, _10255_);
  or _77910_ (_27313_, _27312_, _03516_);
  or _77911_ (_27315_, _27313_, _27311_);
  nand _77912_ (_27316_, _10016_, _03516_);
  and _77913_ (_27317_, _27316_, _03203_);
  and _77914_ (_27318_, _27317_, _27315_);
  nor _77915_ (_27319_, _06195_, _03203_);
  or _77916_ (_27320_, _27319_, _03568_);
  or _77917_ (_27321_, _27320_, _27318_);
  nand _77918_ (_27322_, _10016_, _03568_);
  and _77919_ (_27323_, _27322_, _27321_);
  or _77920_ (_27324_, _27323_, _26212_);
  and _77921_ (_27326_, _27324_, _27274_);
  or _77922_ (_27327_, _27326_, _03575_);
  nand _77923_ (_27328_, _10016_, _03575_);
  and _77924_ (_27329_, _27328_, _10316_);
  and _77925_ (_27330_, _27329_, _27327_);
  nor _77926_ (_27331_, _27268_, _10316_);
  or _77927_ (_27332_, _27331_, _03512_);
  or _77928_ (_27333_, _27332_, _27330_);
  and _77929_ (_27334_, _27333_, _27273_);
  or _77930_ (_27335_, _27334_, _10249_);
  nand _77931_ (_27337_, _06195_, _10249_);
  and _77932_ (_27338_, _27337_, _04887_);
  and _77933_ (_27339_, _27338_, _27335_);
  nand _77934_ (_27340_, _10015_, _03511_);
  nand _77935_ (_27341_, _27340_, _10325_);
  or _77936_ (_27342_, _27341_, _27339_);
  and _77937_ (_27343_, _10360_, _10178_);
  not _77938_ (_27344_, _27305_);
  nor _77939_ (_27345_, _27344_, _10360_);
  or _77940_ (_27346_, _27345_, _27343_);
  or _77941_ (_27348_, _27346_, _10325_);
  and _77942_ (_27349_, _27348_, _27342_);
  or _77943_ (_27350_, _27349_, _27272_);
  and _77944_ (_27351_, _10178_, _10116_);
  nor _77945_ (_27352_, _27344_, _10116_);
  or _77946_ (_27353_, _27352_, _27351_);
  or _77947_ (_27354_, _27353_, _10328_);
  and _77948_ (_27355_, _27354_, _27350_);
  or _77949_ (_27356_, _27355_, _03527_);
  nor _77950_ (_27357_, _27344_, _10382_);
  and _77951_ (_27359_, _10382_, _10178_);
  or _77952_ (_27360_, _27359_, _03998_);
  or _77953_ (_27361_, _27360_, _27357_);
  and _77954_ (_27362_, _27361_, _10085_);
  and _77955_ (_27363_, _27362_, _27356_);
  or _77956_ (_27364_, _27305_, _10398_);
  nand _77957_ (_27365_, _10398_, _10179_);
  and _77958_ (_27366_, _27365_, _03638_);
  and _77959_ (_27367_, _27366_, _27364_);
  or _77960_ (_27368_, _27367_, _10083_);
  or _77961_ (_27370_, _27368_, _27363_);
  and _77962_ (_27371_, _27370_, _27271_);
  or _77963_ (_27372_, _27371_, _03505_);
  nand _77964_ (_27373_, _10016_, _03505_);
  and _77965_ (_27374_, _27373_, _03200_);
  and _77966_ (_27375_, _27374_, _27372_);
  nor _77967_ (_27376_, _06195_, _03200_);
  or _77968_ (_27377_, _27376_, _26282_);
  or _77969_ (_27378_, _27377_, _27375_);
  and _77970_ (_27379_, _27378_, _27264_);
  or _77971_ (_27381_, _27379_, _25991_);
  or _77972_ (_27382_, _27267_, _10415_);
  and _77973_ (_27383_, _27382_, _10419_);
  and _77974_ (_27384_, _27383_, _27381_);
  and _77975_ (_27385_, _10015_, _03607_);
  or _77976_ (_27386_, _27385_, _10420_);
  or _77977_ (_27387_, _27386_, _27384_);
  nand _77978_ (_27388_, _06195_, _10420_);
  and _77979_ (_27389_, _27388_, _27387_);
  or _77980_ (_27390_, _27389_, _03606_);
  nand _77981_ (_27392_, _10016_, _03606_);
  and _77982_ (_27393_, _27392_, _10426_);
  and _77983_ (_27394_, _27393_, _27390_);
  nor _77984_ (_27395_, _27268_, _10426_);
  or _77985_ (_27396_, _27395_, _10431_);
  or _77986_ (_27397_, _27396_, _27394_);
  or _77987_ (_27398_, _10015_, _10430_);
  and _77988_ (_27399_, _27398_, _03254_);
  and _77989_ (_27400_, _27399_, _27397_);
  nor _77990_ (_27401_, _27268_, _03254_);
  or _77991_ (_27403_, _27401_, _03499_);
  or _77992_ (_27404_, _27403_, _27400_);
  nand _77993_ (_27405_, _10016_, _03499_);
  and _77994_ (_27406_, _27405_, _27404_);
  or _77995_ (_27407_, _27406_, _03223_);
  nand _77996_ (_27408_, _06195_, _03223_);
  and _77997_ (_27409_, _27408_, _09755_);
  and _77998_ (_27410_, _27409_, _27407_);
  nand _77999_ (_27411_, _10178_, _03632_);
  nand _78000_ (_27412_, _27411_, _03493_);
  or _78001_ (_27414_, _27412_, _27410_);
  or _78002_ (_27415_, _10015_, _03493_);
  and _78003_ (_27416_, _27415_, _03474_);
  and _78004_ (_27417_, _27416_, _27414_);
  nand _78005_ (_27418_, _10178_, _03221_);
  nand _78006_ (_27419_, _27418_, _10081_);
  or _78007_ (_27420_, _27419_, _27417_);
  not _78008_ (_27421_, _03745_);
  or _78009_ (_27422_, _27267_, _10081_);
  and _78010_ (_27423_, _27422_, _27421_);
  and _78011_ (_27425_, _27423_, _27420_);
  and _78012_ (_27426_, _10015_, _03745_);
  or _78013_ (_27427_, _27426_, _03187_);
  or _78014_ (_27428_, _27427_, _27425_);
  nand _78015_ (_27429_, _06195_, _03187_);
  and _78016_ (_27430_, _27429_, _10459_);
  and _78017_ (_27431_, _27430_, _27428_);
  and _78018_ (_27432_, _27259_, _10458_);
  or _78019_ (_27433_, _27432_, _06055_);
  or _78020_ (_27434_, _27433_, _27431_);
  or _78021_ (_27436_, _10015_, _05775_);
  and _78022_ (_27437_, _27436_, _03438_);
  and _78023_ (_27438_, _27437_, _27434_);
  and _78024_ (_27439_, _10178_, _03437_);
  or _78025_ (_27440_, _27439_, _08385_);
  or _78026_ (_27441_, _27440_, _27438_);
  and _78027_ (_27442_, _10016_, _08385_);
  nor _78028_ (_27443_, _27442_, _10472_);
  and _78029_ (_27444_, _27443_, _27441_);
  nor _78030_ (_27445_, _10490_, _10488_);
  nor _78031_ (_27447_, _27445_, _10491_);
  and _78032_ (_27448_, _27447_, _10472_);
  or _78033_ (_27449_, _27448_, _03744_);
  or _78034_ (_27450_, _27449_, _27444_);
  nand _78035_ (_27451_, _10016_, _03744_);
  and _78036_ (_27452_, _27451_, _27450_);
  or _78037_ (_27453_, _27452_, _03189_);
  nand _78038_ (_27454_, _06195_, _03189_);
  and _78039_ (_27455_, _27454_, _10515_);
  and _78040_ (_27456_, _27455_, _27453_);
  or _78041_ (_27458_, _27259_, _08698_);
  nand _78042_ (_27459_, _10016_, _08698_);
  and _78043_ (_27460_, _27459_, _10076_);
  and _78044_ (_27461_, _27460_, _27458_);
  or _78045_ (_27462_, _27461_, _27456_);
  and _78046_ (_27463_, _27462_, _10520_);
  nor _78047_ (_27464_, _27268_, _10520_);
  or _78048_ (_27465_, _27464_, _10524_);
  or _78049_ (_27466_, _27465_, _27463_);
  or _78050_ (_27467_, _10523_, _10015_);
  and _78051_ (_27469_, _27467_, _04499_);
  and _78052_ (_27470_, _27469_, _27466_);
  and _78053_ (_27471_, _10178_, _03636_);
  or _78054_ (_27472_, _27471_, _03769_);
  or _78055_ (_27473_, _27472_, _27470_);
  nand _78056_ (_27474_, _10016_, _03769_);
  and _78057_ (_27475_, _27474_, _27473_);
  or _78058_ (_27476_, _27475_, _03194_);
  nand _78059_ (_27477_, _06195_, _03194_);
  and _78060_ (_27478_, _27477_, _10535_);
  and _78061_ (_27480_, _27478_, _27476_);
  or _78062_ (_27481_, _27259_, _10077_);
  or _78063_ (_27482_, _10015_, _08698_);
  and _78064_ (_27483_, _27482_, _10534_);
  and _78065_ (_27484_, _27483_, _27481_);
  or _78066_ (_27485_, _27484_, _27480_);
  and _78067_ (_27486_, _27485_, _10546_);
  and _78068_ (_27487_, _27267_, _10545_);
  or _78069_ (_27488_, _27487_, _10549_);
  or _78070_ (_27489_, _27488_, _27486_);
  or _78071_ (_27491_, _10015_, _10548_);
  and _78072_ (_27492_, _27491_, _05769_);
  and _78073_ (_27493_, _27492_, _27489_);
  and _78074_ (_27494_, _10178_, _03754_);
  or _78075_ (_27495_, _27494_, _03752_);
  or _78076_ (_27496_, _27495_, _27493_);
  nand _78077_ (_27497_, _10016_, _03752_);
  and _78078_ (_27498_, _27497_, _27496_);
  or _78079_ (_27499_, _27498_, _03192_);
  nand _78080_ (_27500_, _06195_, _03192_);
  and _78081_ (_27502_, _27500_, _09959_);
  and _78082_ (_27503_, _27502_, _27499_);
  or _78083_ (_27504_, _27503_, _27263_);
  and _78084_ (_27505_, _27504_, _09956_);
  nor _78085_ (_27506_, _27268_, _09956_);
  or _78086_ (_27507_, _27506_, _08479_);
  or _78087_ (_27508_, _27507_, _27505_);
  or _78088_ (_27509_, _10015_, _08478_);
  and _78089_ (_27510_, _27509_, _03759_);
  and _78090_ (_27511_, _27510_, _27508_);
  and _78091_ (_27513_, _10178_, _03758_);
  or _78092_ (_27514_, _27513_, _03760_);
  or _78093_ (_27515_, _27514_, _27511_);
  nand _78094_ (_27516_, _10016_, _03760_);
  and _78095_ (_27517_, _27516_, _27515_);
  or _78096_ (_27518_, _27517_, _03183_);
  nand _78097_ (_27519_, _06195_, _03183_);
  and _78098_ (_27520_, _27519_, _10577_);
  and _78099_ (_27521_, _27520_, _27518_);
  or _78100_ (_27522_, _27259_, _07888_);
  or _78101_ (_27523_, _10015_, \oc8051_golden_model_1.PSW [7]);
  and _78102_ (_27524_, _27523_, _10576_);
  and _78103_ (_27525_, _27524_, _27522_);
  or _78104_ (_27526_, _27525_, _27521_);
  and _78105_ (_27527_, _27526_, _09951_);
  nor _78106_ (_27528_, _27268_, _09951_);
  or _78107_ (_27529_, _27528_, _08525_);
  or _78108_ (_27530_, _27529_, _27527_);
  or _78109_ (_27531_, _10015_, _08524_);
  and _78110_ (_27532_, _27531_, _08556_);
  and _78111_ (_27535_, _27532_, _27530_);
  and _78112_ (_27536_, _27267_, _08555_);
  or _78113_ (_27537_, _27536_, _03775_);
  or _78114_ (_27538_, _27537_, _27535_);
  or _78115_ (_27539_, _06722_, _11403_);
  and _78116_ (_27540_, _27539_, _27538_);
  or _78117_ (_27541_, _27540_, _03179_);
  nand _78118_ (_27542_, _06195_, _03179_);
  and _78119_ (_27543_, _27542_, _10599_);
  and _78120_ (_27544_, _27543_, _27541_);
  nor _78121_ (_27546_, _10794_, _10179_);
  and _78122_ (_27547_, _27305_, _10794_);
  or _78123_ (_27548_, _27547_, _27546_);
  and _78124_ (_27549_, _27548_, _03627_);
  or _78125_ (_27550_, _27549_, _27544_);
  and _78126_ (_27551_, _27550_, _09949_);
  nor _78127_ (_27552_, _27268_, _09949_);
  or _78128_ (_27553_, _27552_, _09937_);
  or _78129_ (_27554_, _27553_, _27551_);
  or _78130_ (_27555_, _10015_, _09936_);
  and _78131_ (_27557_, _27555_, _10803_);
  and _78132_ (_27558_, _27557_, _27554_);
  and _78133_ (_27559_, _27267_, _07729_);
  or _78134_ (_27560_, _27559_, _03522_);
  or _78135_ (_27561_, _27560_, _27558_);
  or _78136_ (_27562_, _06722_, _03523_);
  and _78137_ (_27563_, _27562_, _25887_);
  and _78138_ (_27564_, _27563_, _27561_);
  nor _78139_ (_27565_, _06195_, _25887_);
  or _78140_ (_27566_, _27565_, _03628_);
  or _78141_ (_27568_, _27566_, _27564_);
  nand _78142_ (_27569_, _10794_, _10179_);
  or _78143_ (_27570_, _27305_, _10794_);
  and _78144_ (_27571_, _27570_, _27569_);
  or _78145_ (_27572_, _27571_, _03791_);
  and _78146_ (_27573_, _27572_, _10821_);
  and _78147_ (_27574_, _27573_, _27568_);
  nor _78148_ (_27575_, _27268_, _10821_);
  or _78149_ (_27576_, _27575_, _03790_);
  or _78150_ (_27577_, _27576_, _27574_);
  nand _78151_ (_27579_, _10016_, _03790_);
  and _78152_ (_27580_, _27579_, _10828_);
  and _78153_ (_27581_, _27580_, _27577_);
  nor _78154_ (_27582_, _27268_, _10828_);
  or _78155_ (_27583_, _27582_, _04947_);
  or _78156_ (_27584_, _27583_, _27581_);
  and _78157_ (_27585_, _27584_, _27257_);
  or _78158_ (_27586_, _27585_, _03151_);
  or _78159_ (_27587_, _27571_, _03152_);
  and _78160_ (_27588_, _27587_, _10844_);
  and _78161_ (_27590_, _27588_, _27586_);
  nor _78162_ (_27591_, _27268_, _10844_);
  or _78163_ (_27592_, _27591_, _03520_);
  or _78164_ (_27593_, _27592_, _27590_);
  nand _78165_ (_27594_, _10016_, _03520_);
  and _78166_ (_27595_, _27594_, _10851_);
  and _78167_ (_27596_, _27595_, _27593_);
  nor _78168_ (_27597_, _27268_, _10851_);
  or _78169_ (_27598_, _27597_, _25883_);
  or _78170_ (_27599_, _27598_, _27596_);
  nand _78171_ (_27601_, _25883_, _06195_);
  and _78172_ (_27602_, _27601_, _10863_);
  and _78173_ (_27603_, _27602_, _27599_);
  and _78174_ (_27604_, _27267_, _10862_);
  or _78175_ (_27605_, _27604_, _27603_);
  or _78176_ (_27606_, _27605_, _42967_);
  or _78177_ (_27607_, _42963_, \oc8051_golden_model_1.PC [4]);
  and _78178_ (_27608_, _27607_, _41755_);
  and _78179_ (_43331_, _27608_, _27606_);
  nor _78180_ (_27609_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor _78181_ (_27611_, _10010_, _02887_);
  nor _78182_ (_27612_, _27611_, _27609_);
  and _78183_ (_27613_, _27612_, _10862_);
  and _78184_ (_27614_, _10010_, _03520_);
  and _78185_ (_27615_, _10010_, _03790_);
  nor _78186_ (_27616_, _27612_, _09949_);
  nor _78187_ (_27617_, _27612_, _09951_);
  nor _78188_ (_27618_, _27612_, _09956_);
  not _78189_ (_27619_, _27612_);
  and _78190_ (_27620_, _27619_, _10545_);
  nor _78191_ (_27622_, _27612_, _10520_);
  and _78192_ (_27623_, _10011_, _03744_);
  and _78193_ (_27624_, _10011_, _03499_);
  nor _78194_ (_27625_, _26281_, _10010_);
  and _78195_ (_27626_, _27619_, _10083_);
  or _78196_ (_27627_, _10176_, _10175_);
  and _78197_ (_27628_, _27627_, _10208_);
  nor _78198_ (_27629_, _27627_, _10208_);
  or _78199_ (_27630_, _27629_, _27628_);
  nor _78200_ (_27631_, _27630_, _10116_);
  and _78201_ (_27633_, _10173_, _10116_);
  nor _78202_ (_27634_, _27633_, _27631_);
  nor _78203_ (_27635_, _27634_, _10328_);
  and _78204_ (_27636_, _10261_, _10173_);
  nor _78205_ (_27637_, _27630_, _10261_);
  or _78206_ (_27638_, _27637_, _27636_);
  or _78207_ (_27639_, _27638_, _04444_);
  and _78208_ (_27640_, _10269_, _10010_);
  or _78209_ (_27641_, _10013_, _10012_);
  not _78210_ (_27642_, _27641_);
  nor _78211_ (_27644_, _27642_, _10038_);
  and _78212_ (_27645_, _27642_, _10038_);
  nor _78213_ (_27646_, _27645_, _27644_);
  nor _78214_ (_27647_, _27646_, _10269_);
  or _78215_ (_27648_, _27647_, _27640_);
  nor _78216_ (_27649_, _27648_, _05831_);
  nor _78217_ (_27650_, _27612_, _10290_);
  nor _78218_ (_27651_, _27612_, _25905_);
  not _78219_ (_27652_, _27651_);
  not _78220_ (_27653_, \oc8051_golden_model_1.PC [5]);
  and _78221_ (_27655_, _26180_, _27653_);
  and _78222_ (_27656_, _10011_, _04426_);
  nor _78223_ (_27657_, _27656_, _03923_);
  not _78224_ (_27658_, _27657_);
  nor _78225_ (_27659_, _27658_, _27655_);
  and _78226_ (_27660_, _27659_, _27652_);
  not _78227_ (_27661_, _10290_);
  nor _78228_ (_27662_, _06164_, _04762_);
  or _78229_ (_27663_, _27662_, _27661_);
  nor _78230_ (_27664_, _27663_, _27660_);
  nor _78231_ (_27666_, _27664_, _27650_);
  nor _78232_ (_27667_, _27666_, _05833_);
  or _78233_ (_27668_, _27667_, _04438_);
  nor _78234_ (_27669_, _27668_, _27649_);
  and _78235_ (_27670_, _27612_, _04438_);
  or _78236_ (_27671_, _27670_, _03570_);
  or _78237_ (_27672_, _27671_, _27669_);
  and _78238_ (_27673_, _27672_, _27639_);
  nor _78239_ (_27674_, _27673_, _10256_);
  nor _78240_ (_27675_, _27612_, _10255_);
  nor _78241_ (_27677_, _27675_, _03516_);
  not _78242_ (_27678_, _27677_);
  nor _78243_ (_27679_, _27678_, _27674_);
  and _78244_ (_27680_, _10010_, _03516_);
  nor _78245_ (_27681_, _27680_, _27679_);
  or _78246_ (_27682_, _27681_, _04746_);
  or _78247_ (_27683_, _06164_, _03203_);
  and _78248_ (_27684_, _27683_, _27682_);
  or _78249_ (_27685_, _27684_, _03568_);
  and _78250_ (_27686_, _10010_, _03568_);
  nor _78251_ (_27688_, _27686_, _26212_);
  nand _78252_ (_27689_, _27688_, _27685_);
  nor _78253_ (_27690_, _27612_, _10307_);
  nor _78254_ (_27691_, _27690_, _03575_);
  nand _78255_ (_27692_, _27691_, _27689_);
  and _78256_ (_27693_, _10010_, _03575_);
  nor _78257_ (_27694_, _27693_, _26220_);
  nand _78258_ (_27695_, _27694_, _27692_);
  nor _78259_ (_27696_, _27612_, _10316_);
  nor _78260_ (_27697_, _27696_, _03512_);
  nand _78261_ (_27699_, _27697_, _27695_);
  and _78262_ (_27700_, _10010_, _03512_);
  nor _78263_ (_27701_, _27700_, _10249_);
  nand _78264_ (_27702_, _27701_, _27699_);
  and _78265_ (_27703_, _06164_, _10249_);
  nor _78266_ (_27704_, _27703_, _03511_);
  nand _78267_ (_27705_, _27704_, _27702_);
  and _78268_ (_27706_, _10010_, _03511_);
  nor _78269_ (_27707_, _27706_, _10326_);
  nand _78270_ (_27708_, _27707_, _27705_);
  and _78271_ (_27710_, _10360_, _10173_);
  nor _78272_ (_27711_, _27630_, _10360_);
  or _78273_ (_27712_, _27711_, _27710_);
  nor _78274_ (_27713_, _27712_, _10325_);
  nor _78275_ (_27714_, _27713_, _03657_);
  nand _78276_ (_27715_, _27714_, _27708_);
  nand _78277_ (_27716_, _27715_, _03998_);
  or _78278_ (_27717_, _27716_, _27635_);
  nor _78279_ (_27718_, _27630_, _10382_);
  not _78280_ (_27719_, _27718_);
  and _78281_ (_27721_, _10382_, _10173_);
  nor _78282_ (_27722_, _27721_, _03998_);
  and _78283_ (_27723_, _27722_, _27719_);
  nor _78284_ (_27724_, _27723_, _03638_);
  nand _78285_ (_27725_, _27724_, _27717_);
  and _78286_ (_27726_, _27630_, _10399_);
  and _78287_ (_27727_, _10398_, _10174_);
  or _78288_ (_27728_, _27727_, _10085_);
  or _78289_ (_27729_, _27728_, _27726_);
  and _78290_ (_27730_, _27729_, _10084_);
  and _78291_ (_27732_, _27730_, _27725_);
  or _78292_ (_27733_, _27732_, _27626_);
  nand _78293_ (_27734_, _27733_, _03506_);
  and _78294_ (_27735_, _10011_, _03505_);
  nor _78295_ (_27736_, _27735_, _04743_);
  nand _78296_ (_27737_, _27736_, _27734_);
  nor _78297_ (_27738_, _06164_, _03200_);
  nor _78298_ (_27739_, _27738_, _26282_);
  and _78299_ (_27740_, _27739_, _27737_);
  or _78300_ (_27741_, _27740_, _27625_);
  nand _78301_ (_27743_, _27741_, _10415_);
  nor _78302_ (_27744_, _27612_, _10415_);
  nor _78303_ (_27745_, _27744_, _03607_);
  nand _78304_ (_27746_, _27745_, _27743_);
  and _78305_ (_27747_, _10010_, _03607_);
  nor _78306_ (_27748_, _27747_, _10420_);
  nand _78307_ (_27749_, _27748_, _27746_);
  and _78308_ (_27750_, _06164_, _10420_);
  nor _78309_ (_27751_, _27750_, _03606_);
  nand _78310_ (_27752_, _27751_, _27749_);
  and _78311_ (_27754_, _10010_, _03606_);
  nor _78312_ (_27755_, _27754_, _26302_);
  and _78313_ (_27756_, _27755_, _27752_);
  nor _78314_ (_27757_, _27612_, _10426_);
  or _78315_ (_27758_, _27757_, _27756_);
  nand _78316_ (_27759_, _27758_, _10430_);
  nor _78317_ (_27760_, _10010_, _10430_);
  nor _78318_ (_27761_, _27760_, _03311_);
  nand _78319_ (_27762_, _27761_, _27759_);
  nor _78320_ (_27763_, _27619_, _03254_);
  nor _78321_ (_27765_, _27763_, _03499_);
  and _78322_ (_27766_, _27765_, _27762_);
  or _78323_ (_27767_, _27766_, _27624_);
  nand _78324_ (_27768_, _27767_, _04853_);
  and _78325_ (_27769_, _06164_, _03223_);
  nor _78326_ (_27770_, _27769_, _03632_);
  nand _78327_ (_27771_, _27770_, _27768_);
  and _78328_ (_27772_, _10173_, _03632_);
  nor _78329_ (_27773_, _27772_, _26322_);
  nand _78330_ (_27774_, _27773_, _27771_);
  nor _78331_ (_27776_, _10010_, _03493_);
  nor _78332_ (_27777_, _27776_, _03221_);
  nand _78333_ (_27778_, _27777_, _27774_);
  and _78334_ (_27779_, _10173_, _03221_);
  nor _78335_ (_27780_, _27779_, _26330_);
  nand _78336_ (_27781_, _27780_, _27778_);
  nor _78337_ (_27782_, _27612_, _10081_);
  nor _78338_ (_27783_, _27782_, _03745_);
  and _78339_ (_27784_, _27783_, _27781_);
  and _78340_ (_27785_, _10010_, _03745_);
  or _78341_ (_27787_, _27785_, _03187_);
  or _78342_ (_27788_, _27787_, _27784_);
  and _78343_ (_27789_, _06164_, _03187_);
  nor _78344_ (_27790_, _27789_, _10458_);
  nand _78345_ (_27791_, _27790_, _27788_);
  nor _78346_ (_27792_, _27646_, _10459_);
  nor _78347_ (_27793_, _27792_, _06055_);
  nand _78348_ (_27794_, _27793_, _27791_);
  nor _78349_ (_27795_, _10010_, _05775_);
  nor _78350_ (_27796_, _27795_, _03437_);
  nand _78351_ (_27798_, _27796_, _27794_);
  and _78352_ (_27799_, _10173_, _03437_);
  nor _78353_ (_27800_, _27799_, _08385_);
  nand _78354_ (_27801_, _27800_, _27798_);
  and _78355_ (_27802_, _10011_, _08385_);
  nor _78356_ (_27803_, _27802_, _10472_);
  nand _78357_ (_27804_, _27803_, _27801_);
  and _78358_ (_27805_, _10492_, _10485_);
  not _78359_ (_27806_, _27805_);
  nor _78360_ (_27807_, _10493_, _25897_);
  and _78361_ (_27808_, _27807_, _27806_);
  nor _78362_ (_27809_, _27808_, _03744_);
  and _78363_ (_27810_, _27809_, _27804_);
  or _78364_ (_27811_, _27810_, _27623_);
  nand _78365_ (_27812_, _27811_, _11376_);
  and _78366_ (_27813_, _06164_, _03189_);
  nor _78367_ (_27814_, _27813_, _10076_);
  nand _78368_ (_27815_, _27814_, _27812_);
  and _78369_ (_27816_, _10010_, _08698_);
  nor _78370_ (_27817_, _27646_, _08698_);
  or _78371_ (_27820_, _27817_, _27816_);
  and _78372_ (_27821_, _27820_, _10076_);
  nor _78373_ (_27822_, _27821_, _26754_);
  and _78374_ (_27823_, _27822_, _27815_);
  or _78375_ (_27824_, _27823_, _27622_);
  nand _78376_ (_27825_, _27824_, _10523_);
  nor _78377_ (_27826_, _10523_, _10010_);
  nor _78378_ (_27827_, _27826_, _03636_);
  and _78379_ (_27828_, _27827_, _27825_);
  and _78380_ (_27829_, _10173_, _03636_);
  or _78381_ (_27831_, _27829_, _03769_);
  nor _78382_ (_27832_, _27831_, _27828_);
  and _78383_ (_27833_, _10011_, _03769_);
  or _78384_ (_27834_, _27833_, _27832_);
  nand _78385_ (_27835_, _27834_, _25894_);
  and _78386_ (_27836_, _06164_, _03194_);
  nor _78387_ (_27837_, _27836_, _10534_);
  nand _78388_ (_27838_, _27837_, _27835_);
  and _78389_ (_27839_, _27646_, _08698_);
  nor _78390_ (_27840_, _10010_, _08698_);
  nor _78391_ (_27842_, _27840_, _10535_);
  not _78392_ (_27843_, _27842_);
  nor _78393_ (_27844_, _27843_, _27839_);
  nor _78394_ (_27845_, _27844_, _10545_);
  and _78395_ (_27846_, _27845_, _27838_);
  or _78396_ (_27847_, _27846_, _27620_);
  nand _78397_ (_27848_, _27847_, _10548_);
  nor _78398_ (_27849_, _10010_, _10548_);
  nor _78399_ (_27850_, _27849_, _04504_);
  nand _78400_ (_27851_, _27850_, _27848_);
  and _78401_ (_27853_, _10173_, _03754_);
  nor _78402_ (_27854_, _27853_, _03752_);
  and _78403_ (_27855_, _27854_, _27851_);
  and _78404_ (_27856_, _10011_, _03752_);
  or _78405_ (_27857_, _27856_, _27855_);
  nand _78406_ (_27858_, _27857_, _25891_);
  and _78407_ (_27859_, _06164_, _03192_);
  nor _78408_ (_27860_, _27859_, _09958_);
  nand _78409_ (_27861_, _27860_, _27858_);
  and _78410_ (_27862_, _27646_, _07888_);
  nor _78411_ (_27864_, _10010_, _07888_);
  nor _78412_ (_27865_, _27864_, _09959_);
  not _78413_ (_27866_, _27865_);
  nor _78414_ (_27867_, _27866_, _27862_);
  nor _78415_ (_27868_, _27867_, _10560_);
  and _78416_ (_27869_, _27868_, _27861_);
  or _78417_ (_27870_, _27869_, _27618_);
  nand _78418_ (_27871_, _27870_, _08478_);
  nor _78419_ (_27872_, _10010_, _08478_);
  nor _78420_ (_27873_, _27872_, _03758_);
  and _78421_ (_27875_, _27873_, _27871_);
  and _78422_ (_27876_, _10173_, _03758_);
  or _78423_ (_27877_, _27876_, _03760_);
  nor _78424_ (_27878_, _27877_, _27875_);
  and _78425_ (_27879_, _10011_, _03760_);
  or _78426_ (_27880_, _27879_, _27878_);
  nand _78427_ (_27881_, _27880_, _26082_);
  and _78428_ (_27882_, _06164_, _03183_);
  nor _78429_ (_27883_, _27882_, _10576_);
  nand _78430_ (_27884_, _27883_, _27881_);
  and _78431_ (_27886_, _27646_, \oc8051_golden_model_1.PSW [7]);
  nor _78432_ (_27887_, _10010_, \oc8051_golden_model_1.PSW [7]);
  nor _78433_ (_27888_, _27887_, _10577_);
  not _78434_ (_27889_, _27888_);
  nor _78435_ (_27890_, _27889_, _27886_);
  nor _78436_ (_27891_, _27890_, _10581_);
  and _78437_ (_27892_, _27891_, _27884_);
  or _78438_ (_27893_, _27892_, _27617_);
  nand _78439_ (_27894_, _27893_, _08524_);
  nor _78440_ (_27895_, _10010_, _08524_);
  nor _78441_ (_27897_, _27895_, _08555_);
  and _78442_ (_27898_, _27897_, _27894_);
  and _78443_ (_27899_, _27612_, _08555_);
  or _78444_ (_27900_, _27899_, _03775_);
  nor _78445_ (_27901_, _27900_, _27898_);
  and _78446_ (_27902_, _06616_, _03775_);
  or _78447_ (_27903_, _27902_, _27901_);
  nand _78448_ (_27904_, _27903_, _06328_);
  and _78449_ (_27905_, _06164_, _03179_);
  nor _78450_ (_27906_, _27905_, _03627_);
  nand _78451_ (_27908_, _27906_, _27904_);
  and _78452_ (_27909_, _27630_, _10794_);
  nor _78453_ (_27910_, _10794_, _10173_);
  or _78454_ (_27911_, _27910_, _10599_);
  or _78455_ (_27912_, _27911_, _27909_);
  and _78456_ (_27913_, _27912_, _09949_);
  and _78457_ (_27914_, _27913_, _27908_);
  or _78458_ (_27915_, _27914_, _27616_);
  nand _78459_ (_27916_, _27915_, _09936_);
  nor _78460_ (_27917_, _10010_, _09936_);
  nor _78461_ (_27919_, _27917_, _07729_);
  and _78462_ (_27920_, _27919_, _27916_);
  and _78463_ (_27921_, _27612_, _07729_);
  or _78464_ (_27922_, _27921_, _03522_);
  nor _78465_ (_27923_, _27922_, _27920_);
  and _78466_ (_27924_, _06616_, _03522_);
  or _78467_ (_27925_, _27924_, _27923_);
  nand _78468_ (_27926_, _27925_, _25887_);
  and _78469_ (_27927_, _06164_, _03172_);
  nor _78470_ (_27928_, _27927_, _03628_);
  nand _78471_ (_27930_, _27928_, _27926_);
  and _78472_ (_27931_, _10794_, _10173_);
  nor _78473_ (_27932_, _27630_, _10794_);
  or _78474_ (_27933_, _27932_, _27931_);
  and _78475_ (_27934_, _27933_, _03628_);
  nor _78476_ (_27935_, _27934_, _10822_);
  nand _78477_ (_27936_, _27935_, _27930_);
  nor _78478_ (_27937_, _27612_, _10821_);
  nor _78479_ (_27938_, _27937_, _03790_);
  and _78480_ (_27939_, _27938_, _27936_);
  or _78481_ (_27941_, _27939_, _27615_);
  nand _78482_ (_27942_, _27941_, _10828_);
  nor _78483_ (_27943_, _27619_, _10828_);
  nor _78484_ (_27944_, _27943_, _04947_);
  nand _78485_ (_27945_, _27944_, _27942_);
  and _78486_ (_27946_, _06164_, _04947_);
  nor _78487_ (_27947_, _27946_, _03151_);
  nand _78488_ (_27948_, _27947_, _27945_);
  and _78489_ (_27949_, _27933_, _03151_);
  nor _78490_ (_27950_, _27949_, _10845_);
  nand _78491_ (_27952_, _27950_, _27948_);
  nor _78492_ (_27953_, _27612_, _10844_);
  nor _78493_ (_27954_, _27953_, _03520_);
  and _78494_ (_27955_, _27954_, _27952_);
  or _78495_ (_27956_, _27955_, _27614_);
  nand _78496_ (_27957_, _27956_, _10851_);
  nor _78497_ (_27958_, _27619_, _10851_);
  nor _78498_ (_27959_, _27958_, _25883_);
  nand _78499_ (_27960_, _27959_, _27957_);
  and _78500_ (_27961_, _25883_, _06164_);
  nor _78501_ (_27963_, _27961_, _10862_);
  and _78502_ (_27964_, _27963_, _27960_);
  or _78503_ (_27965_, _27964_, _27613_);
  or _78504_ (_27966_, _27965_, _42967_);
  or _78505_ (_27967_, _42963_, \oc8051_golden_model_1.PC [5]);
  and _78506_ (_27968_, _27967_, _41755_);
  and _78507_ (_43334_, _27968_, _27966_);
  nand _78508_ (_27969_, _06132_, _04947_);
  and _78509_ (_27970_, _05836_, _09938_);
  nor _78510_ (_27971_, _27970_, \oc8051_golden_model_1.PC [6]);
  nor _78511_ (_27973_, _27971_, _09939_);
  not _78512_ (_27974_, _27973_);
  nand _78513_ (_27975_, _27974_, _07729_);
  nand _78514_ (_27976_, _10166_, _03758_);
  nand _78515_ (_27977_, _10166_, _03636_);
  nor _78516_ (_27978_, _10041_, _10007_);
  nor _78517_ (_27979_, _27978_, _10042_);
  and _78518_ (_27980_, _27979_, _10458_);
  nand _78519_ (_27981_, _27974_, _10083_);
  and _78520_ (_27982_, _10210_, _10170_);
  nor _78521_ (_27984_, _27982_, _10211_);
  or _78522_ (_27985_, _27984_, _10116_);
  nand _78523_ (_27986_, _10166_, _10116_);
  and _78524_ (_27987_, _27986_, _27985_);
  or _78525_ (_27988_, _27987_, _10328_);
  or _78526_ (_27989_, _27973_, _10303_);
  and _78527_ (_27990_, _10261_, _10165_);
  not _78528_ (_27991_, _10261_);
  and _78529_ (_27992_, _27984_, _27991_);
  or _78530_ (_27993_, _27992_, _04444_);
  or _78531_ (_27995_, _27993_, _27990_);
  nand _78532_ (_27996_, _06132_, _03923_);
  and _78533_ (_27997_, _10003_, _04426_);
  and _78534_ (_27998_, _04427_, \oc8051_golden_model_1.PC [6]);
  and _78535_ (_27999_, _27998_, _10278_);
  or _78536_ (_28000_, _27999_, _27997_);
  and _78537_ (_28001_, _28000_, _26578_);
  nor _78538_ (_28002_, _27974_, _25905_);
  or _78539_ (_28003_, _28002_, _28001_);
  and _78540_ (_28004_, _28003_, _10290_);
  or _78541_ (_28006_, _28004_, _03923_);
  and _78542_ (_28007_, _28006_, _27996_);
  nor _78543_ (_28008_, _27974_, _10290_);
  or _78544_ (_28009_, _28008_, _05833_);
  or _78545_ (_28010_, _28009_, _28007_);
  and _78546_ (_28011_, _27979_, _10271_);
  and _78547_ (_28012_, _10269_, _10003_);
  or _78548_ (_28013_, _28012_, _05831_);
  or _78549_ (_28014_, _28013_, _28011_);
  and _78550_ (_28015_, _28014_, _28010_);
  or _78551_ (_28017_, _28015_, _10297_);
  and _78552_ (_28018_, _28017_, _27995_);
  or _78553_ (_28019_, _28018_, _10256_);
  and _78554_ (_28020_, _28019_, _27989_);
  or _78555_ (_28021_, _28020_, _03516_);
  nand _78556_ (_28022_, _10004_, _03516_);
  and _78557_ (_28023_, _28022_, _03203_);
  and _78558_ (_28024_, _28023_, _28021_);
  nor _78559_ (_28025_, _06132_, _03203_);
  or _78560_ (_28026_, _28025_, _03568_);
  or _78561_ (_28028_, _28026_, _28024_);
  nand _78562_ (_28029_, _10004_, _03568_);
  and _78563_ (_28030_, _28029_, _10307_);
  and _78564_ (_28031_, _28030_, _28028_);
  nor _78565_ (_28032_, _27974_, _10307_);
  or _78566_ (_28033_, _28032_, _03575_);
  or _78567_ (_28034_, _28033_, _28031_);
  nand _78568_ (_28035_, _10004_, _03575_);
  and _78569_ (_28036_, _28035_, _10316_);
  and _78570_ (_28037_, _28036_, _28034_);
  nor _78571_ (_28039_, _27974_, _10316_);
  or _78572_ (_28040_, _28039_, _03512_);
  or _78573_ (_28041_, _28040_, _28037_);
  nand _78574_ (_28042_, _10004_, _03512_);
  and _78575_ (_28043_, _28042_, _03206_);
  and _78576_ (_28044_, _28043_, _28041_);
  nor _78577_ (_28045_, _06132_, _03206_);
  or _78578_ (_28046_, _28045_, _28044_);
  and _78579_ (_28047_, _28046_, _04887_);
  nand _78580_ (_28048_, _10003_, _03511_);
  nand _78581_ (_28050_, _28048_, _10325_);
  or _78582_ (_28051_, _28050_, _28047_);
  or _78583_ (_28052_, _27984_, _10360_);
  nand _78584_ (_28053_, _10360_, _10166_);
  and _78585_ (_28054_, _28053_, _28052_);
  or _78586_ (_28055_, _28054_, _10325_);
  and _78587_ (_28056_, _28055_, _28051_);
  or _78588_ (_28057_, _28056_, _27272_);
  and _78589_ (_28058_, _28057_, _27988_);
  or _78590_ (_28059_, _28058_, _03527_);
  not _78591_ (_28061_, _27984_);
  nor _78592_ (_28062_, _28061_, _10382_);
  and _78593_ (_28063_, _10382_, _10165_);
  or _78594_ (_28064_, _28063_, _03998_);
  or _78595_ (_28065_, _28064_, _28062_);
  and _78596_ (_28066_, _28065_, _10085_);
  and _78597_ (_28067_, _28066_, _28059_);
  or _78598_ (_28068_, _27984_, _10398_);
  nand _78599_ (_28069_, _10398_, _10166_);
  and _78600_ (_28070_, _28069_, _03638_);
  and _78601_ (_28072_, _28070_, _28068_);
  or _78602_ (_28073_, _28072_, _10083_);
  or _78603_ (_28074_, _28073_, _28067_);
  and _78604_ (_28075_, _28074_, _27981_);
  or _78605_ (_28076_, _28075_, _03505_);
  nand _78606_ (_28077_, _10004_, _03505_);
  and _78607_ (_28078_, _28077_, _03200_);
  and _78608_ (_28079_, _28078_, _28076_);
  nor _78609_ (_28080_, _06132_, _03200_);
  or _78610_ (_28081_, _28080_, _26282_);
  or _78611_ (_28083_, _28081_, _28079_);
  or _78612_ (_28084_, _26281_, _10003_);
  and _78613_ (_28085_, _28084_, _28083_);
  or _78614_ (_28086_, _28085_, _25991_);
  or _78615_ (_28087_, _27973_, _10415_);
  and _78616_ (_28088_, _28087_, _10419_);
  and _78617_ (_28089_, _28088_, _28086_);
  and _78618_ (_28090_, _10003_, _03607_);
  or _78619_ (_28091_, _28090_, _10420_);
  or _78620_ (_28092_, _28091_, _28089_);
  nand _78621_ (_28094_, _06132_, _10420_);
  and _78622_ (_28095_, _28094_, _11467_);
  and _78623_ (_28096_, _28095_, _28092_);
  nand _78624_ (_28097_, _10003_, _03606_);
  nand _78625_ (_28098_, _28097_, _10426_);
  or _78626_ (_28099_, _28098_, _28096_);
  or _78627_ (_28100_, _27973_, _10426_);
  and _78628_ (_28101_, _28100_, _10430_);
  and _78629_ (_28102_, _28101_, _28099_);
  nor _78630_ (_28103_, _10004_, _10430_);
  or _78631_ (_28105_, _28103_, _03311_);
  or _78632_ (_28106_, _28105_, _28102_);
  or _78633_ (_28107_, _27973_, _03254_);
  and _78634_ (_28108_, _28107_, _28106_);
  or _78635_ (_28109_, _28108_, _03499_);
  nand _78636_ (_28110_, _10004_, _03499_);
  and _78637_ (_28111_, _28110_, _04853_);
  and _78638_ (_28112_, _28111_, _28109_);
  nor _78639_ (_28113_, _06132_, _04853_);
  or _78640_ (_28114_, _28113_, _03632_);
  or _78641_ (_28116_, _28114_, _28112_);
  nand _78642_ (_28117_, _10166_, _03632_);
  and _78643_ (_28118_, _28117_, _28116_);
  or _78644_ (_28119_, _28118_, _26322_);
  or _78645_ (_28120_, _10003_, _03493_);
  and _78646_ (_28121_, _28120_, _28119_);
  or _78647_ (_28122_, _28121_, _03221_);
  nand _78648_ (_28123_, _10166_, _03221_);
  and _78649_ (_28124_, _28123_, _10081_);
  and _78650_ (_28125_, _28124_, _28122_);
  nor _78651_ (_28127_, _27974_, _10081_);
  or _78652_ (_28128_, _28127_, _03745_);
  or _78653_ (_28129_, _28128_, _28125_);
  nand _78654_ (_28130_, _10004_, _03745_);
  and _78655_ (_28131_, _28130_, _26022_);
  and _78656_ (_28132_, _28131_, _28129_);
  nor _78657_ (_28133_, _06132_, _26022_);
  or _78658_ (_28134_, _28133_, _28132_);
  and _78659_ (_28135_, _28134_, _10459_);
  or _78660_ (_28136_, _28135_, _27980_);
  and _78661_ (_28138_, _28136_, _05775_);
  nor _78662_ (_28139_, _10004_, _05775_);
  or _78663_ (_28140_, _28139_, _03437_);
  or _78664_ (_28141_, _28140_, _28138_);
  nand _78665_ (_28142_, _10166_, _03437_);
  and _78666_ (_28143_, _28142_, _08386_);
  and _78667_ (_28144_, _28143_, _28141_);
  and _78668_ (_28145_, _10003_, _08385_);
  or _78669_ (_28146_, _28145_, _10472_);
  or _78670_ (_28147_, _28146_, _28144_);
  nor _78671_ (_28149_, _10495_, _10481_);
  nor _78672_ (_28150_, _28149_, _10496_);
  or _78673_ (_28151_, _28150_, _25897_);
  and _78674_ (_28152_, _28151_, _04118_);
  and _78675_ (_28153_, _28152_, _28147_);
  and _78676_ (_28154_, _10003_, _03744_);
  or _78677_ (_28155_, _28154_, _03189_);
  or _78678_ (_28156_, _28155_, _28153_);
  nand _78679_ (_28157_, _06132_, _03189_);
  and _78680_ (_28158_, _28157_, _10515_);
  and _78681_ (_28160_, _28158_, _28156_);
  or _78682_ (_28161_, _27979_, _08698_);
  or _78683_ (_28162_, _10003_, _10077_);
  and _78684_ (_28163_, _28162_, _10076_);
  and _78685_ (_28164_, _28163_, _28161_);
  or _78686_ (_28165_, _28164_, _26754_);
  or _78687_ (_28166_, _28165_, _28160_);
  or _78688_ (_28167_, _27973_, _10520_);
  and _78689_ (_28168_, _28167_, _10523_);
  and _78690_ (_28169_, _28168_, _28166_);
  nor _78691_ (_28171_, _10523_, _10004_);
  or _78692_ (_28172_, _28171_, _03636_);
  or _78693_ (_28173_, _28172_, _28169_);
  and _78694_ (_28174_, _28173_, _27977_);
  or _78695_ (_28175_, _28174_, _03769_);
  nand _78696_ (_28176_, _10004_, _03769_);
  and _78697_ (_28177_, _28176_, _25894_);
  and _78698_ (_28178_, _28177_, _28175_);
  nor _78699_ (_28179_, _06132_, _25894_);
  or _78700_ (_28180_, _28179_, _28178_);
  and _78701_ (_28182_, _28180_, _10535_);
  or _78702_ (_28183_, _27979_, _10077_);
  or _78703_ (_28184_, _10003_, _08698_);
  and _78704_ (_28185_, _28184_, _10534_);
  and _78705_ (_28186_, _28185_, _28183_);
  or _78706_ (_28187_, _28186_, _10545_);
  or _78707_ (_28188_, _28187_, _28182_);
  nand _78708_ (_28189_, _27974_, _10545_);
  and _78709_ (_28190_, _28189_, _10548_);
  and _78710_ (_28191_, _28190_, _28188_);
  nor _78711_ (_28193_, _10004_, _10548_);
  or _78712_ (_28194_, _28193_, _03754_);
  or _78713_ (_28195_, _28194_, _28191_);
  nand _78714_ (_28196_, _10166_, _03754_);
  and _78715_ (_28197_, _28196_, _28195_);
  or _78716_ (_28198_, _28197_, _03752_);
  nand _78717_ (_28199_, _10004_, _03752_);
  and _78718_ (_28200_, _28199_, _25891_);
  and _78719_ (_28201_, _28200_, _28198_);
  nor _78720_ (_28202_, _06132_, _25891_);
  or _78721_ (_28204_, _28202_, _28201_);
  and _78722_ (_28205_, _28204_, _09959_);
  or _78723_ (_28206_, _27979_, \oc8051_golden_model_1.PSW [7]);
  or _78724_ (_28207_, _10003_, _07888_);
  and _78725_ (_28208_, _28207_, _09958_);
  and _78726_ (_28209_, _28208_, _28206_);
  or _78727_ (_28210_, _28209_, _10560_);
  or _78728_ (_28211_, _28210_, _28205_);
  or _78729_ (_28212_, _27973_, _09956_);
  and _78730_ (_28213_, _28212_, _08478_);
  and _78731_ (_28215_, _28213_, _28211_);
  nor _78732_ (_28216_, _10004_, _08478_);
  or _78733_ (_28217_, _28216_, _03758_);
  or _78734_ (_28218_, _28217_, _28215_);
  and _78735_ (_28219_, _28218_, _27976_);
  or _78736_ (_28220_, _28219_, _03760_);
  nand _78737_ (_28221_, _10004_, _03760_);
  and _78738_ (_28222_, _28221_, _26082_);
  and _78739_ (_28223_, _28222_, _28220_);
  nor _78740_ (_28224_, _06132_, _26082_);
  or _78741_ (_28226_, _28224_, _28223_);
  and _78742_ (_28227_, _28226_, _10577_);
  or _78743_ (_28228_, _27979_, _07888_);
  or _78744_ (_28229_, _10003_, \oc8051_golden_model_1.PSW [7]);
  and _78745_ (_28230_, _28229_, _10576_);
  and _78746_ (_28231_, _28230_, _28228_);
  or _78747_ (_28232_, _28231_, _10581_);
  or _78748_ (_28233_, _28232_, _28227_);
  or _78749_ (_28234_, _27973_, _09951_);
  and _78750_ (_28235_, _28234_, _08524_);
  and _78751_ (_28237_, _28235_, _28233_);
  nor _78752_ (_28238_, _10004_, _08524_);
  or _78753_ (_28239_, _28238_, _08555_);
  or _78754_ (_28240_, _28239_, _28237_);
  nand _78755_ (_28241_, _27974_, _08555_);
  and _78756_ (_28242_, _28241_, _11403_);
  and _78757_ (_28243_, _28242_, _28240_);
  and _78758_ (_28244_, _06713_, _03775_);
  or _78759_ (_28245_, _28244_, _03179_);
  or _78760_ (_28246_, _28245_, _28243_);
  nand _78761_ (_28247_, _06132_, _03179_);
  and _78762_ (_28248_, _28247_, _10599_);
  and _78763_ (_28249_, _28248_, _28246_);
  nand _78764_ (_28250_, _28061_, _10794_);
  or _78765_ (_28251_, _10794_, _10165_);
  and _78766_ (_28252_, _28251_, _03627_);
  and _78767_ (_28253_, _28252_, _28250_);
  or _78768_ (_28254_, _28253_, _10603_);
  or _78769_ (_28255_, _28254_, _28249_);
  or _78770_ (_28256_, _27973_, _09949_);
  and _78771_ (_28259_, _28256_, _09936_);
  and _78772_ (_28260_, _28259_, _28255_);
  nor _78773_ (_28261_, _10004_, _09936_);
  or _78774_ (_28262_, _28261_, _07729_);
  or _78775_ (_28263_, _28262_, _28260_);
  and _78776_ (_28264_, _28263_, _27975_);
  or _78777_ (_28265_, _28264_, _03522_);
  or _78778_ (_28266_, _06713_, _03523_);
  and _78779_ (_28267_, _28266_, _25887_);
  and _78780_ (_28268_, _28267_, _28265_);
  nor _78781_ (_28270_, _06132_, _25887_);
  or _78782_ (_28271_, _28270_, _03628_);
  or _78783_ (_28272_, _28271_, _28268_);
  or _78784_ (_28273_, _27984_, _10794_);
  nand _78785_ (_28274_, _10794_, _10166_);
  and _78786_ (_28275_, _28274_, _28273_);
  or _78787_ (_28276_, _28275_, _03791_);
  and _78788_ (_28277_, _28276_, _28272_);
  or _78789_ (_28278_, _28277_, _10822_);
  or _78790_ (_28279_, _27973_, _10821_);
  and _78791_ (_28281_, _28279_, _28278_);
  or _78792_ (_28282_, _28281_, _03790_);
  nand _78793_ (_28283_, _10004_, _03790_);
  and _78794_ (_28284_, _28283_, _10828_);
  and _78795_ (_28285_, _28284_, _28282_);
  nor _78796_ (_28286_, _27974_, _10828_);
  or _78797_ (_28287_, _28286_, _04947_);
  or _78798_ (_28288_, _28287_, _28285_);
  and _78799_ (_28289_, _28288_, _27969_);
  or _78800_ (_28290_, _28289_, _03151_);
  or _78801_ (_28292_, _28275_, _03152_);
  and _78802_ (_28293_, _28292_, _10844_);
  and _78803_ (_28294_, _28293_, _28290_);
  nor _78804_ (_28295_, _27974_, _10844_);
  nor _78805_ (_28296_, _28295_, _03520_);
  not _78806_ (_28297_, _28296_);
  nor _78807_ (_28298_, _28297_, _28294_);
  not _78808_ (_28299_, _10851_);
  and _78809_ (_28300_, _10004_, _03520_);
  nor _78810_ (_28301_, _28300_, _28299_);
  not _78811_ (_28303_, _28301_);
  nor _78812_ (_28304_, _28303_, _28298_);
  nor _78813_ (_28305_, _27974_, _10851_);
  nor _78814_ (_28306_, _28305_, _25883_);
  not _78815_ (_28307_, _28306_);
  nor _78816_ (_28308_, _28307_, _28304_);
  and _78817_ (_28309_, _25883_, _06132_);
  or _78818_ (_28310_, _28309_, _10862_);
  nor _78819_ (_28311_, _28310_, _28308_);
  and _78820_ (_28312_, _27973_, _10862_);
  nor _78821_ (_28314_, _28312_, _28311_);
  nand _78822_ (_28315_, _28314_, _42963_);
  or _78823_ (_28316_, _42963_, \oc8051_golden_model_1.PC [6]);
  and _78824_ (_28317_, _28316_, _41755_);
  and _78825_ (_43335_, _28317_, _28315_);
  and _78826_ (_28318_, _05841_, _03520_);
  and _78827_ (_28319_, _05841_, _03790_);
  nor _78828_ (_28320_, _09939_, \oc8051_golden_model_1.PC [7]);
  nor _78829_ (_28321_, _28320_, _09940_);
  nor _78830_ (_28322_, _28321_, _09949_);
  nor _78831_ (_28324_, _28321_, _09956_);
  not _78832_ (_28325_, _28321_);
  and _78833_ (_28326_, _28325_, _10545_);
  nor _78834_ (_28327_, _28321_, _10520_);
  nor _78835_ (_28328_, _28321_, _10426_);
  and _78836_ (_28329_, _05841_, _03606_);
  nor _78837_ (_28330_, _28321_, _10415_);
  nor _78838_ (_28331_, _06086_, _03200_);
  nand _78839_ (_28332_, _10261_, _06680_);
  or _78840_ (_28333_, _10161_, _10162_);
  and _78841_ (_28335_, _28333_, _10212_);
  nor _78842_ (_28336_, _28333_, _10212_);
  nor _78843_ (_28337_, _28336_, _28335_);
  or _78844_ (_28338_, _28337_, _10261_);
  and _78845_ (_28339_, _28338_, _28332_);
  or _78846_ (_28340_, _28339_, _04444_);
  and _78847_ (_28341_, _10269_, _05841_);
  or _78848_ (_28342_, _09999_, _10000_);
  and _78849_ (_28343_, _28342_, _10043_);
  nor _78850_ (_28344_, _28342_, _10043_);
  nor _78851_ (_28346_, _28344_, _28343_);
  and _78852_ (_28347_, _28346_, _10271_);
  or _78853_ (_28348_, _28347_, _28341_);
  or _78854_ (_28349_, _28348_, _05831_);
  nand _78855_ (_28350_, _06086_, _03923_);
  or _78856_ (_28351_, _28321_, _10290_);
  or _78857_ (_28352_, _28321_, _25905_);
  nand _78858_ (_28353_, _05994_, _03922_);
  nor _78859_ (_28354_, _04426_, \oc8051_golden_model_1.PC [7]);
  nand _78860_ (_28355_, _28354_, _10278_);
  and _78861_ (_28357_, _28355_, _28353_);
  or _78862_ (_28358_, _28357_, _26577_);
  nand _78863_ (_28359_, _28358_, _28352_);
  nand _78864_ (_28360_, _28359_, _25909_);
  and _78865_ (_28361_, _28360_, _28351_);
  and _78866_ (_28362_, _28361_, _28350_);
  or _78867_ (_28363_, _28362_, _05833_);
  and _78868_ (_28364_, _28363_, _05847_);
  and _78869_ (_28365_, _28364_, _28349_);
  and _78870_ (_28366_, _28321_, _04438_);
  or _78871_ (_28368_, _28366_, _03570_);
  or _78872_ (_28369_, _28368_, _28365_);
  and _78873_ (_28370_, _28369_, _28340_);
  or _78874_ (_28371_, _28370_, _10256_);
  or _78875_ (_28372_, _28321_, _10255_);
  and _78876_ (_28373_, _28372_, _03517_);
  and _78877_ (_28374_, _28373_, _28371_);
  and _78878_ (_28375_, _05841_, _03516_);
  or _78879_ (_28376_, _28375_, _04746_);
  or _78880_ (_28377_, _28376_, _28374_);
  nand _78881_ (_28379_, _06086_, _04746_);
  and _78882_ (_28380_, _28379_, _03983_);
  and _78883_ (_28381_, _28380_, _28377_);
  nand _78884_ (_28382_, _05841_, _03568_);
  nand _78885_ (_28383_, _28382_, _10307_);
  or _78886_ (_28384_, _28383_, _28381_);
  or _78887_ (_28385_, _28321_, _10307_);
  and _78888_ (_28386_, _28385_, _03583_);
  and _78889_ (_28387_, _28386_, _28384_);
  nand _78890_ (_28388_, _05841_, _03575_);
  nand _78891_ (_28390_, _28388_, _10316_);
  or _78892_ (_28391_, _28390_, _28387_);
  or _78893_ (_28392_, _28321_, _10316_);
  and _78894_ (_28393_, _28392_, _03513_);
  and _78895_ (_28394_, _28393_, _28391_);
  and _78896_ (_28395_, _05841_, _03512_);
  or _78897_ (_28396_, _28395_, _10249_);
  or _78898_ (_28397_, _28396_, _28394_);
  nand _78899_ (_28398_, _06086_, _10249_);
  and _78900_ (_28399_, _28398_, _04887_);
  and _78901_ (_28401_, _28399_, _28397_);
  nand _78902_ (_28402_, _05841_, _03511_);
  nand _78903_ (_28403_, _28402_, _10325_);
  or _78904_ (_28404_, _28403_, _28401_);
  not _78905_ (_28405_, _28337_);
  nor _78906_ (_28406_, _28405_, _10360_);
  and _78907_ (_28407_, _10360_, _06679_);
  or _78908_ (_28408_, _28407_, _10325_);
  or _78909_ (_28409_, _28408_, _28406_);
  and _78910_ (_28410_, _28409_, _28404_);
  or _78911_ (_28412_, _28410_, _03657_);
  nand _78912_ (_28413_, _10116_, _06680_);
  or _78913_ (_28414_, _28337_, _10116_);
  and _78914_ (_28415_, _28414_, _28413_);
  or _78915_ (_28416_, _28415_, _10328_);
  and _78916_ (_28417_, _28416_, _11596_);
  and _78917_ (_28418_, _28417_, _28412_);
  and _78918_ (_28419_, _10382_, _06679_);
  nor _78919_ (_28420_, _28405_, _10382_);
  nor _78920_ (_28421_, _28420_, _28419_);
  nor _78921_ (_28423_, _28421_, _03998_);
  nor _78922_ (_28424_, _28337_, _10398_);
  and _78923_ (_28425_, _10398_, _06680_);
  nor _78924_ (_28426_, _28425_, _10085_);
  not _78925_ (_28427_, _28426_);
  nor _78926_ (_28428_, _28427_, _28424_);
  nor _78927_ (_28429_, _28428_, _28423_);
  and _78928_ (_28430_, _28321_, _10083_);
  nor _78929_ (_28431_, _28430_, _03505_);
  and _78930_ (_28432_, _28431_, _28429_);
  not _78931_ (_28433_, _28432_);
  nor _78932_ (_28434_, _28433_, _28418_);
  and _78933_ (_28435_, _05994_, _03505_);
  nor _78934_ (_28436_, _28435_, _04743_);
  not _78935_ (_28437_, _28436_);
  nor _78936_ (_28438_, _28437_, _28434_);
  nor _78937_ (_28439_, _28438_, _28331_);
  or _78938_ (_28440_, _28439_, _26282_);
  or _78939_ (_28441_, _26281_, _05994_);
  and _78940_ (_28442_, _28441_, _10415_);
  and _78941_ (_28445_, _28442_, _28440_);
  or _78942_ (_28446_, _28445_, _03607_);
  nor _78943_ (_28447_, _28446_, _28330_);
  and _78944_ (_28448_, _05841_, _03607_);
  or _78945_ (_28449_, _28448_, _28447_);
  and _78946_ (_28450_, _28449_, _03213_);
  nor _78947_ (_28451_, _06086_, _03213_);
  or _78948_ (_28452_, _28451_, _28450_);
  and _78949_ (_28453_, _28452_, _11467_);
  or _78950_ (_28454_, _28453_, _26302_);
  nor _78951_ (_28456_, _28454_, _28329_);
  or _78952_ (_28457_, _28456_, _28328_);
  nand _78953_ (_28458_, _28457_, _10430_);
  nor _78954_ (_28459_, _10430_, _05841_);
  nor _78955_ (_28460_, _28459_, _03311_);
  and _78956_ (_28461_, _28460_, _28458_);
  nor _78957_ (_28462_, _28325_, _03254_);
  or _78958_ (_28463_, _28462_, _03499_);
  nor _78959_ (_28464_, _28463_, _28461_);
  and _78960_ (_28465_, _05994_, _03499_);
  or _78961_ (_28467_, _28465_, _28464_);
  nand _78962_ (_28468_, _28467_, _04853_);
  and _78963_ (_28469_, _06086_, _03223_);
  nor _78964_ (_28470_, _28469_, _03632_);
  nand _78965_ (_28471_, _28470_, _28468_);
  and _78966_ (_28472_, _06679_, _03632_);
  nor _78967_ (_28473_, _28472_, _26322_);
  nand _78968_ (_28474_, _28473_, _28471_);
  nor _78969_ (_28475_, _05841_, _03493_);
  nor _78970_ (_28476_, _28475_, _03221_);
  nand _78971_ (_28478_, _28476_, _28474_);
  and _78972_ (_28479_, _06679_, _03221_);
  nor _78973_ (_28480_, _28479_, _26330_);
  nand _78974_ (_28481_, _28480_, _28478_);
  nor _78975_ (_28482_, _28321_, _10081_);
  nor _78976_ (_28483_, _28482_, _03745_);
  nand _78977_ (_28484_, _28483_, _28481_);
  and _78978_ (_28485_, _05841_, _03745_);
  nor _78979_ (_28486_, _28485_, _03187_);
  nand _78980_ (_28487_, _28486_, _28484_);
  and _78981_ (_28489_, _06086_, _03187_);
  nor _78982_ (_28490_, _28489_, _10458_);
  nand _78983_ (_28491_, _28490_, _28487_);
  and _78984_ (_28492_, _28346_, _10458_);
  nor _78985_ (_28493_, _28492_, _06055_);
  nand _78986_ (_28494_, _28493_, _28491_);
  nor _78987_ (_28495_, _05841_, _05775_);
  nor _78988_ (_28496_, _28495_, _03437_);
  nand _78989_ (_28497_, _28496_, _28494_);
  and _78990_ (_28498_, _06679_, _03437_);
  nor _78991_ (_28500_, _28498_, _08385_);
  nand _78992_ (_28501_, _28500_, _28497_);
  and _78993_ (_28502_, _08385_, _05994_);
  nor _78994_ (_28503_, _28502_, _10472_);
  and _78995_ (_28504_, _28503_, _28501_);
  or _78996_ (_28505_, _10478_, _10477_);
  nor _78997_ (_28506_, _28505_, _10497_);
  and _78998_ (_28507_, _28505_, _10497_);
  nor _78999_ (_28508_, _28507_, _28506_);
  and _79000_ (_28509_, _28508_, _10472_);
  or _79001_ (_28511_, _28509_, _03744_);
  nor _79002_ (_28512_, _28511_, _28504_);
  and _79003_ (_28513_, _05994_, _03744_);
  or _79004_ (_28514_, _28513_, _28512_);
  nand _79005_ (_28515_, _28514_, _11376_);
  and _79006_ (_28516_, _06086_, _03189_);
  nor _79007_ (_28517_, _28516_, _10076_);
  nand _79008_ (_28518_, _28517_, _28515_);
  and _79009_ (_28519_, _08698_, _05841_);
  and _79010_ (_28520_, _28346_, _10077_);
  or _79011_ (_28522_, _28520_, _28519_);
  and _79012_ (_28523_, _28522_, _10076_);
  nor _79013_ (_28524_, _28523_, _26754_);
  and _79014_ (_28525_, _28524_, _28518_);
  or _79015_ (_28526_, _28525_, _28327_);
  nand _79016_ (_28527_, _28526_, _10523_);
  nor _79017_ (_28528_, _10523_, _05841_);
  nor _79018_ (_28529_, _28528_, _03636_);
  and _79019_ (_28530_, _28529_, _28527_);
  and _79020_ (_28531_, _06679_, _03636_);
  or _79021_ (_28533_, _28531_, _03769_);
  nor _79022_ (_28534_, _28533_, _28530_);
  and _79023_ (_28535_, _05994_, _03769_);
  or _79024_ (_28536_, _28535_, _28534_);
  nand _79025_ (_28537_, _28536_, _25894_);
  and _79026_ (_28538_, _06086_, _03194_);
  nor _79027_ (_28539_, _28538_, _10534_);
  nand _79028_ (_28540_, _28539_, _28537_);
  nor _79029_ (_28541_, _28346_, _10077_);
  nor _79030_ (_28542_, _08698_, _05841_);
  nor _79031_ (_28544_, _28542_, _10535_);
  not _79032_ (_28545_, _28544_);
  nor _79033_ (_28546_, _28545_, _28541_);
  nor _79034_ (_28547_, _28546_, _10545_);
  and _79035_ (_28548_, _28547_, _28540_);
  or _79036_ (_28549_, _28548_, _28326_);
  nand _79037_ (_28550_, _28549_, _10548_);
  nor _79038_ (_28551_, _10548_, _05841_);
  nor _79039_ (_28552_, _28551_, _04504_);
  nand _79040_ (_28553_, _28552_, _28550_);
  and _79041_ (_28555_, _06679_, _03754_);
  nor _79042_ (_28556_, _28555_, _03752_);
  and _79043_ (_28557_, _28556_, _28553_);
  and _79044_ (_28558_, _05994_, _03752_);
  or _79045_ (_28559_, _28558_, _28557_);
  nand _79046_ (_28560_, _28559_, _25891_);
  and _79047_ (_28561_, _06086_, _03192_);
  nor _79048_ (_28562_, _28561_, _09958_);
  nand _79049_ (_28563_, _28562_, _28560_);
  and _79050_ (_28564_, _05841_, \oc8051_golden_model_1.PSW [7]);
  and _79051_ (_28566_, _28346_, _07888_);
  or _79052_ (_28567_, _28566_, _28564_);
  and _79053_ (_28568_, _28567_, _09958_);
  nor _79054_ (_28569_, _28568_, _10560_);
  and _79055_ (_28570_, _28569_, _28563_);
  or _79056_ (_28571_, _28570_, _28324_);
  nand _79057_ (_28572_, _28571_, _08478_);
  nor _79058_ (_28573_, _08478_, _05841_);
  nor _79059_ (_28574_, _28573_, _03758_);
  nand _79060_ (_28575_, _28574_, _28572_);
  and _79061_ (_28577_, _06679_, _03758_);
  nor _79062_ (_28578_, _28577_, _03760_);
  and _79063_ (_28579_, _28578_, _28575_);
  and _79064_ (_28580_, _05994_, _03760_);
  nor _79065_ (_28581_, _28580_, _28579_);
  nand _79066_ (_28582_, _28581_, _26077_);
  nor _79067_ (_28583_, _06086_, _26082_);
  nor _79068_ (_28584_, _28346_, _07888_);
  nor _79069_ (_28585_, _05841_, \oc8051_golden_model_1.PSW [7]);
  nor _79070_ (_28586_, _28585_, _10577_);
  not _79071_ (_28588_, _28586_);
  nor _79072_ (_28589_, _28588_, _28584_);
  nor _79073_ (_28590_, _28589_, _28583_);
  and _79074_ (_28591_, _28590_, _28582_);
  or _79075_ (_28592_, _28591_, _10581_);
  or _79076_ (_28593_, _28325_, _09951_);
  and _79077_ (_28594_, _28593_, _08524_);
  nand _79078_ (_28595_, _28594_, _28592_);
  nor _79079_ (_28596_, _08524_, _05841_);
  nor _79080_ (_28597_, _28596_, _08555_);
  and _79081_ (_28599_, _28597_, _28595_);
  and _79082_ (_28600_, _28321_, _08555_);
  or _79083_ (_28601_, _28600_, _03775_);
  nor _79084_ (_28602_, _28601_, _28599_);
  and _79085_ (_28603_, _06004_, _03775_);
  or _79086_ (_28604_, _28603_, _28602_);
  nand _79087_ (_28605_, _28604_, _06328_);
  and _79088_ (_28606_, _06086_, _03179_);
  nor _79089_ (_28607_, _28606_, _03627_);
  nand _79090_ (_28608_, _28607_, _28605_);
  and _79091_ (_28610_, _28405_, _10794_);
  nor _79092_ (_28611_, _10794_, _06679_);
  or _79093_ (_28612_, _28611_, _10599_);
  or _79094_ (_28613_, _28612_, _28610_);
  and _79095_ (_28614_, _28613_, _09949_);
  and _79096_ (_28615_, _28614_, _28608_);
  or _79097_ (_28616_, _28615_, _28322_);
  nand _79098_ (_28617_, _28616_, _09936_);
  nor _79099_ (_28618_, _09936_, _05841_);
  nor _79100_ (_28619_, _28618_, _07729_);
  and _79101_ (_28621_, _28619_, _28617_);
  and _79102_ (_28622_, _28321_, _07729_);
  or _79103_ (_28623_, _28622_, _03522_);
  nor _79104_ (_28624_, _28623_, _28621_);
  and _79105_ (_28625_, _06004_, _03522_);
  or _79106_ (_28626_, _28625_, _28624_);
  nand _79107_ (_28627_, _28626_, _25887_);
  and _79108_ (_28628_, _06086_, _03172_);
  nor _79109_ (_28629_, _28628_, _03628_);
  nand _79110_ (_28630_, _28629_, _28627_);
  and _79111_ (_28632_, _10794_, _06680_);
  nor _79112_ (_28633_, _28337_, _10794_);
  nor _79113_ (_28634_, _28633_, _28632_);
  and _79114_ (_28635_, _28634_, _03628_);
  nor _79115_ (_28636_, _28635_, _10822_);
  nand _79116_ (_28637_, _28636_, _28630_);
  nor _79117_ (_28638_, _28321_, _10821_);
  nor _79118_ (_28639_, _28638_, _03790_);
  and _79119_ (_28640_, _28639_, _28637_);
  or _79120_ (_28641_, _28640_, _28319_);
  nand _79121_ (_28642_, _28641_, _10828_);
  nor _79122_ (_28643_, _28325_, _10828_);
  nor _79123_ (_28644_, _28643_, _04947_);
  nand _79124_ (_28645_, _28644_, _28642_);
  and _79125_ (_28646_, _06086_, _04947_);
  nor _79126_ (_28647_, _28646_, _03151_);
  nand _79127_ (_28648_, _28647_, _28645_);
  and _79128_ (_28649_, _28634_, _03151_);
  nor _79129_ (_28650_, _28649_, _10845_);
  nand _79130_ (_28651_, _28650_, _28648_);
  nor _79131_ (_28653_, _28321_, _10844_);
  nor _79132_ (_28654_, _28653_, _03520_);
  and _79133_ (_28655_, _28654_, _28651_);
  or _79134_ (_28656_, _28655_, _28318_);
  nand _79135_ (_28657_, _28656_, _10851_);
  nor _79136_ (_28658_, _28325_, _10851_);
  nor _79137_ (_28659_, _28658_, _25883_);
  nand _79138_ (_28660_, _28659_, _28657_);
  and _79139_ (_28661_, _25883_, _06086_);
  nor _79140_ (_28662_, _28661_, _10862_);
  and _79141_ (_28664_, _28662_, _28660_);
  and _79142_ (_28665_, _28321_, _10862_);
  or _79143_ (_28666_, _28665_, _28664_);
  or _79144_ (_28667_, _28666_, _42967_);
  or _79145_ (_28668_, _42963_, \oc8051_golden_model_1.PC [7]);
  and _79146_ (_28669_, _28668_, _41755_);
  and _79147_ (_43336_, _28669_, _28667_);
  nor _79148_ (_28670_, _10855_, _03471_);
  nor _79149_ (_28671_, _10832_, _03471_);
  and _79150_ (_28672_, _09940_, \oc8051_golden_model_1.PC [8]);
  nor _79151_ (_28674_, _09940_, \oc8051_golden_model_1.PC [8]);
  nor _79152_ (_28675_, _28674_, _28672_);
  and _79153_ (_28676_, _28675_, _07729_);
  nor _79154_ (_28677_, _28675_, _09949_);
  and _79155_ (_28678_, _28675_, _08555_);
  nor _79156_ (_28679_, _28675_, _09951_);
  nor _79157_ (_28680_, _28675_, _09956_);
  not _79158_ (_28681_, _28675_);
  and _79159_ (_28682_, _28681_, _10545_);
  and _79160_ (_28683_, _10216_, _03636_);
  nor _79161_ (_28685_, _28675_, _10520_);
  nor _79162_ (_28686_, _10458_, _03187_);
  not _79163_ (_28687_, _28686_);
  and _79164_ (_28688_, _10047_, _03745_);
  not _79165_ (_28689_, _28688_);
  nor _79166_ (_28690_, _28675_, _10081_);
  nor _79167_ (_28691_, _10047_, _10430_);
  nor _79168_ (_28692_, _28675_, _10415_);
  nor _79169_ (_28693_, _26281_, _10047_);
  and _79170_ (_28694_, _28675_, _10083_);
  not _79171_ (_28696_, _28694_);
  and _79172_ (_28697_, _10382_, _10216_);
  nor _79173_ (_28698_, _10220_, _10214_);
  nor _79174_ (_28699_, _28698_, _10221_);
  not _79175_ (_28700_, _28699_);
  nor _79176_ (_28701_, _28700_, _10382_);
  nor _79177_ (_28702_, _28701_, _28697_);
  nor _79178_ (_28703_, _28702_, _03998_);
  and _79179_ (_28704_, _10398_, _10216_);
  and _79180_ (_28705_, _28699_, _10399_);
  or _79181_ (_28707_, _28705_, _28704_);
  and _79182_ (_28708_, _28707_, _03638_);
  nor _79183_ (_28709_, _28708_, _28703_);
  nand _79184_ (_28710_, _28709_, _28696_);
  and _79185_ (_28711_, _10047_, _03512_);
  or _79186_ (_28712_, _03568_, _04746_);
  nand _79187_ (_28713_, _10047_, _03516_);
  and _79188_ (_28714_, _10261_, _10217_);
  nor _79189_ (_28715_, _28699_, _10261_);
  or _79190_ (_28716_, _28715_, _28714_);
  and _79191_ (_28718_, _28716_, _03570_);
  or _79192_ (_28719_, _10271_, _12052_);
  nor _79193_ (_28720_, _10050_, _10045_);
  nor _79194_ (_28721_, _28720_, _10051_);
  nand _79195_ (_28722_, _28721_, _10271_);
  and _79196_ (_28723_, _28722_, _28719_);
  and _79197_ (_28724_, _28723_, _05833_);
  nand _79198_ (_28725_, _10290_, _10278_);
  and _79199_ (_28726_, _28725_, _28681_);
  and _79200_ (_28727_, _12052_, _03922_);
  or _79201_ (_28729_, _28727_, _26577_);
  nor _79202_ (_28730_, _04426_, \oc8051_golden_model_1.PC [8]);
  and _79203_ (_28731_, _28730_, _10278_);
  or _79204_ (_28732_, _28731_, _28729_);
  and _79205_ (_28733_, _28732_, _25909_);
  or _79206_ (_28734_, _28733_, _28726_);
  nand _79207_ (_28735_, _28675_, _26577_);
  and _79208_ (_28736_, _28735_, _05831_);
  and _79209_ (_28737_, _28736_, _28734_);
  or _79210_ (_28738_, _28737_, _04438_);
  or _79211_ (_28740_, _28738_, _28724_);
  nand _79212_ (_28741_, _28675_, _04438_);
  and _79213_ (_28742_, _28741_, _04444_);
  and _79214_ (_28743_, _28742_, _28740_);
  or _79215_ (_28744_, _28743_, _28718_);
  and _79216_ (_28745_, _28744_, _10255_);
  nor _79217_ (_28746_, _28675_, _10255_);
  or _79218_ (_28747_, _28746_, _03516_);
  or _79219_ (_28748_, _28747_, _28745_);
  and _79220_ (_28749_, _28748_, _28713_);
  nor _79221_ (_28751_, _28749_, _28712_);
  nand _79222_ (_28752_, _10047_, _03568_);
  nand _79223_ (_28753_, _28752_, _10307_);
  or _79224_ (_28754_, _28753_, _28751_);
  or _79225_ (_28755_, _28675_, _10307_);
  and _79226_ (_28756_, _28755_, _03583_);
  and _79227_ (_28757_, _28756_, _28754_);
  nand _79228_ (_28758_, _10047_, _03575_);
  nand _79229_ (_28759_, _28758_, _10316_);
  or _79230_ (_28760_, _28759_, _28757_);
  or _79231_ (_28762_, _28675_, _10316_);
  and _79232_ (_28763_, _28762_, _03513_);
  and _79233_ (_28764_, _28763_, _28760_);
  or _79234_ (_28765_, _28764_, _28711_);
  and _79235_ (_28766_, _28765_, _10250_);
  nand _79236_ (_28767_, _10047_, _03511_);
  nand _79237_ (_28768_, _28767_, _10325_);
  or _79238_ (_28769_, _28768_, _28766_);
  nor _79239_ (_28770_, _28700_, _10360_);
  and _79240_ (_28771_, _10360_, _10216_);
  or _79241_ (_28773_, _28771_, _10325_);
  or _79242_ (_28774_, _28773_, _28770_);
  and _79243_ (_28775_, _28774_, _28769_);
  or _79244_ (_28776_, _28775_, _03657_);
  nand _79245_ (_28777_, _10217_, _10116_);
  or _79246_ (_28778_, _28699_, _10116_);
  and _79247_ (_28779_, _28778_, _28777_);
  or _79248_ (_28780_, _28779_, _10328_);
  and _79249_ (_28781_, _28780_, _11596_);
  and _79250_ (_28782_, _28781_, _28776_);
  nor _79251_ (_28784_, _28782_, _28710_);
  nor _79252_ (_28785_, _28784_, _03505_);
  and _79253_ (_28786_, _26281_, _03200_);
  and _79254_ (_28787_, _10047_, _03505_);
  not _79255_ (_28788_, _28787_);
  and _79256_ (_28789_, _28788_, _28786_);
  not _79257_ (_28790_, _28789_);
  nor _79258_ (_28791_, _28790_, _28785_);
  nor _79259_ (_28792_, _28791_, _28693_);
  nor _79260_ (_28793_, _28792_, _25991_);
  or _79261_ (_28795_, _28793_, _03607_);
  nor _79262_ (_28796_, _28795_, _28692_);
  and _79263_ (_28797_, _10047_, _03607_);
  or _79264_ (_28798_, _28797_, _10420_);
  nor _79265_ (_28799_, _28798_, _28796_);
  nor _79266_ (_28800_, _28799_, _03606_);
  and _79267_ (_28801_, _10047_, _03606_);
  nor _79268_ (_28802_, _28801_, _26302_);
  not _79269_ (_28803_, _28802_);
  nor _79270_ (_28804_, _28803_, _28800_);
  nor _79271_ (_28806_, _28675_, _10426_);
  nor _79272_ (_28807_, _28806_, _28804_);
  nor _79273_ (_28808_, _28807_, _10431_);
  or _79274_ (_28809_, _28808_, _03311_);
  nor _79275_ (_28810_, _28809_, _28691_);
  nor _79276_ (_28811_, _28681_, _03254_);
  or _79277_ (_28812_, _28811_, _28810_);
  and _79278_ (_28813_, _28812_, _03500_);
  and _79279_ (_28814_, _10047_, _03499_);
  or _79280_ (_28815_, _28814_, _28813_);
  and _79281_ (_28817_, _28815_, _04853_);
  and _79282_ (_28818_, _28817_, _09755_);
  and _79283_ (_28819_, _10216_, _03632_);
  nor _79284_ (_28820_, _28819_, _26322_);
  not _79285_ (_28821_, _28820_);
  nor _79286_ (_28822_, _28821_, _28818_);
  nor _79287_ (_28823_, _10047_, _03493_);
  nor _79288_ (_28824_, _28823_, _03221_);
  not _79289_ (_28825_, _28824_);
  nor _79290_ (_28826_, _28825_, _28822_);
  and _79291_ (_28828_, _10216_, _03221_);
  nor _79292_ (_28829_, _28828_, _26330_);
  not _79293_ (_28830_, _28829_);
  nor _79294_ (_28831_, _28830_, _28826_);
  or _79295_ (_28832_, _28831_, _03745_);
  or _79296_ (_28833_, _28832_, _28690_);
  and _79297_ (_28834_, _28833_, _28689_);
  or _79298_ (_28835_, _28834_, _28687_);
  and _79299_ (_28836_, _28721_, _10458_);
  nor _79300_ (_28837_, _28836_, _06055_);
  and _79301_ (_28839_, _28837_, _28835_);
  nor _79302_ (_28840_, _10047_, _05775_);
  nor _79303_ (_28841_, _28840_, _03437_);
  not _79304_ (_28842_, _28841_);
  or _79305_ (_28843_, _28842_, _28839_);
  and _79306_ (_28844_, _10216_, _03437_);
  nor _79307_ (_28845_, _28844_, _08385_);
  nand _79308_ (_28846_, _28845_, _28843_);
  and _79309_ (_28847_, _12052_, _08385_);
  nor _79310_ (_28848_, _28847_, _10472_);
  and _79311_ (_28850_, _28848_, _28846_);
  and _79312_ (_28851_, _10499_, _10476_);
  not _79313_ (_28852_, _28851_);
  nor _79314_ (_28853_, _10500_, _25897_);
  and _79315_ (_28854_, _28853_, _28852_);
  or _79316_ (_28855_, _28854_, _28850_);
  nand _79317_ (_28856_, _28855_, _04118_);
  and _79318_ (_28857_, _10047_, _03744_);
  nor _79319_ (_28858_, _28857_, _03189_);
  nand _79320_ (_28859_, _28858_, _28856_);
  nand _79321_ (_28861_, _28859_, _10515_);
  and _79322_ (_28862_, _10047_, _08698_);
  and _79323_ (_28863_, _28721_, _10077_);
  or _79324_ (_28864_, _28863_, _28862_);
  and _79325_ (_28865_, _28864_, _10076_);
  nor _79326_ (_28866_, _28865_, _26754_);
  and _79327_ (_28867_, _28866_, _28861_);
  or _79328_ (_28868_, _28867_, _28685_);
  nand _79329_ (_28869_, _28868_, _10523_);
  nor _79330_ (_28870_, _10523_, _10047_);
  nor _79331_ (_28872_, _28870_, _03636_);
  and _79332_ (_28873_, _28872_, _28869_);
  or _79333_ (_28874_, _28873_, _28683_);
  nand _79334_ (_28875_, _28874_, _04501_);
  and _79335_ (_28876_, _10047_, _03769_);
  nor _79336_ (_28877_, _28876_, _03194_);
  nand _79337_ (_28878_, _28877_, _28875_);
  nand _79338_ (_28879_, _28878_, _10535_);
  nor _79339_ (_28880_, _28721_, _10077_);
  nor _79340_ (_28881_, _10047_, _08698_);
  nor _79341_ (_28883_, _28881_, _10535_);
  not _79342_ (_28884_, _28883_);
  nor _79343_ (_28885_, _28884_, _28880_);
  nor _79344_ (_28886_, _28885_, _10545_);
  and _79345_ (_28887_, _28886_, _28879_);
  or _79346_ (_28888_, _28887_, _28682_);
  nand _79347_ (_28889_, _28888_, _10548_);
  nor _79348_ (_28890_, _10047_, _10548_);
  nor _79349_ (_28891_, _28890_, _03754_);
  nand _79350_ (_28892_, _28891_, _28889_);
  and _79351_ (_28894_, _10216_, _03754_);
  nor _79352_ (_28895_, _28894_, _03752_);
  nand _79353_ (_28896_, _28895_, _28892_);
  nor _79354_ (_28897_, _09958_, _03192_);
  not _79355_ (_28898_, _28897_);
  and _79356_ (_28899_, _12052_, _03752_);
  nor _79357_ (_28900_, _28899_, _28898_);
  nand _79358_ (_28901_, _28900_, _28896_);
  and _79359_ (_28902_, _10047_, \oc8051_golden_model_1.PSW [7]);
  and _79360_ (_28903_, _28721_, _07888_);
  or _79361_ (_28905_, _28903_, _28902_);
  and _79362_ (_28906_, _28905_, _09958_);
  nor _79363_ (_28907_, _28906_, _10560_);
  and _79364_ (_28908_, _28907_, _28901_);
  or _79365_ (_28909_, _28908_, _28680_);
  nand _79366_ (_28910_, _28909_, _08478_);
  nor _79367_ (_28911_, _10047_, _08478_);
  nor _79368_ (_28912_, _28911_, _03758_);
  nand _79369_ (_28913_, _28912_, _28910_);
  and _79370_ (_28914_, _10216_, _03758_);
  nor _79371_ (_28916_, _28914_, _03760_);
  nand _79372_ (_28917_, _28916_, _28913_);
  and _79373_ (_28918_, _12052_, _03760_);
  nor _79374_ (_28919_, _28918_, _26078_);
  nand _79375_ (_28920_, _28919_, _28917_);
  nor _79376_ (_28921_, _28721_, _07888_);
  nor _79377_ (_28922_, _10047_, \oc8051_golden_model_1.PSW [7]);
  nor _79378_ (_28923_, _28922_, _10577_);
  not _79379_ (_28924_, _28923_);
  nor _79380_ (_28925_, _28924_, _28921_);
  nor _79381_ (_28927_, _28925_, _10581_);
  and _79382_ (_28928_, _28927_, _28920_);
  or _79383_ (_28929_, _28928_, _28679_);
  nand _79384_ (_28930_, _28929_, _08524_);
  nor _79385_ (_28931_, _10047_, _08524_);
  nor _79386_ (_28932_, _28931_, _08555_);
  and _79387_ (_28933_, _28932_, _28930_);
  or _79388_ (_28934_, _28933_, _28678_);
  nand _79389_ (_28935_, _28934_, _11403_);
  and _79390_ (_28936_, _04419_, _03775_);
  nor _79391_ (_28938_, _28936_, _03179_);
  nand _79392_ (_28939_, _28938_, _28935_);
  nand _79393_ (_28940_, _28939_, _10599_);
  and _79394_ (_28941_, _28700_, _10794_);
  nor _79395_ (_28942_, _10794_, _10216_);
  or _79396_ (_28943_, _28942_, _10599_);
  or _79397_ (_28944_, _28943_, _28941_);
  and _79398_ (_28945_, _28944_, _09949_);
  and _79399_ (_28946_, _28945_, _28940_);
  or _79400_ (_28947_, _28946_, _28677_);
  nand _79401_ (_28949_, _28947_, _09936_);
  nor _79402_ (_28950_, _10047_, _09936_);
  nor _79403_ (_28951_, _28950_, _07729_);
  and _79404_ (_28952_, _28951_, _28949_);
  or _79405_ (_28953_, _28952_, _28676_);
  nand _79406_ (_28954_, _28953_, _03523_);
  and _79407_ (_28955_, _04419_, _03522_);
  nor _79408_ (_28956_, _28955_, _03172_);
  nand _79409_ (_28957_, _28956_, _28954_);
  nand _79410_ (_28958_, _28957_, _03791_);
  and _79411_ (_28960_, _10794_, _10217_);
  nor _79412_ (_28961_, _28699_, _10794_);
  nor _79413_ (_28962_, _28961_, _28960_);
  and _79414_ (_28963_, _28962_, _03628_);
  nor _79415_ (_28964_, _28963_, _10822_);
  nand _79416_ (_28965_, _28964_, _28958_);
  nor _79417_ (_28966_, _28675_, _10821_);
  nor _79418_ (_28967_, _28966_, _03790_);
  nand _79419_ (_28968_, _28967_, _28965_);
  and _79420_ (_28969_, _10047_, _03790_);
  nor _79421_ (_28970_, _28969_, _27228_);
  nand _79422_ (_28971_, _28970_, _28968_);
  nor _79423_ (_28972_, _28675_, _10828_);
  nor _79424_ (_28973_, _28972_, _03641_);
  and _79425_ (_28974_, _28973_, _28971_);
  or _79426_ (_28975_, _28974_, _28671_);
  nor _79427_ (_28976_, _03160_, _03151_);
  nand _79428_ (_28977_, _28976_, _28975_);
  and _79429_ (_28978_, _28962_, _03151_);
  nor _79430_ (_28979_, _28978_, _10845_);
  nand _79431_ (_28982_, _28979_, _28977_);
  nor _79432_ (_28983_, _28675_, _10844_);
  nor _79433_ (_28984_, _28983_, _03520_);
  nand _79434_ (_28985_, _28984_, _28982_);
  and _79435_ (_28986_, _10047_, _03520_);
  nor _79436_ (_28987_, _28986_, _28299_);
  nand _79437_ (_28988_, _28987_, _28985_);
  nor _79438_ (_28989_, _28675_, _10851_);
  nor _79439_ (_28990_, _28989_, _03645_);
  and _79440_ (_28991_, _28990_, _28988_);
  or _79441_ (_28993_, _28991_, _28670_);
  nor _79442_ (_28994_, _10862_, _03166_);
  and _79443_ (_28995_, _28994_, _28993_);
  and _79444_ (_28996_, _28675_, _10862_);
  or _79445_ (_28997_, _28996_, _28995_);
  or _79446_ (_28998_, _28997_, _42967_);
  or _79447_ (_28999_, _42963_, \oc8051_golden_model_1.PC [8]);
  and _79448_ (_29000_, _28999_, _41755_);
  and _79449_ (_43337_, _29000_, _28998_);
  nor _79450_ (_29001_, _04284_, _10855_);
  nor _79451_ (_29003_, _04284_, _10832_);
  and _79452_ (_29004_, _28672_, \oc8051_golden_model_1.PC [9]);
  nor _79453_ (_29005_, _28672_, \oc8051_golden_model_1.PC [9]);
  nor _79454_ (_29006_, _29005_, _29004_);
  nor _79455_ (_29007_, _29006_, _09949_);
  nor _79456_ (_29008_, _29006_, _09951_);
  and _79457_ (_29009_, _10156_, _03758_);
  nor _79458_ (_29010_, _29006_, _09956_);
  not _79459_ (_29011_, _29006_);
  and _79460_ (_29012_, _29011_, _10545_);
  and _79461_ (_29014_, _10156_, _03636_);
  nor _79462_ (_29015_, _29006_, _10520_);
  and _79463_ (_29016_, _09995_, _03745_);
  and _79464_ (_29017_, _09995_, _03606_);
  and _79465_ (_29018_, _09995_, _03607_);
  not _79466_ (_29019_, _11596_);
  nand _79467_ (_29020_, _29006_, _04012_);
  nand _79468_ (_29021_, _29011_, _28725_);
  and _79469_ (_29022_, _12260_, _03922_);
  nor _79470_ (_29023_, _29022_, _26577_);
  nor _79471_ (_29025_, _04426_, \oc8051_golden_model_1.PC [9]);
  nand _79472_ (_29026_, _29025_, _10278_);
  nand _79473_ (_29027_, _29026_, _29023_);
  nand _79474_ (_29028_, _29027_, _25909_);
  and _79475_ (_29029_, _29028_, _29021_);
  nor _79476_ (_29030_, _29029_, _05833_);
  and _79477_ (_29031_, _29030_, _29020_);
  and _79478_ (_29032_, _10269_, _09995_);
  nor _79479_ (_29033_, _10051_, _10048_);
  and _79480_ (_29034_, _29033_, _09998_);
  nor _79481_ (_29036_, _29033_, _09998_);
  nor _79482_ (_29037_, _29036_, _29034_);
  nor _79483_ (_29038_, _29037_, _10269_);
  or _79484_ (_29039_, _29038_, _29032_);
  nor _79485_ (_29040_, _29039_, _05831_);
  nor _79486_ (_29041_, _29040_, _29031_);
  nor _79487_ (_29042_, _29041_, _04438_);
  and _79488_ (_29043_, _29011_, _04438_);
  nor _79489_ (_29044_, _29043_, _29042_);
  and _79490_ (_29045_, _29044_, _04444_);
  nor _79491_ (_29047_, _10221_, _10218_);
  and _79492_ (_29048_, _29047_, _10160_);
  nor _79493_ (_29049_, _29047_, _10160_);
  nor _79494_ (_29050_, _29049_, _29048_);
  and _79495_ (_29051_, _29050_, _27991_);
  nor _79496_ (_29052_, _25937_, _10156_);
  or _79497_ (_29053_, _29052_, _04444_);
  nor _79498_ (_29054_, _29053_, _29051_);
  or _79499_ (_29055_, _29054_, _10256_);
  nor _79500_ (_29056_, _29055_, _29045_);
  nor _79501_ (_29058_, _29006_, _10255_);
  nor _79502_ (_29059_, _29058_, _03516_);
  not _79503_ (_29060_, _29059_);
  nor _79504_ (_29061_, _29060_, _29056_);
  and _79505_ (_29062_, _09995_, _03516_);
  or _79506_ (_29063_, _29062_, _04746_);
  nor _79507_ (_29064_, _29063_, _29061_);
  nor _79508_ (_29065_, _29064_, _03568_);
  and _79509_ (_29066_, _09995_, _03568_);
  nor _79510_ (_29067_, _29066_, _26212_);
  not _79511_ (_29069_, _29067_);
  nor _79512_ (_29070_, _29069_, _29065_);
  nor _79513_ (_29071_, _29006_, _10307_);
  nor _79514_ (_29072_, _29071_, _03575_);
  not _79515_ (_29073_, _29072_);
  nor _79516_ (_29074_, _29073_, _29070_);
  and _79517_ (_29075_, _09995_, _03575_);
  nor _79518_ (_29076_, _29075_, _26220_);
  not _79519_ (_29077_, _29076_);
  nor _79520_ (_29078_, _29077_, _29074_);
  nor _79521_ (_29080_, _29006_, _10316_);
  nor _79522_ (_29081_, _29080_, _03512_);
  not _79523_ (_29082_, _29081_);
  nor _79524_ (_29083_, _29082_, _29078_);
  and _79525_ (_29084_, _09995_, _03512_);
  or _79526_ (_29085_, _29084_, _10249_);
  nor _79527_ (_29086_, _29085_, _29083_);
  nor _79528_ (_29087_, _29086_, _03511_);
  and _79529_ (_29088_, _09995_, _03511_);
  nor _79530_ (_29089_, _29088_, _10326_);
  not _79531_ (_29091_, _29089_);
  nor _79532_ (_29092_, _29091_, _29087_);
  and _79533_ (_29093_, _10360_, _10156_);
  nor _79534_ (_29094_, _29050_, _10360_);
  or _79535_ (_29095_, _29094_, _10325_);
  nor _79536_ (_29096_, _29095_, _29093_);
  or _79537_ (_29097_, _29096_, _03657_);
  nor _79538_ (_29098_, _29097_, _29092_);
  and _79539_ (_29099_, _10156_, _10116_);
  nor _79540_ (_29100_, _29050_, _10116_);
  nor _79541_ (_29102_, _29100_, _29099_);
  nor _79542_ (_29103_, _29102_, _11574_);
  nor _79543_ (_29104_, _29103_, _29098_);
  nor _79544_ (_29105_, _29104_, _29019_);
  and _79545_ (_29106_, _10398_, _10156_);
  nor _79546_ (_29107_, _29050_, _10398_);
  or _79547_ (_29108_, _29107_, _29106_);
  and _79548_ (_29109_, _29108_, _03638_);
  nor _79549_ (_29110_, _29050_, _10382_);
  and _79550_ (_29111_, _10382_, _10156_);
  nor _79551_ (_29113_, _29111_, _29110_);
  nor _79552_ (_29114_, _29113_, _03998_);
  nor _79553_ (_29115_, _29114_, _29109_);
  and _79554_ (_29116_, _29006_, _10083_);
  nor _79555_ (_29117_, _29116_, _03505_);
  and _79556_ (_29118_, _29117_, _29115_);
  not _79557_ (_29119_, _29118_);
  nor _79558_ (_29120_, _29119_, _29105_);
  and _79559_ (_29121_, _12260_, _03505_);
  not _79560_ (_29122_, _29121_);
  nand _79561_ (_29124_, _29122_, _28786_);
  or _79562_ (_29125_, _29124_, _29120_);
  nor _79563_ (_29126_, _26281_, _12260_);
  nor _79564_ (_29127_, _29126_, _25991_);
  nand _79565_ (_29128_, _29127_, _29125_);
  nor _79566_ (_29129_, _29006_, _10415_);
  nor _79567_ (_29130_, _29129_, _03607_);
  and _79568_ (_29131_, _29130_, _29128_);
  or _79569_ (_29132_, _29131_, _29018_);
  and _79570_ (_29133_, _29132_, _10421_);
  or _79571_ (_29135_, _29133_, _29017_);
  nand _79572_ (_29136_, _29135_, _10426_);
  nor _79573_ (_29137_, _29011_, _10426_);
  nor _79574_ (_29138_, _29137_, _10431_);
  nand _79575_ (_29139_, _29138_, _29136_);
  nor _79576_ (_29140_, _09995_, _10430_);
  nor _79577_ (_29141_, _29140_, _03311_);
  nand _79578_ (_29142_, _29141_, _29139_);
  nor _79579_ (_29143_, _29011_, _03254_);
  nor _79580_ (_29144_, _29143_, _03499_);
  nand _79581_ (_29146_, _29144_, _29142_);
  nor _79582_ (_29147_, _03632_, _03223_);
  not _79583_ (_29148_, _29147_);
  and _79584_ (_29149_, _12260_, _03499_);
  nor _79585_ (_29150_, _29149_, _29148_);
  nand _79586_ (_29151_, _29150_, _29146_);
  and _79587_ (_29152_, _10156_, _03632_);
  nor _79588_ (_29153_, _29152_, _26322_);
  nand _79589_ (_29154_, _29153_, _29151_);
  nor _79590_ (_29155_, _09995_, _03493_);
  nor _79591_ (_29157_, _29155_, _03221_);
  nand _79592_ (_29158_, _29157_, _29154_);
  and _79593_ (_29159_, _10156_, _03221_);
  nor _79594_ (_29160_, _29159_, _26330_);
  nand _79595_ (_29161_, _29160_, _29158_);
  nor _79596_ (_29162_, _29006_, _10081_);
  nor _79597_ (_29163_, _29162_, _03745_);
  and _79598_ (_29164_, _29163_, _29161_);
  or _79599_ (_29165_, _29164_, _29016_);
  nand _79600_ (_29166_, _29165_, _28686_);
  nor _79601_ (_29168_, _29037_, _10459_);
  nor _79602_ (_29169_, _29168_, _06055_);
  nand _79603_ (_29170_, _29169_, _29166_);
  nor _79604_ (_29171_, _09995_, _05775_);
  nor _79605_ (_29172_, _29171_, _03437_);
  nand _79606_ (_29173_, _29172_, _29170_);
  and _79607_ (_29174_, _10156_, _03437_);
  nor _79608_ (_29175_, _29174_, _08385_);
  nand _79609_ (_29176_, _29175_, _29173_);
  and _79610_ (_29177_, _12260_, _08385_);
  nor _79611_ (_29179_, _29177_, _10472_);
  and _79612_ (_29180_, _29179_, _29176_);
  nor _79613_ (_29181_, _10500_, \oc8051_golden_model_1.DPH [1]);
  not _79614_ (_29182_, _29181_);
  nor _79615_ (_29183_, _10501_, _25897_);
  and _79616_ (_29184_, _29183_, _29182_);
  or _79617_ (_29185_, _29184_, _29180_);
  nand _79618_ (_29186_, _29185_, _04118_);
  and _79619_ (_29187_, _09995_, _03744_);
  nor _79620_ (_29188_, _29187_, _03189_);
  nand _79621_ (_29190_, _29188_, _29186_);
  nand _79622_ (_29191_, _29190_, _10515_);
  and _79623_ (_29192_, _09995_, _08698_);
  nor _79624_ (_29193_, _29037_, _08698_);
  or _79625_ (_29194_, _29193_, _29192_);
  and _79626_ (_29195_, _29194_, _10076_);
  nor _79627_ (_29196_, _29195_, _26754_);
  and _79628_ (_29197_, _29196_, _29191_);
  or _79629_ (_29198_, _29197_, _29015_);
  nand _79630_ (_29199_, _29198_, _10523_);
  nor _79631_ (_29200_, _10523_, _09995_);
  nor _79632_ (_29201_, _29200_, _03636_);
  and _79633_ (_29202_, _29201_, _29199_);
  or _79634_ (_29203_, _29202_, _29014_);
  nand _79635_ (_29204_, _29203_, _04501_);
  and _79636_ (_29205_, _09995_, _03769_);
  nor _79637_ (_29206_, _29205_, _03194_);
  nand _79638_ (_29207_, _29206_, _29204_);
  nand _79639_ (_29208_, _29207_, _10535_);
  and _79640_ (_29209_, _29037_, _08698_);
  nor _79641_ (_29211_, _09995_, _08698_);
  nor _79642_ (_29212_, _29211_, _10535_);
  not _79643_ (_29213_, _29212_);
  nor _79644_ (_29214_, _29213_, _29209_);
  nor _79645_ (_29215_, _29214_, _10545_);
  and _79646_ (_29216_, _29215_, _29208_);
  or _79647_ (_29217_, _29216_, _29012_);
  nand _79648_ (_29218_, _29217_, _10548_);
  nor _79649_ (_29219_, _09995_, _10548_);
  nor _79650_ (_29220_, _29219_, _04504_);
  nand _79651_ (_29222_, _29220_, _29218_);
  nand _79652_ (_29223_, _10156_, _04504_);
  nand _79653_ (_29224_, _29223_, _29222_);
  nand _79654_ (_29225_, _29224_, _03753_);
  and _79655_ (_29226_, _09995_, _03752_);
  nor _79656_ (_29227_, _29226_, _03192_);
  nand _79657_ (_29228_, _29227_, _29225_);
  nand _79658_ (_29229_, _29228_, _09959_);
  and _79659_ (_29230_, _09995_, \oc8051_golden_model_1.PSW [7]);
  nor _79660_ (_29231_, _29037_, \oc8051_golden_model_1.PSW [7]);
  or _79661_ (_29233_, _29231_, _29230_);
  and _79662_ (_29234_, _29233_, _09958_);
  nor _79663_ (_29235_, _29234_, _10560_);
  and _79664_ (_29236_, _29235_, _29229_);
  or _79665_ (_29237_, _29236_, _29010_);
  nand _79666_ (_29238_, _29237_, _08478_);
  nor _79667_ (_29239_, _09995_, _08478_);
  nor _79668_ (_29240_, _29239_, _03758_);
  and _79669_ (_29241_, _29240_, _29238_);
  or _79670_ (_29242_, _29241_, _29009_);
  nand _79671_ (_29244_, _29242_, _04517_);
  and _79672_ (_29245_, _09995_, _03760_);
  nor _79673_ (_29246_, _29245_, _03183_);
  nand _79674_ (_29247_, _29246_, _29244_);
  nand _79675_ (_29248_, _29247_, _10577_);
  and _79676_ (_29249_, _29037_, \oc8051_golden_model_1.PSW [7]);
  nor _79677_ (_29250_, _09995_, \oc8051_golden_model_1.PSW [7]);
  nor _79678_ (_29251_, _29250_, _10577_);
  not _79679_ (_29252_, _29251_);
  nor _79680_ (_29253_, _29252_, _29249_);
  nor _79681_ (_29255_, _29253_, _10581_);
  and _79682_ (_29256_, _29255_, _29248_);
  or _79683_ (_29257_, _29256_, _29008_);
  nand _79684_ (_29258_, _29257_, _08524_);
  nor _79685_ (_29259_, _09995_, _08524_);
  nor _79686_ (_29260_, _29259_, _08555_);
  nand _79687_ (_29261_, _29260_, _29258_);
  and _79688_ (_29262_, _29006_, _08555_);
  nor _79689_ (_29263_, _29262_, _03775_);
  nand _79690_ (_29264_, _29263_, _29261_);
  nor _79691_ (_29266_, _03627_, _03179_);
  not _79692_ (_29267_, _29266_);
  and _79693_ (_29268_, _04603_, _03775_);
  nor _79694_ (_29269_, _29268_, _29267_);
  nand _79695_ (_29270_, _29269_, _29264_);
  nor _79696_ (_29271_, _10794_, _10156_);
  and _79697_ (_29272_, _29050_, _10794_);
  or _79698_ (_29273_, _29272_, _10599_);
  nor _79699_ (_29274_, _29273_, _29271_);
  nor _79700_ (_29275_, _29274_, _10603_);
  and _79701_ (_29277_, _29275_, _29270_);
  or _79702_ (_29278_, _29277_, _29007_);
  nand _79703_ (_29279_, _29278_, _09936_);
  nor _79704_ (_29280_, _09995_, _09936_);
  nor _79705_ (_29281_, _29280_, _07729_);
  nand _79706_ (_29282_, _29281_, _29279_);
  and _79707_ (_29283_, _29006_, _07729_);
  nor _79708_ (_29284_, _29283_, _03522_);
  nand _79709_ (_29285_, _29284_, _29282_);
  and _79710_ (_29286_, _04603_, _03522_);
  nor _79711_ (_29288_, _03628_, _03172_);
  not _79712_ (_29289_, _29288_);
  nor _79713_ (_29290_, _29289_, _29286_);
  nand _79714_ (_29291_, _29290_, _29285_);
  and _79715_ (_29292_, _10794_, _10156_);
  nor _79716_ (_29293_, _29050_, _10794_);
  or _79717_ (_29294_, _29293_, _29292_);
  and _79718_ (_29295_, _29294_, _03628_);
  nor _79719_ (_29296_, _29295_, _10822_);
  nand _79720_ (_29297_, _29296_, _29291_);
  nor _79721_ (_29299_, _29006_, _10821_);
  nor _79722_ (_29300_, _29299_, _03790_);
  nand _79723_ (_29301_, _29300_, _29297_);
  and _79724_ (_29302_, _09995_, _03790_);
  nor _79725_ (_29303_, _29302_, _27228_);
  nand _79726_ (_29304_, _29303_, _29301_);
  nor _79727_ (_29305_, _29006_, _10828_);
  nor _79728_ (_29306_, _29305_, _03641_);
  and _79729_ (_29307_, _29306_, _29304_);
  or _79730_ (_29308_, _29307_, _29003_);
  nand _79731_ (_29310_, _29308_, _28976_);
  and _79732_ (_29311_, _29294_, _03151_);
  nor _79733_ (_29312_, _29311_, _10845_);
  nand _79734_ (_29313_, _29312_, _29310_);
  nor _79735_ (_29314_, _29006_, _10844_);
  nor _79736_ (_29315_, _29314_, _03520_);
  nand _79737_ (_29316_, _29315_, _29313_);
  and _79738_ (_29317_, _09995_, _03520_);
  nor _79739_ (_29318_, _29317_, _28299_);
  nand _79740_ (_29319_, _29318_, _29316_);
  nor _79741_ (_29321_, _29006_, _10851_);
  nor _79742_ (_29322_, _29321_, _03645_);
  and _79743_ (_29323_, _29322_, _29319_);
  or _79744_ (_29324_, _29323_, _29001_);
  and _79745_ (_29325_, _29324_, _28994_);
  and _79746_ (_29326_, _29006_, _10862_);
  or _79747_ (_29327_, _29326_, _29325_);
  or _79748_ (_29328_, _29327_, _42967_);
  or _79749_ (_29329_, _42963_, \oc8051_golden_model_1.PC [9]);
  and _79750_ (_29330_, _29329_, _41755_);
  and _79751_ (_43338_, _29330_, _29328_);
  and _79752_ (_29332_, _29004_, \oc8051_golden_model_1.PC [10]);
  nor _79753_ (_29333_, _29004_, \oc8051_golden_model_1.PC [10]);
  nor _79754_ (_29334_, _29333_, _29332_);
  and _79755_ (_29335_, _29334_, _10862_);
  and _79756_ (_29336_, _03877_, _03645_);
  nor _79757_ (_29337_, _29334_, _10844_);
  and _79758_ (_29338_, _03877_, _03641_);
  not _79759_ (_29339_, _29334_);
  and _79760_ (_29340_, _29339_, _07729_);
  and _79761_ (_29342_, _29339_, _08555_);
  and _79762_ (_29343_, _10143_, _03758_);
  and _79763_ (_29344_, _10143_, _03636_);
  nor _79764_ (_29345_, _10076_, _03189_);
  nor _79765_ (_29346_, _29339_, _10426_);
  and _79766_ (_29347_, _29334_, _10083_);
  and _79767_ (_29348_, _10398_, _10142_);
  not _79768_ (_29349_, _10153_);
  nor _79769_ (_29350_, _10225_, _10222_);
  nor _79770_ (_29351_, _29350_, _29349_);
  and _79771_ (_29353_, _29350_, _29349_);
  nor _79772_ (_29354_, _29353_, _29351_);
  and _79773_ (_29355_, _29354_, _10399_);
  or _79774_ (_29356_, _29355_, _29348_);
  and _79775_ (_29357_, _29356_, _03638_);
  nand _79776_ (_29358_, _10382_, _10143_);
  or _79777_ (_29359_, _29354_, _10382_);
  and _79778_ (_29360_, _29359_, _03527_);
  and _79779_ (_29361_, _29360_, _29358_);
  or _79780_ (_29362_, _29361_, _29357_);
  or _79781_ (_29364_, _29362_, _29347_);
  nor _79782_ (_29365_, _29339_, _10316_);
  nor _79783_ (_29366_, _29334_, _10307_);
  nor _79784_ (_29367_, _29339_, _10303_);
  or _79785_ (_29368_, _29354_, _10261_);
  nand _79786_ (_29369_, _10261_, _10143_);
  and _79787_ (_29370_, _29369_, _03570_);
  and _79788_ (_29371_, _29370_, _29368_);
  and _79789_ (_29372_, _10269_, _09989_);
  not _79790_ (_29373_, _09992_);
  nor _79791_ (_29375_, _10055_, _10052_);
  nor _79792_ (_29376_, _29375_, _29373_);
  and _79793_ (_29377_, _29375_, _29373_);
  nor _79794_ (_29378_, _29377_, _29376_);
  and _79795_ (_29379_, _29378_, _10271_);
  nor _79796_ (_29380_, _29379_, _29372_);
  nand _79797_ (_29381_, _29380_, _05833_);
  and _79798_ (_29382_, _25905_, _10290_);
  nor _79799_ (_29383_, _29382_, _29334_);
  and _79800_ (_29384_, _12464_, _03922_);
  nor _79801_ (_29386_, _04426_, \oc8051_golden_model_1.PC [10]);
  and _79802_ (_29387_, _29386_, _10278_);
  or _79803_ (_29388_, _29387_, _29384_);
  and _79804_ (_29389_, _29388_, _26578_);
  or _79805_ (_29390_, _29389_, _29383_);
  nor _79806_ (_29391_, _29339_, _10290_);
  or _79807_ (_29392_, _05833_, _03923_);
  nor _79808_ (_29393_, _29392_, _29391_);
  and _79809_ (_29394_, _29393_, _29390_);
  nor _79810_ (_29395_, _29394_, _10297_);
  and _79811_ (_29397_, _29395_, _29381_);
  or _79812_ (_29398_, _29397_, _29371_);
  and _79813_ (_29399_, _29398_, _10255_);
  or _79814_ (_29400_, _29399_, _29367_);
  and _79815_ (_29401_, _29400_, _03576_);
  nor _79816_ (_29402_, _12464_, _03576_);
  nor _79817_ (_29403_, _29402_, _04746_);
  nand _79818_ (_29404_, _29403_, _10307_);
  nor _79819_ (_29405_, _29404_, _29401_);
  or _79820_ (_29406_, _29405_, _29366_);
  nand _79821_ (_29408_, _29406_, _03583_);
  and _79822_ (_29409_, _12464_, _03575_);
  nor _79823_ (_29410_, _29409_, _26220_);
  and _79824_ (_29411_, _29410_, _29408_);
  or _79825_ (_29412_, _29411_, _29365_);
  nand _79826_ (_29413_, _29412_, _03513_);
  and _79827_ (_29414_, _09989_, _03512_);
  nor _79828_ (_29415_, _29414_, _10249_);
  nand _79829_ (_29416_, _29415_, _29413_);
  nand _79830_ (_29417_, _29416_, _04887_);
  and _79831_ (_29419_, _09989_, _03511_);
  nor _79832_ (_29420_, _29419_, _10326_);
  nand _79833_ (_29421_, _29420_, _29417_);
  and _79834_ (_29422_, _10360_, _10142_);
  not _79835_ (_29423_, _29354_);
  nor _79836_ (_29424_, _29423_, _10360_);
  or _79837_ (_29425_, _29424_, _10325_);
  nor _79838_ (_29426_, _29425_, _29422_);
  nor _79839_ (_29427_, _29426_, _03657_);
  nand _79840_ (_29428_, _29427_, _29421_);
  nor _79841_ (_29430_, _29423_, _10116_);
  and _79842_ (_29431_, _10142_, _10116_);
  nor _79843_ (_29432_, _29431_, _29430_);
  or _79844_ (_29433_, _29432_, _10328_);
  nand _79845_ (_29434_, _29433_, _29428_);
  and _79846_ (_29435_, _29434_, _11596_);
  or _79847_ (_29436_, _29435_, _29364_);
  and _79848_ (_29437_, _26281_, _03506_);
  and _79849_ (_29438_, _29437_, _29436_);
  nor _79850_ (_29439_, _29437_, _12464_);
  nand _79851_ (_29441_, _10415_, _03200_);
  or _79852_ (_29442_, _29441_, _29439_);
  or _79853_ (_29443_, _29442_, _29438_);
  nor _79854_ (_29444_, _29334_, _10415_);
  nor _79855_ (_29445_, _29444_, _03607_);
  and _79856_ (_29446_, _29445_, _29443_);
  and _79857_ (_29447_, _09989_, _03607_);
  nor _79858_ (_29448_, _29447_, _29446_);
  nand _79859_ (_29449_, _29448_, _10421_);
  and _79860_ (_29450_, _12464_, _03606_);
  nor _79861_ (_29452_, _29450_, _26302_);
  and _79862_ (_29453_, _29452_, _29449_);
  nor _79863_ (_29454_, _29453_, _29346_);
  or _79864_ (_29455_, _29454_, _10431_);
  or _79865_ (_29456_, _12464_, _10430_);
  and _79866_ (_29457_, _29456_, _03254_);
  nand _79867_ (_29458_, _29457_, _29455_);
  nor _79868_ (_29459_, _29334_, _03254_);
  nor _79869_ (_29460_, _29459_, _03499_);
  and _79870_ (_29461_, _29460_, _29458_);
  and _79871_ (_29463_, _09989_, _03499_);
  nor _79872_ (_29464_, _29463_, _29461_);
  and _79873_ (_29465_, _29464_, _29147_);
  and _79874_ (_29466_, _10143_, _03632_);
  or _79875_ (_29467_, _29466_, _29465_);
  and _79876_ (_29468_, _29467_, _03493_);
  nor _79877_ (_29469_, _09989_, _03493_);
  or _79878_ (_29470_, _29469_, _29468_);
  nand _79879_ (_29471_, _29470_, _03474_);
  and _79880_ (_29472_, _10143_, _03221_);
  nor _79881_ (_29474_, _29472_, _26330_);
  and _79882_ (_29475_, _29474_, _29471_);
  nor _79883_ (_29476_, _29339_, _10081_);
  or _79884_ (_29477_, _29476_, _29475_);
  nand _79885_ (_29478_, _29477_, _27421_);
  and _79886_ (_29479_, _09989_, _03745_);
  nor _79887_ (_29480_, _29479_, _28687_);
  nand _79888_ (_29481_, _29480_, _29478_);
  nor _79889_ (_29482_, _29378_, _10459_);
  nor _79890_ (_29483_, _29482_, _06055_);
  and _79891_ (_29485_, _29483_, _29481_);
  nor _79892_ (_29486_, _12464_, _05775_);
  or _79893_ (_29487_, _29486_, _03437_);
  or _79894_ (_29488_, _29487_, _29485_);
  and _79895_ (_29489_, _10143_, _03437_);
  nor _79896_ (_29490_, _29489_, _08385_);
  nand _79897_ (_29491_, _29490_, _29488_);
  and _79898_ (_29492_, _09989_, _08385_);
  nor _79899_ (_29493_, _29492_, _10472_);
  nand _79900_ (_29494_, _29493_, _29491_);
  nor _79901_ (_29496_, _10501_, \oc8051_golden_model_1.DPH [2]);
  nor _79902_ (_29497_, _29496_, _10502_);
  nor _79903_ (_29498_, _29497_, _25897_);
  nor _79904_ (_29499_, _29498_, _03744_);
  and _79905_ (_29500_, _29499_, _29494_);
  and _79906_ (_29501_, _09989_, _03744_);
  or _79907_ (_29502_, _29501_, _29500_);
  nand _79908_ (_29503_, _29502_, _29345_);
  nor _79909_ (_29504_, _29378_, _08698_);
  or _79910_ (_29505_, _09989_, _10077_);
  nand _79911_ (_29507_, _29505_, _10076_);
  or _79912_ (_29508_, _29507_, _29504_);
  and _79913_ (_29509_, _29508_, _10520_);
  nand _79914_ (_29510_, _29509_, _29503_);
  nor _79915_ (_29511_, _29334_, _10520_);
  nor _79916_ (_29512_, _29511_, _10524_);
  nand _79917_ (_29513_, _29512_, _29510_);
  nor _79918_ (_29514_, _10523_, _12464_);
  nor _79919_ (_29515_, _29514_, _03636_);
  and _79920_ (_29516_, _29515_, _29513_);
  or _79921_ (_29517_, _29516_, _29344_);
  or _79922_ (_29518_, _29517_, _03769_);
  nand _79923_ (_29519_, _09989_, _03769_);
  and _79924_ (_29520_, _29519_, _29518_);
  or _79925_ (_29521_, _29520_, _03194_);
  or _79926_ (_29522_, _29521_, _10534_);
  nor _79927_ (_29523_, _29378_, _10077_);
  nor _79928_ (_29524_, _09989_, _08698_);
  nor _79929_ (_29525_, _29524_, _10535_);
  not _79930_ (_29526_, _29525_);
  nor _79931_ (_29529_, _29526_, _29523_);
  nor _79932_ (_29530_, _29529_, _10545_);
  nand _79933_ (_29531_, _29530_, _29522_);
  and _79934_ (_29532_, _29339_, _10545_);
  nor _79935_ (_29533_, _29532_, _10549_);
  nand _79936_ (_29534_, _29533_, _29531_);
  nor _79937_ (_29535_, _12464_, _10548_);
  nor _79938_ (_29536_, _29535_, _04504_);
  nand _79939_ (_29537_, _29536_, _29534_);
  nand _79940_ (_29538_, _10143_, _04504_);
  nand _79941_ (_29540_, _29538_, _29537_);
  nand _79942_ (_29541_, _29540_, _03753_);
  and _79943_ (_29542_, _12464_, _03752_);
  nor _79944_ (_29543_, _29542_, _28898_);
  nand _79945_ (_29544_, _29543_, _29541_);
  and _79946_ (_29545_, _09989_, \oc8051_golden_model_1.PSW [7]);
  and _79947_ (_29546_, _29378_, _07888_);
  or _79948_ (_29547_, _29546_, _29545_);
  and _79949_ (_29548_, _29547_, _09958_);
  nor _79950_ (_29549_, _29548_, _10560_);
  nand _79951_ (_29551_, _29549_, _29544_);
  nor _79952_ (_29552_, _29334_, _09956_);
  nor _79953_ (_29553_, _29552_, _08479_);
  nand _79954_ (_29554_, _29553_, _29551_);
  nor _79955_ (_29555_, _12464_, _08478_);
  nor _79956_ (_29556_, _29555_, _03758_);
  and _79957_ (_29557_, _29556_, _29554_);
  or _79958_ (_29558_, _29557_, _29343_);
  nand _79959_ (_29559_, _29558_, _04517_);
  and _79960_ (_29560_, _12464_, _03760_);
  nor _79961_ (_29562_, _29560_, _26078_);
  nand _79962_ (_29563_, _29562_, _29559_);
  nor _79963_ (_29564_, _29378_, _07888_);
  nor _79964_ (_29565_, _09989_, \oc8051_golden_model_1.PSW [7]);
  nor _79965_ (_29566_, _29565_, _10577_);
  not _79966_ (_29567_, _29566_);
  nor _79967_ (_29568_, _29567_, _29564_);
  nor _79968_ (_29569_, _29568_, _10581_);
  nand _79969_ (_29570_, _29569_, _29563_);
  nor _79970_ (_29571_, _29334_, _09951_);
  nor _79971_ (_29573_, _29571_, _08525_);
  nand _79972_ (_29574_, _29573_, _29570_);
  nor _79973_ (_29575_, _12464_, _08524_);
  nor _79974_ (_29576_, _29575_, _08555_);
  and _79975_ (_29577_, _29576_, _29574_);
  or _79976_ (_29578_, _29577_, _29342_);
  nand _79977_ (_29579_, _29578_, _11403_);
  and _79978_ (_29580_, _05026_, _03775_);
  nor _79979_ (_29581_, _29580_, _29267_);
  nand _79980_ (_29582_, _29581_, _29579_);
  and _79981_ (_29584_, _29423_, _10794_);
  nor _79982_ (_29585_, _10794_, _10142_);
  or _79983_ (_29586_, _29585_, _10599_);
  nor _79984_ (_29587_, _29586_, _29584_);
  nor _79985_ (_29588_, _29587_, _10603_);
  nand _79986_ (_29589_, _29588_, _29582_);
  nor _79987_ (_29590_, _29334_, _09949_);
  nor _79988_ (_29591_, _29590_, _09937_);
  nand _79989_ (_29592_, _29591_, _29589_);
  nor _79990_ (_29593_, _12464_, _09936_);
  nor _79991_ (_29595_, _29593_, _07729_);
  and _79992_ (_29596_, _29595_, _29592_);
  or _79993_ (_29597_, _29596_, _29340_);
  nand _79994_ (_29598_, _29597_, _03523_);
  and _79995_ (_29599_, _05026_, _03522_);
  nor _79996_ (_29600_, _29599_, _29289_);
  nand _79997_ (_29601_, _29600_, _29598_);
  and _79998_ (_29602_, _10794_, _10143_);
  nor _79999_ (_29603_, _29354_, _10794_);
  nor _80000_ (_29604_, _29603_, _29602_);
  and _80001_ (_29606_, _29604_, _03628_);
  nor _80002_ (_29607_, _29606_, _10822_);
  and _80003_ (_29608_, _29607_, _29601_);
  nor _80004_ (_29609_, _29334_, _10821_);
  or _80005_ (_29610_, _29609_, _29608_);
  nand _80006_ (_29611_, _29610_, _04192_);
  and _80007_ (_29612_, _12464_, _03790_);
  nor _80008_ (_29613_, _29612_, _27228_);
  nand _80009_ (_29614_, _29613_, _29611_);
  nor _80010_ (_29615_, _29339_, _10828_);
  nor _80011_ (_29617_, _29615_, _03641_);
  nand _80012_ (_29618_, _29617_, _29614_);
  nand _80013_ (_29619_, _29618_, _28976_);
  or _80014_ (_29620_, _29619_, _29338_);
  and _80015_ (_29621_, _29604_, _03151_);
  nor _80016_ (_29622_, _29621_, _10845_);
  and _80017_ (_29623_, _29622_, _29620_);
  or _80018_ (_29624_, _29623_, _29337_);
  nand _80019_ (_29625_, _29624_, _03521_);
  and _80020_ (_29626_, _12464_, _03520_);
  nor _80021_ (_29628_, _29626_, _28299_);
  nand _80022_ (_29629_, _29628_, _29625_);
  nor _80023_ (_29630_, _29339_, _10851_);
  nor _80024_ (_29631_, _29630_, _03645_);
  nand _80025_ (_29632_, _29631_, _29629_);
  nand _80026_ (_29633_, _29632_, _28994_);
  nor _80027_ (_29634_, _29633_, _29336_);
  or _80028_ (_29635_, _29634_, _29335_);
  or _80029_ (_29636_, _29635_, _42967_);
  or _80030_ (_29637_, _42963_, \oc8051_golden_model_1.PC [10]);
  and _80031_ (_29639_, _29637_, _41755_);
  and _80032_ (_43339_, _29639_, _29636_);
  and _80033_ (_29640_, _29332_, \oc8051_golden_model_1.PC [11]);
  nor _80034_ (_29641_, _29332_, \oc8051_golden_model_1.PC [11]);
  nor _80035_ (_29642_, _29641_, _29640_);
  or _80036_ (_29643_, _29642_, _09949_);
  or _80037_ (_29644_, _29642_, _09951_);
  or _80038_ (_29645_, _10573_, _09984_);
  and _80039_ (_29646_, _29645_, _10577_);
  or _80040_ (_29647_, _29642_, _09956_);
  or _80041_ (_29649_, _09984_, _09960_);
  and _80042_ (_29650_, _29649_, _09959_);
  or _80043_ (_29651_, _29642_, _10520_);
  or _80044_ (_29652_, _09984_, _05775_);
  and _80045_ (_29653_, _10147_, _03221_);
  or _80046_ (_29654_, _29642_, _10426_);
  and _80047_ (_29655_, _29642_, _25991_);
  nor _80048_ (_29656_, _29351_, _10144_);
  and _80049_ (_29657_, _29656_, _10151_);
  nor _80050_ (_29658_, _29656_, _10151_);
  nor _80051_ (_29660_, _29658_, _29657_);
  nor _80052_ (_29661_, _29660_, _10116_);
  and _80053_ (_29662_, _10147_, _10116_);
  or _80054_ (_29663_, _29662_, _29661_);
  and _80055_ (_29664_, _29663_, _03657_);
  and _80056_ (_29665_, _09984_, _03575_);
  not _80057_ (_29666_, _29660_);
  or _80058_ (_29667_, _29666_, _10261_);
  nand _80059_ (_29668_, _10261_, _10148_);
  and _80060_ (_29669_, _29668_, _29667_);
  or _80061_ (_29671_, _29669_, _04444_);
  and _80062_ (_29672_, _10269_, _09984_);
  nor _80063_ (_29673_, _29376_, _09990_);
  and _80064_ (_29674_, _29673_, _09987_);
  nor _80065_ (_29675_, _29673_, _09987_);
  or _80066_ (_29676_, _29675_, _29674_);
  and _80067_ (_29677_, _29676_, _10271_);
  or _80068_ (_29678_, _29677_, _29672_);
  or _80069_ (_29679_, _29678_, _05831_);
  or _80070_ (_29680_, _27282_, \oc8051_golden_model_1.PC [11]);
  and _80071_ (_29682_, _29680_, _04427_);
  and _80072_ (_29683_, _09984_, _04426_);
  or _80073_ (_29684_, _29683_, _26577_);
  or _80074_ (_29685_, _29684_, _29682_);
  or _80075_ (_29686_, _29642_, _25905_);
  and _80076_ (_29687_, _29686_, _25909_);
  and _80077_ (_29688_, _29687_, _29685_);
  and _80078_ (_29689_, _09984_, _03923_);
  and _80079_ (_29690_, _29642_, _27661_);
  or _80080_ (_29691_, _29690_, _05833_);
  or _80081_ (_29693_, _29691_, _29689_);
  or _80082_ (_29694_, _29693_, _29688_);
  and _80083_ (_29695_, _29694_, _05847_);
  and _80084_ (_29696_, _29695_, _29679_);
  and _80085_ (_29697_, _29642_, _04438_);
  or _80086_ (_29698_, _29697_, _03570_);
  or _80087_ (_29699_, _29698_, _29696_);
  and _80088_ (_29700_, _29699_, _29671_);
  or _80089_ (_29701_, _29700_, _10256_);
  or _80090_ (_29702_, _29642_, _10255_);
  and _80091_ (_29704_, _29702_, _10302_);
  and _80092_ (_29705_, _29704_, _29701_);
  not _80093_ (_29706_, _10302_);
  nand _80094_ (_29707_, _29706_, _09984_);
  nand _80095_ (_29708_, _29707_, _10307_);
  or _80096_ (_29709_, _29708_, _29705_);
  or _80097_ (_29710_, _29642_, _10307_);
  and _80098_ (_29711_, _29710_, _03583_);
  and _80099_ (_29712_, _29711_, _29709_);
  or _80100_ (_29713_, _29712_, _29665_);
  and _80101_ (_29715_, _29713_, _10316_);
  not _80102_ (_29716_, _10251_);
  and _80103_ (_29717_, _29642_, _26220_);
  or _80104_ (_29718_, _29717_, _29716_);
  or _80105_ (_29719_, _29718_, _29715_);
  or _80106_ (_29720_, _10251_, _09984_);
  and _80107_ (_29721_, _29720_, _29719_);
  or _80108_ (_29722_, _29721_, _10326_);
  and _80109_ (_29723_, _10360_, _10147_);
  nor _80110_ (_29724_, _29660_, _10360_);
  or _80111_ (_29726_, _29724_, _29723_);
  or _80112_ (_29727_, _29726_, _10325_);
  and _80113_ (_29728_, _29727_, _10328_);
  and _80114_ (_29729_, _29728_, _29722_);
  or _80115_ (_29730_, _29729_, _29664_);
  and _80116_ (_29731_, _29730_, _11596_);
  nand _80117_ (_29732_, _29660_, _10399_);
  nand _80118_ (_29733_, _10398_, _10148_);
  and _80119_ (_29734_, _29733_, _03638_);
  and _80120_ (_29735_, _29734_, _29732_);
  or _80121_ (_29737_, _29666_, _10382_);
  nand _80122_ (_29738_, _10382_, _10148_);
  and _80123_ (_29739_, _29738_, _03527_);
  and _80124_ (_29740_, _29739_, _29737_);
  or _80125_ (_29741_, _29740_, _29735_);
  nand _80126_ (_29742_, _29642_, _10083_);
  nand _80127_ (_29743_, _29742_, _10408_);
  or _80128_ (_29744_, _29743_, _29741_);
  or _80129_ (_29745_, _29744_, _29731_);
  or _80130_ (_29746_, _10408_, _09984_);
  and _80131_ (_29748_, _29746_, _10415_);
  and _80132_ (_29749_, _29748_, _29745_);
  or _80133_ (_29750_, _29749_, _29655_);
  and _80134_ (_29751_, _29750_, _10422_);
  and _80135_ (_29752_, _10423_, _09984_);
  or _80136_ (_29753_, _29752_, _26302_);
  or _80137_ (_29754_, _29753_, _29751_);
  and _80138_ (_29755_, _29754_, _29654_);
  or _80139_ (_29756_, _29755_, _10431_);
  or _80140_ (_29757_, _09984_, _10430_);
  and _80141_ (_29759_, _29757_, _03254_);
  and _80142_ (_29760_, _29759_, _29756_);
  nand _80143_ (_29761_, _29642_, _03311_);
  nand _80144_ (_29762_, _29761_, _10439_);
  or _80145_ (_29763_, _29762_, _29760_);
  or _80146_ (_29764_, _10439_, _09984_);
  and _80147_ (_29765_, _29764_, _09755_);
  and _80148_ (_29766_, _29765_, _29763_);
  nand _80149_ (_29767_, _10147_, _03632_);
  nand _80150_ (_29768_, _29767_, _03493_);
  or _80151_ (_29770_, _29768_, _29766_);
  or _80152_ (_29771_, _09984_, _03493_);
  and _80153_ (_29772_, _29771_, _03474_);
  and _80154_ (_29773_, _29772_, _29770_);
  or _80155_ (_29774_, _29773_, _29653_);
  and _80156_ (_29775_, _29774_, _10081_);
  and _80157_ (_29776_, _29642_, _26330_);
  or _80158_ (_29777_, _29776_, _10454_);
  or _80159_ (_29778_, _29777_, _29775_);
  or _80160_ (_29779_, _10453_, _09984_);
  and _80161_ (_29780_, _29779_, _10459_);
  and _80162_ (_29781_, _29780_, _29778_);
  and _80163_ (_29782_, _29676_, _10458_);
  or _80164_ (_29783_, _29782_, _06055_);
  or _80165_ (_29784_, _29783_, _29781_);
  and _80166_ (_29785_, _29784_, _29652_);
  or _80167_ (_29786_, _29785_, _03437_);
  nand _80168_ (_29787_, _10148_, _03437_);
  and _80169_ (_29788_, _29787_, _08386_);
  and _80170_ (_29789_, _29788_, _29786_);
  and _80171_ (_29792_, _09984_, _08385_);
  or _80172_ (_29793_, _29792_, _29789_);
  and _80173_ (_29794_, _29793_, _25897_);
  or _80174_ (_29795_, _10502_, \oc8051_golden_model_1.DPH [3]);
  nor _80175_ (_29796_, _10503_, _25897_);
  and _80176_ (_29797_, _29796_, _29795_);
  or _80177_ (_29798_, _29797_, _10512_);
  or _80178_ (_29799_, _29798_, _29794_);
  or _80179_ (_29800_, _10511_, _09984_);
  and _80180_ (_29801_, _29800_, _10515_);
  and _80181_ (_29803_, _29801_, _29799_);
  or _80182_ (_29804_, _29676_, _08698_);
  or _80183_ (_29805_, _09984_, _10077_);
  and _80184_ (_29806_, _29805_, _10076_);
  and _80185_ (_29807_, _29806_, _29804_);
  or _80186_ (_29808_, _29807_, _26754_);
  or _80187_ (_29809_, _29808_, _29803_);
  and _80188_ (_29810_, _29809_, _29651_);
  or _80189_ (_29811_, _29810_, _10524_);
  or _80190_ (_29812_, _10523_, _09984_);
  and _80191_ (_29814_, _29812_, _04499_);
  and _80192_ (_29815_, _29814_, _29811_);
  nand _80193_ (_29816_, _10147_, _03636_);
  nand _80194_ (_29817_, _29816_, _10531_);
  or _80195_ (_29818_, _29817_, _29815_);
  or _80196_ (_29819_, _10531_, _09984_);
  and _80197_ (_29820_, _29819_, _10535_);
  and _80198_ (_29821_, _29820_, _29818_);
  or _80199_ (_29822_, _29676_, _10077_);
  or _80200_ (_29823_, _09984_, _08698_);
  and _80201_ (_29825_, _29823_, _10534_);
  and _80202_ (_29826_, _29825_, _29822_);
  or _80203_ (_29827_, _29826_, _29821_);
  and _80204_ (_29828_, _29827_, _10546_);
  and _80205_ (_29829_, _29642_, _10545_);
  or _80206_ (_29830_, _29829_, _10549_);
  or _80207_ (_29831_, _29830_, _29828_);
  or _80208_ (_29832_, _09984_, _10548_);
  and _80209_ (_29833_, _29832_, _05769_);
  and _80210_ (_29834_, _29833_, _29831_);
  nand _80211_ (_29836_, _10147_, _03754_);
  nand _80212_ (_29837_, _29836_, _09960_);
  or _80213_ (_29838_, _29837_, _29834_);
  and _80214_ (_29839_, _29838_, _29650_);
  or _80215_ (_29840_, _29676_, \oc8051_golden_model_1.PSW [7]);
  or _80216_ (_29841_, _09984_, _07888_);
  and _80217_ (_29842_, _29841_, _09958_);
  and _80218_ (_29843_, _29842_, _29840_);
  or _80219_ (_29844_, _29843_, _10560_);
  or _80220_ (_29845_, _29844_, _29839_);
  and _80221_ (_29847_, _29845_, _29647_);
  or _80222_ (_29848_, _29847_, _08479_);
  or _80223_ (_29849_, _09984_, _08478_);
  and _80224_ (_29850_, _29849_, _03759_);
  and _80225_ (_29851_, _29850_, _29848_);
  nand _80226_ (_29852_, _10147_, _03758_);
  nand _80227_ (_29853_, _29852_, _10573_);
  or _80228_ (_29854_, _29853_, _29851_);
  and _80229_ (_29855_, _29854_, _29646_);
  or _80230_ (_29856_, _29676_, _07888_);
  or _80231_ (_29858_, _09984_, \oc8051_golden_model_1.PSW [7]);
  and _80232_ (_29859_, _29858_, _10576_);
  and _80233_ (_29860_, _29859_, _29856_);
  or _80234_ (_29861_, _29860_, _10581_);
  or _80235_ (_29862_, _29861_, _29855_);
  and _80236_ (_29863_, _29862_, _29644_);
  or _80237_ (_29864_, _29863_, _08525_);
  or _80238_ (_29865_, _09984_, _08524_);
  and _80239_ (_29866_, _29865_, _08556_);
  and _80240_ (_29867_, _29866_, _29864_);
  and _80241_ (_29869_, _29642_, _08555_);
  or _80242_ (_29870_, _29869_, _03775_);
  or _80243_ (_29871_, _29870_, _29867_);
  nand _80244_ (_29872_, _04843_, _03775_);
  and _80245_ (_29873_, _29872_, _29871_);
  or _80246_ (_29874_, _29873_, _03179_);
  or _80247_ (_29875_, _09984_, _06328_);
  and _80248_ (_29876_, _29875_, _10599_);
  and _80249_ (_29877_, _29876_, _29874_);
  nand _80250_ (_29878_, _29660_, _10794_);
  or _80251_ (_29880_, _10794_, _10147_);
  and _80252_ (_29881_, _29880_, _03627_);
  and _80253_ (_29882_, _29881_, _29878_);
  or _80254_ (_29883_, _29882_, _10603_);
  or _80255_ (_29884_, _29883_, _29877_);
  and _80256_ (_29885_, _29884_, _29643_);
  or _80257_ (_29886_, _29885_, _09937_);
  or _80258_ (_29887_, _09984_, _09936_);
  and _80259_ (_29888_, _29887_, _10803_);
  and _80260_ (_29889_, _29888_, _29886_);
  and _80261_ (_29891_, _29642_, _07729_);
  or _80262_ (_29892_, _29891_, _03522_);
  or _80263_ (_29893_, _29892_, _29889_);
  nand _80264_ (_29894_, _04843_, _03522_);
  and _80265_ (_29895_, _29894_, _29893_);
  or _80266_ (_29896_, _29895_, _03172_);
  or _80267_ (_29897_, _09984_, _25887_);
  and _80268_ (_29898_, _29897_, _03791_);
  and _80269_ (_29899_, _29898_, _29896_);
  or _80270_ (_29900_, _29666_, _10794_);
  nand _80271_ (_29902_, _10794_, _10148_);
  and _80272_ (_29903_, _29902_, _29900_);
  and _80273_ (_29904_, _29903_, _03628_);
  or _80274_ (_29905_, _29904_, _10822_);
  or _80275_ (_29906_, _29905_, _29899_);
  or _80276_ (_29907_, _29642_, _10821_);
  and _80277_ (_29908_, _29907_, _04192_);
  and _80278_ (_29909_, _29908_, _29906_);
  nand _80279_ (_29910_, _09984_, _03790_);
  nand _80280_ (_29911_, _29910_, _10828_);
  or _80281_ (_29912_, _29911_, _29909_);
  or _80282_ (_29913_, _29642_, _10828_);
  and _80283_ (_29914_, _29913_, _10832_);
  and _80284_ (_29915_, _29914_, _29912_);
  nor _80285_ (_29916_, _10832_, _03432_);
  or _80286_ (_29917_, _29916_, _03160_);
  or _80287_ (_29918_, _29917_, _29915_);
  or _80288_ (_29919_, _09984_, _03161_);
  and _80289_ (_29920_, _29919_, _03152_);
  and _80290_ (_29921_, _29920_, _29918_);
  and _80291_ (_29923_, _29903_, _03151_);
  or _80292_ (_29924_, _29923_, _10845_);
  or _80293_ (_29925_, _29924_, _29921_);
  or _80294_ (_29926_, _29642_, _10844_);
  and _80295_ (_29927_, _29926_, _03521_);
  and _80296_ (_29928_, _29927_, _29925_);
  nand _80297_ (_29929_, _09984_, _03520_);
  nand _80298_ (_29930_, _29929_, _10851_);
  or _80299_ (_29931_, _29930_, _29928_);
  or _80300_ (_29932_, _29642_, _10851_);
  and _80301_ (_29934_, _29932_, _10855_);
  and _80302_ (_29935_, _29934_, _29931_);
  not _80303_ (_29936_, _03166_);
  nand _80304_ (_29937_, _03432_, _29936_);
  and _80305_ (_29938_, _29937_, _25883_);
  or _80306_ (_29939_, _29938_, _29935_);
  or _80307_ (_29940_, _09984_, _29936_);
  and _80308_ (_29941_, _29940_, _10863_);
  and _80309_ (_29942_, _29941_, _29939_);
  and _80310_ (_29943_, _29642_, _10862_);
  or _80311_ (_29945_, _29943_, _29942_);
  or _80312_ (_29946_, _29945_, _42967_);
  or _80313_ (_29947_, _42963_, \oc8051_golden_model_1.PC [11]);
  and _80314_ (_29948_, _29947_, _41755_);
  and _80315_ (_43340_, _29948_, _29946_);
  and _80316_ (_29949_, _29640_, \oc8051_golden_model_1.PC [12]);
  nor _80317_ (_29950_, _29640_, \oc8051_golden_model_1.PC [12]);
  nor _80318_ (_29951_, _29950_, _29949_);
  not _80319_ (_29952_, _29951_);
  and _80320_ (_29953_, _29952_, _07729_);
  nor _80321_ (_29955_, _10573_, _12901_);
  nor _80322_ (_29956_, _12901_, _09960_);
  nor _80323_ (_29957_, _10531_, _12901_);
  nor _80324_ (_29958_, _10511_, _12901_);
  nor _80325_ (_29959_, _10408_, _09981_);
  nor _80326_ (_29960_, _29952_, _10316_);
  nor _80327_ (_29961_, _29951_, _10307_);
  and _80328_ (_29962_, _10261_, _10139_);
  and _80329_ (_29963_, _10232_, _10229_);
  nor _80330_ (_29964_, _29963_, _10233_);
  nor _80331_ (_29966_, _29964_, _10261_);
  nor _80332_ (_29967_, _29966_, _29962_);
  or _80333_ (_29968_, _29967_, _04444_);
  and _80334_ (_29969_, _10269_, _09981_);
  and _80335_ (_29970_, _10062_, _10059_);
  nor _80336_ (_29971_, _29970_, _10063_);
  and _80337_ (_29972_, _29971_, _10271_);
  or _80338_ (_29973_, _29972_, _05831_);
  nor _80339_ (_29974_, _29973_, _29969_);
  nor _80340_ (_29975_, _29952_, _29382_);
  not _80341_ (_29977_, _29975_);
  and _80342_ (_29978_, _09981_, _03923_);
  not _80343_ (_29979_, _29978_);
  and _80344_ (_29980_, _09981_, _04426_);
  and _80345_ (_29981_, _04427_, \oc8051_golden_model_1.PC [12]);
  and _80346_ (_29982_, _29981_, _10278_);
  nor _80347_ (_29983_, _29982_, _29980_);
  nor _80348_ (_29984_, _29983_, _26577_);
  and _80349_ (_29985_, _29984_, _25909_);
  nor _80350_ (_29986_, _29985_, _05833_);
  and _80351_ (_29988_, _29986_, _29979_);
  and _80352_ (_29989_, _29988_, _29977_);
  nor _80353_ (_29990_, _29989_, _04438_);
  not _80354_ (_29991_, _29990_);
  nor _80355_ (_29992_, _29991_, _29974_);
  and _80356_ (_29993_, _29951_, _04438_);
  or _80357_ (_29994_, _29993_, _03570_);
  or _80358_ (_29995_, _29994_, _29992_);
  and _80359_ (_29996_, _29995_, _29968_);
  nor _80360_ (_29997_, _29996_, _10256_);
  nor _80361_ (_29999_, _29951_, _10255_);
  nor _80362_ (_30000_, _29999_, _29706_);
  not _80363_ (_30001_, _30000_);
  nor _80364_ (_30002_, _30001_, _29997_);
  nor _80365_ (_30003_, _10302_, _12901_);
  or _80366_ (_30004_, _30003_, _26212_);
  nor _80367_ (_30005_, _30004_, _30002_);
  nor _80368_ (_30006_, _30005_, _29961_);
  nor _80369_ (_30007_, _30006_, _03575_);
  and _80370_ (_30008_, _12901_, _03575_);
  nor _80371_ (_30010_, _30008_, _26220_);
  not _80372_ (_30011_, _30010_);
  nor _80373_ (_30012_, _30011_, _30007_);
  nor _80374_ (_30013_, _30012_, _29960_);
  nor _80375_ (_30014_, _30013_, _29716_);
  nor _80376_ (_30015_, _10251_, _12901_);
  nor _80377_ (_30016_, _30015_, _10326_);
  not _80378_ (_30017_, _30016_);
  nor _80379_ (_30018_, _30017_, _30014_);
  and _80380_ (_30019_, _10360_, _10138_);
  not _80381_ (_30021_, _29964_);
  nor _80382_ (_30022_, _30021_, _10360_);
  or _80383_ (_30023_, _30022_, _10325_);
  nor _80384_ (_30024_, _30023_, _30019_);
  nor _80385_ (_30025_, _30024_, _03657_);
  not _80386_ (_30026_, _30025_);
  nor _80387_ (_30027_, _30026_, _30018_);
  nor _80388_ (_30028_, _30021_, _10116_);
  and _80389_ (_30029_, _10138_, _10116_);
  nor _80390_ (_30030_, _30029_, _30028_);
  nor _80391_ (_30032_, _30030_, _10328_);
  nor _80392_ (_30033_, _30032_, _30027_);
  nor _80393_ (_30034_, _30033_, _29019_);
  and _80394_ (_30035_, _10398_, _10138_);
  and _80395_ (_30036_, _29964_, _10399_);
  or _80396_ (_30037_, _30036_, _30035_);
  and _80397_ (_30038_, _30037_, _03638_);
  and _80398_ (_30039_, _10382_, _10139_);
  nor _80399_ (_30040_, _29964_, _10382_);
  or _80400_ (_30041_, _30040_, _03998_);
  nor _80401_ (_30043_, _30041_, _30039_);
  nor _80402_ (_30044_, _30043_, _30038_);
  and _80403_ (_30045_, _29951_, _10083_);
  not _80404_ (_30046_, _30045_);
  and _80405_ (_30047_, _30046_, _10408_);
  and _80406_ (_30048_, _30047_, _30044_);
  not _80407_ (_30049_, _30048_);
  nor _80408_ (_30050_, _30049_, _30034_);
  nor _80409_ (_30051_, _30050_, _29959_);
  nor _80410_ (_30052_, _30051_, _25991_);
  nor _80411_ (_30054_, _29951_, _10415_);
  nor _80412_ (_30055_, _30054_, _10423_);
  not _80413_ (_30056_, _30055_);
  or _80414_ (_30057_, _30056_, _30052_);
  nor _80415_ (_30058_, _10422_, _12901_);
  nor _80416_ (_30059_, _30058_, _26302_);
  nand _80417_ (_30060_, _30059_, _30057_);
  nor _80418_ (_30061_, _29951_, _10426_);
  nor _80419_ (_30062_, _30061_, _10431_);
  nand _80420_ (_30063_, _30062_, _30060_);
  nor _80421_ (_30065_, _12901_, _10430_);
  nor _80422_ (_30066_, _30065_, _03311_);
  nand _80423_ (_30067_, _30066_, _30063_);
  not _80424_ (_30068_, _10439_);
  nor _80425_ (_30069_, _29951_, _03254_);
  nor _80426_ (_30070_, _30069_, _30068_);
  nand _80427_ (_30071_, _30070_, _30067_);
  nor _80428_ (_30072_, _10439_, _12901_);
  nor _80429_ (_30073_, _30072_, _03632_);
  nand _80430_ (_30074_, _30073_, _30071_);
  and _80431_ (_30076_, _10139_, _03632_);
  nor _80432_ (_30077_, _30076_, _26322_);
  nand _80433_ (_30078_, _30077_, _30074_);
  nor _80434_ (_30079_, _12901_, _03493_);
  nor _80435_ (_30080_, _30079_, _03221_);
  nand _80436_ (_30081_, _30080_, _30078_);
  and _80437_ (_30082_, _10139_, _03221_);
  nor _80438_ (_30083_, _30082_, _26330_);
  nand _80439_ (_30084_, _30083_, _30081_);
  nor _80440_ (_30085_, _29952_, _10081_);
  nor _80441_ (_30086_, _30085_, _10454_);
  nand _80442_ (_30087_, _30086_, _30084_);
  nor _80443_ (_30088_, _10453_, _09981_);
  nor _80444_ (_30089_, _30088_, _10458_);
  and _80445_ (_30090_, _30089_, _30087_);
  and _80446_ (_30091_, _29971_, _10458_);
  nor _80447_ (_30092_, _30091_, _30090_);
  or _80448_ (_30093_, _30092_, _06055_);
  or _80449_ (_30094_, _12901_, _05775_);
  and _80450_ (_30095_, _30094_, _03438_);
  nand _80451_ (_30098_, _30095_, _30093_);
  and _80452_ (_30099_, _10139_, _03437_);
  nor _80453_ (_30100_, _30099_, _08385_);
  nand _80454_ (_30101_, _30100_, _30098_);
  and _80455_ (_30102_, _09981_, _08385_);
  nor _80456_ (_30103_, _30102_, _10472_);
  nand _80457_ (_30104_, _30103_, _30101_);
  nor _80458_ (_30105_, _10503_, \oc8051_golden_model_1.DPH [4]);
  nor _80459_ (_30106_, _30105_, _10504_);
  nor _80460_ (_30107_, _30106_, _25897_);
  nor _80461_ (_30109_, _30107_, _10512_);
  and _80462_ (_30110_, _30109_, _30104_);
  or _80463_ (_30111_, _30110_, _29958_);
  nand _80464_ (_30112_, _30111_, _10515_);
  and _80465_ (_30113_, _09981_, _08698_);
  and _80466_ (_30114_, _29971_, _10077_);
  or _80467_ (_30115_, _30114_, _30113_);
  and _80468_ (_30116_, _30115_, _10076_);
  nor _80469_ (_30117_, _30116_, _26754_);
  nand _80470_ (_30118_, _30117_, _30112_);
  nor _80471_ (_30120_, _29951_, _10520_);
  nor _80472_ (_30121_, _30120_, _10524_);
  nand _80473_ (_30122_, _30121_, _30118_);
  nor _80474_ (_30123_, _10523_, _12901_);
  nor _80475_ (_30124_, _30123_, _03636_);
  nand _80476_ (_30125_, _30124_, _30122_);
  not _80477_ (_30126_, _10531_);
  and _80478_ (_30127_, _10139_, _03636_);
  nor _80479_ (_30128_, _30127_, _30126_);
  and _80480_ (_30129_, _30128_, _30125_);
  or _80481_ (_30131_, _30129_, _29957_);
  nand _80482_ (_30132_, _30131_, _10535_);
  nor _80483_ (_30133_, _29971_, _10077_);
  nor _80484_ (_30134_, _09981_, _08698_);
  nor _80485_ (_30135_, _30134_, _10535_);
  not _80486_ (_30136_, _30135_);
  nor _80487_ (_30137_, _30136_, _30133_);
  nor _80488_ (_30138_, _30137_, _10545_);
  nand _80489_ (_30139_, _30138_, _30132_);
  and _80490_ (_30140_, _29952_, _10545_);
  nor _80491_ (_30142_, _30140_, _10549_);
  nand _80492_ (_30143_, _30142_, _30139_);
  nor _80493_ (_30144_, _12901_, _10548_);
  nor _80494_ (_30145_, _30144_, _04504_);
  nand _80495_ (_30146_, _30145_, _30143_);
  not _80496_ (_30147_, _09960_);
  and _80497_ (_30148_, _10139_, _04504_);
  nor _80498_ (_30149_, _30148_, _30147_);
  and _80499_ (_30150_, _30149_, _30146_);
  or _80500_ (_30151_, _30150_, _29956_);
  nand _80501_ (_30153_, _30151_, _09959_);
  and _80502_ (_30154_, _09981_, \oc8051_golden_model_1.PSW [7]);
  and _80503_ (_30155_, _29971_, _07888_);
  or _80504_ (_30156_, _30155_, _30154_);
  and _80505_ (_30157_, _30156_, _09958_);
  nor _80506_ (_30158_, _30157_, _10560_);
  nand _80507_ (_30159_, _30158_, _30153_);
  nor _80508_ (_30160_, _29951_, _09956_);
  nor _80509_ (_30161_, _30160_, _08479_);
  nand _80510_ (_30162_, _30161_, _30159_);
  nor _80511_ (_30164_, _12901_, _08478_);
  nor _80512_ (_30165_, _30164_, _03758_);
  nand _80513_ (_30166_, _30165_, _30162_);
  not _80514_ (_30167_, _10573_);
  and _80515_ (_30168_, _10139_, _03758_);
  nor _80516_ (_30169_, _30168_, _30167_);
  and _80517_ (_30170_, _30169_, _30166_);
  or _80518_ (_30171_, _30170_, _29955_);
  nand _80519_ (_30172_, _30171_, _10577_);
  nor _80520_ (_30173_, _29971_, _07888_);
  nor _80521_ (_30175_, _09981_, \oc8051_golden_model_1.PSW [7]);
  nor _80522_ (_30176_, _30175_, _10577_);
  not _80523_ (_30177_, _30176_);
  nor _80524_ (_30178_, _30177_, _30173_);
  nor _80525_ (_30179_, _30178_, _10581_);
  nand _80526_ (_30180_, _30179_, _30172_);
  nor _80527_ (_30181_, _29951_, _09951_);
  nor _80528_ (_30182_, _30181_, _08525_);
  nand _80529_ (_30183_, _30182_, _30180_);
  nor _80530_ (_30184_, _12901_, _08524_);
  nor _80531_ (_30186_, _30184_, _08555_);
  nand _80532_ (_30187_, _30186_, _30183_);
  and _80533_ (_30188_, _29952_, _08555_);
  nor _80534_ (_30189_, _30188_, _03775_);
  and _80535_ (_30190_, _30189_, _30187_);
  nor _80536_ (_30191_, _05712_, _11403_);
  or _80537_ (_30192_, _30191_, _03179_);
  or _80538_ (_30193_, _30192_, _30190_);
  and _80539_ (_30194_, _12901_, _03179_);
  nor _80540_ (_30195_, _30194_, _03627_);
  nand _80541_ (_30197_, _30195_, _30193_);
  and _80542_ (_30198_, _30021_, _10794_);
  nor _80543_ (_30199_, _10794_, _10138_);
  or _80544_ (_30200_, _30199_, _10599_);
  or _80545_ (_30201_, _30200_, _30198_);
  and _80546_ (_30202_, _30201_, _09949_);
  nand _80547_ (_30203_, _30202_, _30197_);
  nor _80548_ (_30204_, _29951_, _09949_);
  nor _80549_ (_30205_, _30204_, _09937_);
  nand _80550_ (_30206_, _30205_, _30203_);
  nor _80551_ (_30208_, _12901_, _09936_);
  nor _80552_ (_30209_, _30208_, _07729_);
  and _80553_ (_30210_, _30209_, _30206_);
  or _80554_ (_30211_, _30210_, _29953_);
  nand _80555_ (_30212_, _30211_, _03523_);
  and _80556_ (_30213_, _05712_, _03522_);
  nor _80557_ (_30214_, _30213_, _03172_);
  and _80558_ (_30215_, _30214_, _30212_);
  and _80559_ (_30216_, _09981_, _03172_);
  or _80560_ (_30217_, _30216_, _03628_);
  nor _80561_ (_30219_, _30217_, _30215_);
  nor _80562_ (_30220_, _29964_, _10794_);
  and _80563_ (_30221_, _10794_, _10139_);
  nor _80564_ (_30222_, _30221_, _30220_);
  nor _80565_ (_30223_, _30222_, _03791_);
  or _80566_ (_30224_, _30223_, _30219_);
  and _80567_ (_30225_, _30224_, _10821_);
  nor _80568_ (_30226_, _29951_, _10821_);
  or _80569_ (_30227_, _30226_, _30225_);
  nand _80570_ (_30228_, _30227_, _04192_);
  and _80571_ (_30230_, _12901_, _03790_);
  nor _80572_ (_30231_, _30230_, _27228_);
  nand _80573_ (_30232_, _30231_, _30228_);
  nor _80574_ (_30233_, _29952_, _10828_);
  nor _80575_ (_30234_, _30233_, _03641_);
  nand _80576_ (_30235_, _30234_, _30232_);
  and _80577_ (_30236_, _04249_, _03641_);
  nor _80578_ (_30237_, _30236_, _03160_);
  and _80579_ (_30238_, _30237_, _30235_);
  and _80580_ (_30239_, _09981_, _03160_);
  or _80581_ (_30241_, _30239_, _03151_);
  or _80582_ (_30242_, _30241_, _30238_);
  nor _80583_ (_30243_, _30222_, _03152_);
  nor _80584_ (_30244_, _30243_, _10845_);
  nand _80585_ (_30245_, _30244_, _30242_);
  nor _80586_ (_30246_, _29952_, _10844_);
  nor _80587_ (_30247_, _30246_, _03520_);
  nand _80588_ (_30248_, _30247_, _30245_);
  and _80589_ (_30249_, _12901_, _03520_);
  nor _80590_ (_30250_, _30249_, _28299_);
  nand _80591_ (_30252_, _30250_, _30248_);
  nor _80592_ (_30253_, _29952_, _10851_);
  nor _80593_ (_30254_, _30253_, _03645_);
  nand _80594_ (_30255_, _30254_, _30252_);
  and _80595_ (_30256_, _04249_, _03645_);
  nor _80596_ (_30257_, _30256_, _03166_);
  nand _80597_ (_30258_, _30257_, _30255_);
  and _80598_ (_30259_, _09981_, _03166_);
  nor _80599_ (_30260_, _30259_, _10862_);
  and _80600_ (_30261_, _30260_, _30258_);
  and _80601_ (_30263_, _29952_, _10862_);
  nor _80602_ (_30264_, _30263_, _30261_);
  or _80603_ (_30265_, _30264_, _42967_);
  or _80604_ (_30266_, _42963_, \oc8051_golden_model_1.PC [12]);
  and _80605_ (_30267_, _30266_, _41755_);
  and _80606_ (_43341_, _30267_, _30265_);
  and _80607_ (_30268_, _29949_, \oc8051_golden_model_1.PC [13]);
  nor _80608_ (_30269_, _29949_, \oc8051_golden_model_1.PC [13]);
  nor _80609_ (_30270_, _30269_, _30268_);
  or _80610_ (_30271_, _30270_, _09949_);
  or _80611_ (_30273_, _30270_, _09951_);
  or _80612_ (_30274_, _10573_, _09977_);
  and _80613_ (_30275_, _30274_, _10577_);
  or _80614_ (_30276_, _30270_, _09956_);
  or _80615_ (_30277_, _09977_, _09960_);
  and _80616_ (_30278_, _30277_, _09959_);
  or _80617_ (_30279_, _09979_, _09978_);
  not _80618_ (_30280_, _30279_);
  nor _80619_ (_30281_, _30280_, _10064_);
  and _80620_ (_30282_, _30280_, _10064_);
  or _80621_ (_30284_, _30282_, _30281_);
  or _80622_ (_30285_, _30284_, _08698_);
  or _80623_ (_30286_, _09977_, _10077_);
  and _80624_ (_30287_, _30286_, _10076_);
  and _80625_ (_30288_, _30287_, _30285_);
  or _80626_ (_30289_, _09977_, _05775_);
  and _80627_ (_30290_, _10133_, _03221_);
  or _80628_ (_30291_, _30270_, _10426_);
  or _80629_ (_30292_, _10422_, _09977_);
  and _80630_ (_30293_, _10133_, _10116_);
  or _80631_ (_30295_, _10136_, _10135_);
  not _80632_ (_30296_, _30295_);
  nor _80633_ (_30297_, _30296_, _10234_);
  and _80634_ (_30298_, _30296_, _10234_);
  nor _80635_ (_30299_, _30298_, _30297_);
  nor _80636_ (_30300_, _30299_, _10116_);
  or _80637_ (_30301_, _30300_, _11574_);
  or _80638_ (_30302_, _30301_, _30293_);
  nand _80639_ (_30303_, _10360_, _10134_);
  not _80640_ (_30304_, _30299_);
  or _80641_ (_30306_, _30304_, _10360_);
  and _80642_ (_30307_, _30306_, _10326_);
  and _80643_ (_30308_, _30307_, _30303_);
  and _80644_ (_30309_, _09977_, _03575_);
  or _80645_ (_30310_, _10302_, _09977_);
  nand _80646_ (_30311_, _10261_, _10134_);
  or _80647_ (_30312_, _30304_, _10261_);
  and _80648_ (_30313_, _30312_, _03570_);
  and _80649_ (_30314_, _30313_, _30311_);
  and _80650_ (_30315_, _10269_, _09977_);
  and _80651_ (_30317_, _30284_, _10271_);
  or _80652_ (_30318_, _30317_, _05831_);
  or _80653_ (_30319_, _30318_, _30315_);
  or _80654_ (_30320_, _09977_, _26179_);
  or _80655_ (_30321_, _03923_, \oc8051_golden_model_1.PC [13]);
  nor _80656_ (_30322_, _30321_, _04426_);
  nand _80657_ (_30323_, _30322_, _10278_);
  and _80658_ (_30324_, _30323_, _30320_);
  or _80659_ (_30325_, _30324_, _26577_);
  or _80660_ (_30326_, _09977_, _04762_);
  and _80661_ (_30328_, _30326_, _30325_);
  or _80662_ (_30329_, _30328_, _27661_);
  or _80663_ (_30330_, _30270_, _29382_);
  and _80664_ (_30331_, _30330_, _30329_);
  or _80665_ (_30332_, _30331_, _05833_);
  and _80666_ (_30333_, _30332_, _10296_);
  and _80667_ (_30334_, _30333_, _30319_);
  or _80668_ (_30335_, _30334_, _30314_);
  and _80669_ (_30336_, _30335_, _10255_);
  not _80670_ (_30337_, _30270_);
  nor _80671_ (_30339_, _30337_, _10303_);
  or _80672_ (_30340_, _30339_, _29706_);
  or _80673_ (_30341_, _30340_, _30336_);
  and _80674_ (_30342_, _30341_, _30310_);
  or _80675_ (_30343_, _30342_, _26212_);
  or _80676_ (_30344_, _30270_, _10307_);
  and _80677_ (_30345_, _30344_, _03583_);
  and _80678_ (_30346_, _30345_, _30343_);
  or _80679_ (_30347_, _30346_, _30309_);
  and _80680_ (_30348_, _30347_, _10316_);
  or _80681_ (_30350_, _30337_, _10316_);
  nand _80682_ (_30351_, _30350_, _10251_);
  or _80683_ (_30352_, _30351_, _30348_);
  or _80684_ (_30353_, _10251_, _09977_);
  and _80685_ (_30354_, _30353_, _10325_);
  and _80686_ (_30355_, _30354_, _30352_);
  or _80687_ (_30356_, _30355_, _30308_);
  or _80688_ (_30357_, _30356_, _27272_);
  and _80689_ (_30358_, _30357_, _30302_);
  and _80690_ (_30359_, _30358_, _11596_);
  nand _80691_ (_30361_, _30299_, _10399_);
  nand _80692_ (_30362_, _10398_, _10134_);
  and _80693_ (_30363_, _30362_, _03638_);
  and _80694_ (_30364_, _30363_, _30361_);
  and _80695_ (_30365_, _10382_, _10133_);
  nor _80696_ (_30366_, _30299_, _10382_);
  or _80697_ (_30367_, _30366_, _30365_);
  and _80698_ (_30368_, _30367_, _03527_);
  or _80699_ (_30369_, _30368_, _30364_);
  nand _80700_ (_30370_, _30270_, _10083_);
  nand _80701_ (_30372_, _30370_, _10408_);
  or _80702_ (_30373_, _30372_, _30369_);
  or _80703_ (_30374_, _30373_, _30359_);
  or _80704_ (_30375_, _10408_, _09977_);
  and _80705_ (_30376_, _30375_, _10415_);
  and _80706_ (_30377_, _30376_, _30374_);
  nor _80707_ (_30378_, _30337_, _10415_);
  or _80708_ (_30379_, _30378_, _10423_);
  or _80709_ (_30380_, _30379_, _30377_);
  and _80710_ (_30381_, _30380_, _30292_);
  or _80711_ (_30383_, _30381_, _26302_);
  and _80712_ (_30384_, _30383_, _30291_);
  or _80713_ (_30385_, _30384_, _10431_);
  or _80714_ (_30386_, _09977_, _10430_);
  and _80715_ (_30387_, _30386_, _03254_);
  and _80716_ (_30388_, _30387_, _30385_);
  nand _80717_ (_30389_, _30270_, _03311_);
  nand _80718_ (_30390_, _30389_, _10439_);
  or _80719_ (_30391_, _30390_, _30388_);
  or _80720_ (_30392_, _10439_, _09977_);
  and _80721_ (_30394_, _30392_, _09755_);
  and _80722_ (_30395_, _30394_, _30391_);
  nand _80723_ (_30396_, _10133_, _03632_);
  nand _80724_ (_30397_, _30396_, _03493_);
  or _80725_ (_30398_, _30397_, _30395_);
  or _80726_ (_30399_, _09977_, _03493_);
  and _80727_ (_30400_, _30399_, _03474_);
  and _80728_ (_30401_, _30400_, _30398_);
  or _80729_ (_30402_, _30401_, _30290_);
  and _80730_ (_30403_, _30402_, _10081_);
  nor _80731_ (_30405_, _30337_, _10081_);
  or _80732_ (_30406_, _30405_, _10454_);
  or _80733_ (_30407_, _30406_, _30403_);
  or _80734_ (_30408_, _10453_, _09977_);
  and _80735_ (_30409_, _30408_, _10459_);
  and _80736_ (_30410_, _30409_, _30407_);
  and _80737_ (_30411_, _30284_, _10458_);
  or _80738_ (_30412_, _30411_, _06055_);
  or _80739_ (_30413_, _30412_, _30410_);
  and _80740_ (_30414_, _30413_, _30289_);
  or _80741_ (_30415_, _30414_, _03437_);
  or _80742_ (_30416_, _10133_, _03438_);
  and _80743_ (_30417_, _30416_, _08386_);
  and _80744_ (_30418_, _30417_, _30415_);
  and _80745_ (_30419_, _09977_, _08385_);
  or _80746_ (_30420_, _30419_, _30418_);
  and _80747_ (_30421_, _30420_, _25897_);
  or _80748_ (_30422_, _10504_, \oc8051_golden_model_1.DPH [5]);
  nor _80749_ (_30423_, _10505_, _25897_);
  and _80750_ (_30424_, _30423_, _30422_);
  or _80751_ (_30427_, _30424_, _10512_);
  or _80752_ (_30428_, _30427_, _30421_);
  or _80753_ (_30429_, _10511_, _09977_);
  and _80754_ (_30430_, _30429_, _10515_);
  and _80755_ (_30431_, _30430_, _30428_);
  or _80756_ (_30432_, _30431_, _30288_);
  and _80757_ (_30433_, _30432_, _10520_);
  nor _80758_ (_30434_, _30337_, _10520_);
  or _80759_ (_30435_, _30434_, _10524_);
  or _80760_ (_30436_, _30435_, _30433_);
  or _80761_ (_30438_, _10523_, _09977_);
  and _80762_ (_30439_, _30438_, _04499_);
  and _80763_ (_30440_, _30439_, _30436_);
  nand _80764_ (_30441_, _10133_, _03636_);
  nand _80765_ (_30442_, _30441_, _10531_);
  or _80766_ (_30443_, _30442_, _30440_);
  or _80767_ (_30444_, _10531_, _09977_);
  and _80768_ (_30445_, _30444_, _10535_);
  and _80769_ (_30446_, _30445_, _30443_);
  or _80770_ (_30447_, _30284_, _10077_);
  or _80771_ (_30449_, _09977_, _08698_);
  and _80772_ (_30450_, _30449_, _10534_);
  and _80773_ (_30451_, _30450_, _30447_);
  or _80774_ (_30452_, _30451_, _30446_);
  and _80775_ (_30453_, _30452_, _10546_);
  and _80776_ (_30454_, _30270_, _10545_);
  or _80777_ (_30455_, _30454_, _10549_);
  or _80778_ (_30456_, _30455_, _30453_);
  or _80779_ (_30457_, _09977_, _10548_);
  and _80780_ (_30458_, _30457_, _05769_);
  and _80781_ (_30460_, _30458_, _30456_);
  nand _80782_ (_30461_, _10133_, _03754_);
  nand _80783_ (_30462_, _30461_, _09960_);
  or _80784_ (_30463_, _30462_, _30460_);
  and _80785_ (_30464_, _30463_, _30278_);
  or _80786_ (_30465_, _30284_, \oc8051_golden_model_1.PSW [7]);
  or _80787_ (_30466_, _09977_, _07888_);
  and _80788_ (_30467_, _30466_, _09958_);
  and _80789_ (_30468_, _30467_, _30465_);
  or _80790_ (_30469_, _30468_, _10560_);
  or _80791_ (_30471_, _30469_, _30464_);
  and _80792_ (_30472_, _30471_, _30276_);
  or _80793_ (_30473_, _30472_, _08479_);
  or _80794_ (_30474_, _09977_, _08478_);
  and _80795_ (_30475_, _30474_, _03759_);
  and _80796_ (_30476_, _30475_, _30473_);
  nand _80797_ (_30477_, _10133_, _03758_);
  nand _80798_ (_30478_, _30477_, _10573_);
  or _80799_ (_30479_, _30478_, _30476_);
  and _80800_ (_30480_, _30479_, _30275_);
  or _80801_ (_30482_, _30284_, _07888_);
  or _80802_ (_30483_, _09977_, \oc8051_golden_model_1.PSW [7]);
  and _80803_ (_30484_, _30483_, _10576_);
  and _80804_ (_30485_, _30484_, _30482_);
  or _80805_ (_30486_, _30485_, _10581_);
  or _80806_ (_30487_, _30486_, _30480_);
  and _80807_ (_30488_, _30487_, _30273_);
  or _80808_ (_30489_, _30488_, _08525_);
  or _80809_ (_30490_, _09977_, _08524_);
  and _80810_ (_30492_, _30490_, _08556_);
  and _80811_ (_30495_, _30492_, _30489_);
  and _80812_ (_30497_, _30270_, _08555_);
  or _80813_ (_30499_, _30497_, _03775_);
  or _80814_ (_30501_, _30499_, _30495_);
  nand _80815_ (_30503_, _05422_, _03775_);
  and _80816_ (_30505_, _30503_, _30501_);
  or _80817_ (_30507_, _30505_, _03179_);
  or _80818_ (_30509_, _09977_, _06328_);
  and _80819_ (_30511_, _30509_, _10599_);
  and _80820_ (_30513_, _30511_, _30507_);
  nand _80821_ (_30515_, _30299_, _10794_);
  or _80822_ (_30516_, _10794_, _10133_);
  and _80823_ (_30517_, _30516_, _03627_);
  and _80824_ (_30518_, _30517_, _30515_);
  or _80825_ (_30519_, _30518_, _10603_);
  or _80826_ (_30520_, _30519_, _30513_);
  and _80827_ (_30521_, _30520_, _30271_);
  or _80828_ (_30522_, _30521_, _09937_);
  or _80829_ (_30523_, _09977_, _09936_);
  and _80830_ (_30524_, _30523_, _10803_);
  and _80831_ (_30526_, _30524_, _30522_);
  and _80832_ (_30527_, _30270_, _07729_);
  or _80833_ (_30528_, _30527_, _03522_);
  or _80834_ (_30529_, _30528_, _30526_);
  nand _80835_ (_30530_, _05422_, _03522_);
  and _80836_ (_30531_, _30530_, _30529_);
  or _80837_ (_30532_, _30531_, _03172_);
  or _80838_ (_30533_, _09977_, _25887_);
  and _80839_ (_30534_, _30533_, _03791_);
  and _80840_ (_30535_, _30534_, _30532_);
  nand _80841_ (_30537_, _10794_, _10134_);
  or _80842_ (_30538_, _30304_, _10794_);
  and _80843_ (_30539_, _30538_, _30537_);
  and _80844_ (_30540_, _30539_, _03628_);
  or _80845_ (_30541_, _30540_, _10822_);
  or _80846_ (_30542_, _30541_, _30535_);
  or _80847_ (_30543_, _30270_, _10821_);
  and _80848_ (_30544_, _30543_, _04192_);
  and _80849_ (_30545_, _30544_, _30542_);
  nand _80850_ (_30546_, _09977_, _03790_);
  nand _80851_ (_30548_, _30546_, _10828_);
  or _80852_ (_30549_, _30548_, _30545_);
  or _80853_ (_30550_, _30270_, _10828_);
  and _80854_ (_30551_, _30550_, _10832_);
  and _80855_ (_30552_, _30551_, _30549_);
  nor _80856_ (_30553_, _03834_, _10832_);
  or _80857_ (_30554_, _30553_, _03160_);
  or _80858_ (_30555_, _30554_, _30552_);
  or _80859_ (_30556_, _09977_, _03161_);
  and _80860_ (_30557_, _30556_, _03152_);
  and _80861_ (_30559_, _30557_, _30555_);
  and _80862_ (_30560_, _30539_, _03151_);
  or _80863_ (_30561_, _30560_, _10845_);
  or _80864_ (_30562_, _30561_, _30559_);
  or _80865_ (_30563_, _30270_, _10844_);
  and _80866_ (_30564_, _30563_, _03521_);
  and _80867_ (_30565_, _30564_, _30562_);
  nand _80868_ (_30566_, _09977_, _03520_);
  nand _80869_ (_30567_, _30566_, _10851_);
  or _80870_ (_30568_, _30567_, _30565_);
  or _80871_ (_30570_, _30270_, _10851_);
  and _80872_ (_30571_, _30570_, _10855_);
  and _80873_ (_30572_, _30571_, _30568_);
  nand _80874_ (_30573_, _03834_, _29936_);
  and _80875_ (_30574_, _30573_, _25883_);
  or _80876_ (_30575_, _30574_, _30572_);
  or _80877_ (_30576_, _09977_, _29936_);
  and _80878_ (_30577_, _30576_, _10863_);
  and _80879_ (_30578_, _30577_, _30575_);
  and _80880_ (_30579_, _30270_, _10862_);
  or _80881_ (_30581_, _30579_, _30578_);
  or _80882_ (_30582_, _30581_, _42967_);
  or _80883_ (_30583_, _42963_, \oc8051_golden_model_1.PC [13]);
  and _80884_ (_30584_, _30583_, _41755_);
  and _80885_ (_43342_, _30584_, _30582_);
  and _80886_ (_30585_, _03645_, _03561_);
  and _80887_ (_30586_, _30268_, \oc8051_golden_model_1.PC [14]);
  nor _80888_ (_30587_, _30268_, \oc8051_golden_model_1.PC [14]);
  nor _80889_ (_30588_, _30587_, _30586_);
  nor _80890_ (_30589_, _30588_, _10803_);
  not _80891_ (_30591_, _09971_);
  nor _80892_ (_30592_, _10573_, _30591_);
  nor _80893_ (_30593_, _30591_, _09960_);
  nor _80894_ (_30594_, _10531_, _30591_);
  nor _80895_ (_30595_, _10511_, _30591_);
  nor _80896_ (_30596_, _10408_, _09971_);
  or _80897_ (_30597_, _30588_, _10307_);
  and _80898_ (_30598_, _30588_, _04438_);
  and _80899_ (_30599_, _10269_, _09971_);
  and _80900_ (_30600_, _10066_, _09975_);
  nor _80901_ (_30602_, _30600_, _10067_);
  and _80902_ (_30603_, _30602_, _10271_);
  or _80903_ (_30604_, _30603_, _30599_);
  or _80904_ (_30605_, _30604_, _05831_);
  or _80905_ (_30606_, _09971_, _04762_);
  and _80906_ (_30607_, _30606_, _10290_);
  or _80907_ (_30608_, _09971_, _26179_);
  nor _80908_ (_30609_, _04426_, \oc8051_golden_model_1.PC [14]);
  nand _80909_ (_30610_, _30609_, _10278_);
  and _80910_ (_30611_, _30610_, _30608_);
  or _80911_ (_30613_, _30611_, _26577_);
  or _80912_ (_30614_, _30588_, _25905_);
  and _80913_ (_30615_, _30614_, _30613_);
  or _80914_ (_30616_, _30615_, _03923_);
  and _80915_ (_30617_, _30616_, _30607_);
  not _80916_ (_30618_, _30588_);
  nor _80917_ (_30619_, _30618_, _10290_);
  or _80918_ (_30620_, _30619_, _05833_);
  or _80919_ (_30621_, _30620_, _30617_);
  and _80920_ (_30622_, _30621_, _05847_);
  and _80921_ (_30624_, _30622_, _30605_);
  or _80922_ (_30625_, _30624_, _30598_);
  and _80923_ (_30626_, _30625_, _04444_);
  nand _80924_ (_30627_, _10261_, _10127_);
  and _80925_ (_30628_, _10236_, _10131_);
  nor _80926_ (_30629_, _30628_, _10237_);
  or _80927_ (_30630_, _30629_, _10261_);
  and _80928_ (_30631_, _30630_, _30627_);
  and _80929_ (_30632_, _30631_, _03570_);
  or _80930_ (_30633_, _30632_, _30626_);
  or _80931_ (_30635_, _30633_, _10256_);
  or _80932_ (_30636_, _30588_, _10255_);
  and _80933_ (_30637_, _30636_, _10302_);
  and _80934_ (_30638_, _30637_, _30635_);
  or _80935_ (_30639_, _10302_, _30591_);
  nand _80936_ (_30640_, _30639_, _10307_);
  or _80937_ (_30641_, _30640_, _30638_);
  and _80938_ (_30642_, _30641_, _30597_);
  or _80939_ (_30643_, _30642_, _03575_);
  or _80940_ (_30644_, _09971_, _03583_);
  and _80941_ (_30646_, _30644_, _10316_);
  and _80942_ (_30647_, _30646_, _30643_);
  and _80943_ (_30648_, _30588_, _26220_);
  or _80944_ (_30649_, _30648_, _30647_);
  and _80945_ (_30650_, _30649_, _10251_);
  or _80946_ (_30651_, _10251_, _30591_);
  nand _80947_ (_30652_, _30651_, _10325_);
  or _80948_ (_30653_, _30652_, _30650_);
  and _80949_ (_30654_, _10360_, _10126_);
  not _80950_ (_30655_, _30629_);
  nor _80951_ (_30657_, _30655_, _10360_);
  or _80952_ (_30658_, _30657_, _30654_);
  or _80953_ (_30659_, _30658_, _10325_);
  and _80954_ (_30660_, _30659_, _30653_);
  or _80955_ (_30661_, _30660_, _27272_);
  nor _80956_ (_30662_, _30655_, _10116_);
  and _80957_ (_30663_, _10126_, _10116_);
  or _80958_ (_30664_, _30663_, _10328_);
  or _80959_ (_30665_, _30664_, _30662_);
  and _80960_ (_30666_, _30665_, _11596_);
  and _80961_ (_30668_, _30666_, _30661_);
  not _80962_ (_30669_, _30668_);
  and _80963_ (_30670_, _30588_, _10083_);
  not _80964_ (_30671_, _30670_);
  and _80965_ (_30672_, _30671_, _10408_);
  nor _80966_ (_30673_, _30629_, _10398_);
  and _80967_ (_30674_, _10398_, _10127_);
  nor _80968_ (_30675_, _30674_, _10085_);
  not _80969_ (_30676_, _30675_);
  nor _80970_ (_30677_, _30676_, _30673_);
  and _80971_ (_30678_, _10382_, _10127_);
  nor _80972_ (_30679_, _30629_, _10382_);
  or _80973_ (_30680_, _30679_, _03998_);
  nor _80974_ (_30681_, _30680_, _30678_);
  nor _80975_ (_30682_, _30681_, _30677_);
  and _80976_ (_30683_, _30682_, _30672_);
  and _80977_ (_30684_, _30683_, _30669_);
  nor _80978_ (_30685_, _30684_, _30596_);
  nor _80979_ (_30686_, _30685_, _25991_);
  nor _80980_ (_30687_, _30588_, _10415_);
  nor _80981_ (_30689_, _30687_, _10423_);
  not _80982_ (_30690_, _30689_);
  or _80983_ (_30691_, _30690_, _30686_);
  nor _80984_ (_30692_, _10422_, _30591_);
  nor _80985_ (_30693_, _30692_, _26302_);
  nand _80986_ (_30694_, _30693_, _30691_);
  nor _80987_ (_30695_, _30588_, _10426_);
  nor _80988_ (_30696_, _30695_, _10431_);
  and _80989_ (_30697_, _30696_, _30694_);
  nor _80990_ (_30698_, _30591_, _10430_);
  or _80991_ (_30700_, _30698_, _03311_);
  or _80992_ (_30701_, _30700_, _30697_);
  nor _80993_ (_30702_, _30588_, _03254_);
  nor _80994_ (_30703_, _30702_, _30068_);
  nand _80995_ (_30704_, _30703_, _30701_);
  nor _80996_ (_30705_, _10439_, _30591_);
  nor _80997_ (_30706_, _30705_, _03632_);
  and _80998_ (_30707_, _30706_, _30704_);
  nor _80999_ (_30708_, _10126_, _09755_);
  or _81000_ (_30709_, _30708_, _30707_);
  and _81001_ (_30711_, _30709_, _03493_);
  nor _81002_ (_30712_, _09971_, _03493_);
  or _81003_ (_30713_, _30712_, _30711_);
  nand _81004_ (_30714_, _30713_, _03474_);
  nor _81005_ (_30715_, _10126_, _03474_);
  nor _81006_ (_30716_, _30715_, _26330_);
  nand _81007_ (_30717_, _30716_, _30714_);
  nor _81008_ (_30718_, _30618_, _10081_);
  nor _81009_ (_30719_, _30718_, _10454_);
  nand _81010_ (_30720_, _30719_, _30717_);
  nor _81011_ (_30722_, _10453_, _09971_);
  nor _81012_ (_30723_, _30722_, _10458_);
  and _81013_ (_30724_, _30723_, _30720_);
  and _81014_ (_30725_, _30602_, _10458_);
  nor _81015_ (_30726_, _30725_, _30724_);
  or _81016_ (_30727_, _30726_, _06055_);
  or _81017_ (_30728_, _30591_, _05775_);
  and _81018_ (_30729_, _30728_, _03438_);
  nand _81019_ (_30730_, _30729_, _30727_);
  nor _81020_ (_30731_, _10126_, _03438_);
  nor _81021_ (_30733_, _30731_, _08385_);
  nand _81022_ (_30734_, _30733_, _30730_);
  and _81023_ (_30735_, _09971_, _08385_);
  nor _81024_ (_30736_, _30735_, _10472_);
  nand _81025_ (_30737_, _30736_, _30734_);
  nor _81026_ (_30738_, _10505_, \oc8051_golden_model_1.DPH [6]);
  nor _81027_ (_30739_, _30738_, _10506_);
  nor _81028_ (_30740_, _30739_, _25897_);
  nor _81029_ (_30741_, _30740_, _10512_);
  and _81030_ (_30742_, _30741_, _30737_);
  or _81031_ (_30744_, _30742_, _30595_);
  nand _81032_ (_30745_, _30744_, _10515_);
  and _81033_ (_30746_, _09971_, _08698_);
  and _81034_ (_30747_, _30602_, _10077_);
  or _81035_ (_30748_, _30747_, _30746_);
  and _81036_ (_30749_, _30748_, _10076_);
  nor _81037_ (_30750_, _30749_, _26754_);
  nand _81038_ (_30751_, _30750_, _30745_);
  nor _81039_ (_30752_, _30588_, _10520_);
  nor _81040_ (_30753_, _30752_, _10524_);
  nand _81041_ (_30755_, _30753_, _30751_);
  nor _81042_ (_30756_, _10523_, _30591_);
  nor _81043_ (_30757_, _30756_, _03636_);
  nand _81044_ (_30758_, _30757_, _30755_);
  nor _81045_ (_30759_, _10126_, _04499_);
  nor _81046_ (_30760_, _30759_, _30126_);
  and _81047_ (_30761_, _30760_, _30758_);
  or _81048_ (_30762_, _30761_, _30594_);
  nand _81049_ (_30763_, _30762_, _10535_);
  nor _81050_ (_30764_, _30602_, _10077_);
  nor _81051_ (_30766_, _09971_, _08698_);
  nor _81052_ (_30767_, _30766_, _10535_);
  not _81053_ (_30768_, _30767_);
  nor _81054_ (_30769_, _30768_, _30764_);
  nor _81055_ (_30770_, _30769_, _10545_);
  nand _81056_ (_30771_, _30770_, _30763_);
  and _81057_ (_30772_, _30618_, _10545_);
  nor _81058_ (_30773_, _30772_, _10549_);
  nand _81059_ (_30774_, _30773_, _30771_);
  nor _81060_ (_30775_, _30591_, _10548_);
  nor _81061_ (_30777_, _30775_, _04504_);
  nand _81062_ (_30778_, _30777_, _30774_);
  and _81063_ (_30779_, _10127_, _04504_);
  nor _81064_ (_30780_, _30779_, _30147_);
  and _81065_ (_30781_, _30780_, _30778_);
  or _81066_ (_30782_, _30781_, _30593_);
  nand _81067_ (_30783_, _30782_, _09959_);
  and _81068_ (_30784_, _09971_, \oc8051_golden_model_1.PSW [7]);
  and _81069_ (_30785_, _30602_, _07888_);
  or _81070_ (_30786_, _30785_, _30784_);
  and _81071_ (_30788_, _30786_, _09958_);
  nor _81072_ (_30789_, _30788_, _10560_);
  nand _81073_ (_30790_, _30789_, _30783_);
  nor _81074_ (_30791_, _30588_, _09956_);
  nor _81075_ (_30792_, _30791_, _08479_);
  nand _81076_ (_30793_, _30792_, _30790_);
  nor _81077_ (_30794_, _30591_, _08478_);
  nor _81078_ (_30795_, _30794_, _03758_);
  nand _81079_ (_30796_, _30795_, _30793_);
  nor _81080_ (_30797_, _10126_, _03759_);
  nor _81081_ (_30799_, _30797_, _30167_);
  and _81082_ (_30800_, _30799_, _30796_);
  or _81083_ (_30801_, _30800_, _30592_);
  nand _81084_ (_30802_, _30801_, _10577_);
  nor _81085_ (_30803_, _30602_, _07888_);
  nor _81086_ (_30804_, _09971_, \oc8051_golden_model_1.PSW [7]);
  nor _81087_ (_30805_, _30804_, _10577_);
  not _81088_ (_30806_, _30805_);
  nor _81089_ (_30807_, _30806_, _30803_);
  nor _81090_ (_30808_, _30807_, _10581_);
  nand _81091_ (_30810_, _30808_, _30802_);
  nor _81092_ (_30811_, _30588_, _09951_);
  nor _81093_ (_30812_, _30811_, _08525_);
  nand _81094_ (_30813_, _30812_, _30810_);
  nor _81095_ (_30814_, _30591_, _08524_);
  nor _81096_ (_30815_, _30814_, _08555_);
  nand _81097_ (_30816_, _30815_, _30813_);
  nor _81098_ (_30817_, _30588_, _08556_);
  nor _81099_ (_30818_, _30817_, _03775_);
  and _81100_ (_30819_, _30818_, _30816_);
  nor _81101_ (_30821_, _05327_, _11403_);
  or _81102_ (_30822_, _30821_, _03179_);
  or _81103_ (_30823_, _30822_, _30819_);
  nor _81104_ (_30824_, _09971_, _06328_);
  nor _81105_ (_30825_, _30824_, _03627_);
  nand _81106_ (_30826_, _30825_, _30823_);
  nor _81107_ (_30827_, _10794_, _10126_);
  and _81108_ (_30828_, _30655_, _10794_);
  or _81109_ (_30829_, _30828_, _10599_);
  or _81110_ (_30830_, _30829_, _30827_);
  and _81111_ (_30832_, _30830_, _09949_);
  nand _81112_ (_30833_, _30832_, _30826_);
  nor _81113_ (_30834_, _30588_, _09949_);
  nor _81114_ (_30835_, _30834_, _09937_);
  nand _81115_ (_30836_, _30835_, _30833_);
  nor _81116_ (_30837_, _30591_, _09936_);
  nor _81117_ (_30838_, _30837_, _07729_);
  and _81118_ (_30839_, _30838_, _30836_);
  or _81119_ (_30840_, _30839_, _30589_);
  nand _81120_ (_30841_, _30840_, _03523_);
  and _81121_ (_30843_, _05327_, _03522_);
  nor _81122_ (_30844_, _30843_, _03172_);
  and _81123_ (_30845_, _30844_, _30841_);
  and _81124_ (_30846_, _09971_, _03172_);
  or _81125_ (_30847_, _30846_, _03628_);
  nor _81126_ (_30848_, _30847_, _30845_);
  and _81127_ (_30849_, _10794_, _10127_);
  nor _81128_ (_30850_, _30629_, _10794_);
  nor _81129_ (_30851_, _30850_, _30849_);
  nor _81130_ (_30852_, _30851_, _03791_);
  or _81131_ (_30854_, _30852_, _30848_);
  and _81132_ (_30855_, _30854_, _10821_);
  nor _81133_ (_30856_, _30588_, _10821_);
  or _81134_ (_30857_, _30856_, _30855_);
  nand _81135_ (_30858_, _30857_, _04192_);
  nor _81136_ (_30859_, _09971_, _04192_);
  nor _81137_ (_30860_, _30859_, _27228_);
  nand _81138_ (_30861_, _30860_, _30858_);
  nor _81139_ (_30862_, _30618_, _10828_);
  nor _81140_ (_30863_, _30862_, _03641_);
  nand _81141_ (_30865_, _30863_, _30861_);
  and _81142_ (_30866_, _03641_, _03561_);
  nor _81143_ (_30867_, _30866_, _03160_);
  and _81144_ (_30868_, _30867_, _30865_);
  and _81145_ (_30869_, _09971_, _03160_);
  or _81146_ (_30870_, _30869_, _03151_);
  or _81147_ (_30871_, _30870_, _30868_);
  nor _81148_ (_30872_, _30851_, _03152_);
  nor _81149_ (_30873_, _30872_, _10845_);
  nand _81150_ (_30874_, _30873_, _30871_);
  nor _81151_ (_30876_, _30618_, _10844_);
  nor _81152_ (_30877_, _30876_, _03520_);
  nand _81153_ (_30878_, _30877_, _30874_);
  nor _81154_ (_30879_, _09971_, _03521_);
  nor _81155_ (_30880_, _30879_, _28299_);
  nand _81156_ (_30881_, _30880_, _30878_);
  nor _81157_ (_30882_, _30618_, _10851_);
  nor _81158_ (_30883_, _30882_, _03645_);
  and _81159_ (_30884_, _30883_, _30881_);
  or _81160_ (_30885_, _30884_, _30585_);
  nand _81161_ (_30887_, _30885_, _29936_);
  nor _81162_ (_30888_, _09971_, _29936_);
  nor _81163_ (_30889_, _30888_, _10862_);
  and _81164_ (_30890_, _30889_, _30887_);
  and _81165_ (_30891_, _30588_, _10862_);
  or _81166_ (_30892_, _30891_, _30890_);
  or _81167_ (_30893_, _30892_, _42967_);
  or _81168_ (_30894_, _42963_, \oc8051_golden_model_1.PC [14]);
  and _81169_ (_30895_, _30894_, _41755_);
  and _81170_ (_43343_, _30895_, _30893_);
  nor _81171_ (_30897_, \oc8051_golden_model_1.P2 [0], rst);
  nor _81172_ (_30898_, _30897_, _00000_);
  and _81173_ (_30899_, _10872_, \oc8051_golden_model_1.P2 [0]);
  and _81174_ (_30900_, _11995_, _05210_);
  or _81175_ (_30901_, _30900_, _30899_);
  and _81176_ (_30902_, _30901_, _03769_);
  and _81177_ (_30903_, _05210_, _04419_);
  or _81178_ (_30904_, _30903_, _30899_);
  or _81179_ (_30905_, _30904_, _06039_);
  and _81180_ (_30906_, _05941_, _05210_);
  or _81181_ (_30907_, _30906_, _30899_);
  or _81182_ (_30908_, _30907_, _04444_);
  and _81183_ (_30909_, _05210_, \oc8051_golden_model_1.ACC [0]);
  or _81184_ (_30910_, _30909_, _30899_);
  and _81185_ (_30911_, _30910_, _04426_);
  and _81186_ (_30912_, _04427_, \oc8051_golden_model_1.P2 [0]);
  or _81187_ (_30913_, _30912_, _03570_);
  or _81188_ (_30914_, _30913_, _30911_);
  and _81189_ (_30915_, _30914_, _03517_);
  and _81190_ (_30916_, _30915_, _30908_);
  and _81191_ (_30919_, _10880_, \oc8051_golden_model_1.P2 [0]);
  and _81192_ (_30920_, _11887_, _05801_);
  or _81193_ (_30921_, _30920_, _30919_);
  and _81194_ (_30922_, _30921_, _03516_);
  or _81195_ (_30923_, _30922_, _30916_);
  and _81196_ (_30924_, _30923_, _03983_);
  and _81197_ (_30925_, _30904_, _03568_);
  or _81198_ (_30926_, _30925_, _03575_);
  or _81199_ (_30927_, _30926_, _30924_);
  or _81200_ (_30928_, _30910_, _03583_);
  and _81201_ (_30930_, _30928_, _03513_);
  and _81202_ (_30931_, _30930_, _30927_);
  and _81203_ (_30932_, _30899_, _03512_);
  or _81204_ (_30933_, _30932_, _03505_);
  or _81205_ (_30934_, _30933_, _30931_);
  or _81206_ (_30935_, _30907_, _03506_);
  and _81207_ (_30936_, _30935_, _03500_);
  and _81208_ (_30937_, _30936_, _30934_);
  or _81209_ (_30938_, _11915_, _11875_);
  and _81210_ (_30939_, _30938_, _05801_);
  or _81211_ (_30941_, _30939_, _30919_);
  and _81212_ (_30942_, _30941_, _03499_);
  or _81213_ (_30943_, _30942_, _07314_);
  or _81214_ (_30944_, _30943_, _30937_);
  and _81215_ (_30945_, _30944_, _30905_);
  or _81216_ (_30946_, _30945_, _03479_);
  and _81217_ (_30947_, _06715_, _05210_);
  or _81218_ (_30948_, _30899_, _06044_);
  or _81219_ (_30949_, _30948_, _30947_);
  and _81220_ (_30950_, _30949_, _03474_);
  and _81221_ (_30952_, _30950_, _30946_);
  and _81222_ (_30953_, _06245_, \oc8051_golden_model_1.P1 [0]);
  and _81223_ (_30954_, _06249_, \oc8051_golden_model_1.P3 [0]);
  or _81224_ (_30955_, _30954_, _30953_);
  or _81225_ (_30956_, _30955_, _11952_);
  and _81226_ (_30957_, _06242_, \oc8051_golden_model_1.P0 [0]);
  and _81227_ (_30958_, _06214_, \oc8051_golden_model_1.P2 [0]);
  or _81228_ (_30959_, _30958_, _30957_);
  nor _81229_ (_30960_, _30959_, _30956_);
  and _81230_ (_30961_, _30960_, _11970_);
  and _81231_ (_30963_, _30961_, _11951_);
  nand _81232_ (_30964_, _30963_, _11944_);
  or _81233_ (_30965_, _30964_, _11929_);
  and _81234_ (_30966_, _30965_, _05210_);
  or _81235_ (_30967_, _30966_, _30899_);
  and _81236_ (_30968_, _30967_, _03221_);
  or _81237_ (_30969_, _30968_, _03437_);
  or _81238_ (_30970_, _30969_, _30952_);
  and _81239_ (_30971_, _05210_, _06202_);
  or _81240_ (_30972_, _30971_, _30899_);
  or _81241_ (_30974_, _30972_, _03438_);
  and _81242_ (_30975_, _30974_, _30970_);
  or _81243_ (_30976_, _30975_, _03636_);
  and _81244_ (_30977_, _11990_, _05210_);
  or _81245_ (_30978_, _30977_, _30899_);
  or _81246_ (_30979_, _30978_, _04499_);
  and _81247_ (_30980_, _30979_, _04501_);
  and _81248_ (_30981_, _30980_, _30976_);
  or _81249_ (_30982_, _30981_, _30902_);
  and _81250_ (_30983_, _30982_, _05769_);
  nand _81251_ (_30985_, _30972_, _03754_);
  nor _81252_ (_30986_, _30985_, _30906_);
  or _81253_ (_30987_, _30986_, _30983_);
  and _81254_ (_30988_, _30987_, _03753_);
  or _81255_ (_30989_, _30899_, _05617_);
  and _81256_ (_30990_, _30910_, _03752_);
  and _81257_ (_30991_, _30990_, _30989_);
  or _81258_ (_30992_, _30991_, _03758_);
  or _81259_ (_30993_, _30992_, _30988_);
  nor _81260_ (_30994_, _11988_, _10872_);
  or _81261_ (_30996_, _30899_, _03759_);
  or _81262_ (_30997_, _30996_, _30994_);
  and _81263_ (_30998_, _30997_, _04517_);
  and _81264_ (_30999_, _30998_, _30993_);
  nor _81265_ (_31000_, _11870_, _10872_);
  or _81266_ (_31001_, _31000_, _30899_);
  and _81267_ (_31002_, _31001_, _03760_);
  or _81268_ (_31003_, _31002_, _03790_);
  or _81269_ (_31004_, _31003_, _30999_);
  or _81270_ (_31005_, _30907_, _04192_);
  and _81271_ (_31007_, _31005_, _03152_);
  and _81272_ (_31008_, _31007_, _31004_);
  and _81273_ (_31009_, _30899_, _03151_);
  or _81274_ (_31010_, _31009_, _03520_);
  or _81275_ (_31011_, _31010_, _31008_);
  or _81276_ (_31012_, _30907_, _03521_);
  and _81277_ (_31013_, _31012_, _42963_);
  and _81278_ (_31014_, _31013_, _31011_);
  or _81279_ (_43345_, _31014_, _30898_);
  and _81280_ (_31015_, _10872_, \oc8051_golden_model_1.P2 [1]);
  nor _81281_ (_31017_, _10872_, _04603_);
  or _81282_ (_31018_, _31017_, _31015_);
  and _81283_ (_31019_, _31018_, _03568_);
  and _81284_ (_31020_, _10880_, \oc8051_golden_model_1.P2 [1]);
  and _81285_ (_31021_, _12083_, _05801_);
  or _81286_ (_31022_, _31021_, _31020_);
  or _81287_ (_31023_, _31022_, _03517_);
  or _81288_ (_31024_, _05210_, \oc8051_golden_model_1.P2 [1]);
  and _81289_ (_31025_, _12252_, _05210_);
  not _81290_ (_31026_, _31025_);
  and _81291_ (_31028_, _31026_, _31024_);
  and _81292_ (_31029_, _31028_, _03570_);
  nand _81293_ (_31030_, _05210_, _03233_);
  and _81294_ (_31031_, _31030_, _31024_);
  and _81295_ (_31032_, _31031_, _04426_);
  and _81296_ (_31033_, _04427_, \oc8051_golden_model_1.P2 [1]);
  or _81297_ (_31034_, _31033_, _31032_);
  and _81298_ (_31035_, _31034_, _04444_);
  or _81299_ (_31036_, _31035_, _03516_);
  or _81300_ (_31037_, _31036_, _31029_);
  and _81301_ (_31039_, _31037_, _31023_);
  and _81302_ (_31040_, _31039_, _03983_);
  or _81303_ (_31041_, _31040_, _31019_);
  or _81304_ (_31042_, _31041_, _03575_);
  or _81305_ (_31043_, _31031_, _03583_);
  and _81306_ (_31044_, _31043_, _03513_);
  and _81307_ (_31045_, _31044_, _31042_);
  and _81308_ (_31046_, _12069_, _05801_);
  or _81309_ (_31047_, _31046_, _31020_);
  and _81310_ (_31048_, _31047_, _03512_);
  or _81311_ (_31050_, _31048_, _03505_);
  or _81312_ (_31051_, _31050_, _31045_);
  or _81313_ (_31052_, _31020_, _12098_);
  and _81314_ (_31053_, _31052_, _31022_);
  or _81315_ (_31054_, _31053_, _03506_);
  and _81316_ (_31055_, _31054_, _03500_);
  and _81317_ (_31056_, _31055_, _31051_);
  or _81318_ (_31057_, _12115_, _12069_);
  and _81319_ (_31058_, _31057_, _05801_);
  or _81320_ (_31059_, _31058_, _31020_);
  and _81321_ (_31061_, _31059_, _03499_);
  or _81322_ (_31062_, _31061_, _07314_);
  or _81323_ (_31063_, _31062_, _31056_);
  or _81324_ (_31064_, _31018_, _06039_);
  and _81325_ (_31065_, _31064_, _31063_);
  or _81326_ (_31066_, _31065_, _03479_);
  and _81327_ (_31067_, _06714_, _05210_);
  or _81328_ (_31068_, _31015_, _06044_);
  or _81329_ (_31069_, _31068_, _31067_);
  and _81330_ (_31070_, _31069_, _03474_);
  and _81331_ (_31072_, _31070_, _31066_);
  and _81332_ (_31073_, _06245_, \oc8051_golden_model_1.P1 [1]);
  and _81333_ (_31074_, _06249_, \oc8051_golden_model_1.P3 [1]);
  or _81334_ (_31075_, _31074_, _31073_);
  or _81335_ (_31076_, _31075_, _12155_);
  and _81336_ (_31077_, _06242_, \oc8051_golden_model_1.P0 [1]);
  and _81337_ (_31078_, _06214_, \oc8051_golden_model_1.P2 [1]);
  or _81338_ (_31079_, _31078_, _31077_);
  nor _81339_ (_31080_, _31079_, _31076_);
  and _81340_ (_31081_, _31080_, _12147_);
  and _81341_ (_31083_, _31081_, _12140_);
  nand _81342_ (_31084_, _31083_, _12173_);
  or _81343_ (_31085_, _31084_, _12128_);
  and _81344_ (_31086_, _31085_, _05210_);
  or _81345_ (_31087_, _31086_, _31015_);
  and _81346_ (_31088_, _31087_, _03221_);
  or _81347_ (_31089_, _31088_, _31072_);
  and _81348_ (_31090_, _31089_, _03438_);
  nand _81349_ (_31091_, _05210_, _04317_);
  and _81350_ (_31092_, _31024_, _03437_);
  and _81351_ (_31094_, _31092_, _31091_);
  or _81352_ (_31095_, _31094_, _31090_);
  and _81353_ (_31096_, _31095_, _04499_);
  or _81354_ (_31097_, _12191_, _10872_);
  and _81355_ (_31098_, _31024_, _03636_);
  and _81356_ (_31099_, _31098_, _31097_);
  or _81357_ (_31100_, _31099_, _31096_);
  and _81358_ (_31101_, _31100_, _04501_);
  or _81359_ (_31102_, _12197_, _10872_);
  and _81360_ (_31103_, _31024_, _03769_);
  and _81361_ (_31105_, _31103_, _31102_);
  or _81362_ (_31106_, _31105_, _31101_);
  and _81363_ (_31107_, _31106_, _05769_);
  or _81364_ (_31108_, _12190_, _10872_);
  and _81365_ (_31109_, _31108_, _03754_);
  and _81366_ (_31110_, _31109_, _31024_);
  or _81367_ (_31111_, _31110_, _31107_);
  and _81368_ (_31112_, _31111_, _03753_);
  or _81369_ (_31113_, _31015_, _05569_);
  and _81370_ (_31114_, _31031_, _03752_);
  and _81371_ (_31116_, _31114_, _31113_);
  or _81372_ (_31117_, _31116_, _31112_);
  and _81373_ (_31118_, _31117_, _03759_);
  or _81374_ (_31119_, _31091_, _05569_);
  and _81375_ (_31120_, _31024_, _03758_);
  and _81376_ (_31121_, _31120_, _31119_);
  or _81377_ (_31122_, _31121_, _31118_);
  and _81378_ (_31123_, _31122_, _04517_);
  or _81379_ (_31124_, _31030_, _05569_);
  and _81380_ (_31125_, _31024_, _03760_);
  and _81381_ (_31127_, _31125_, _31124_);
  or _81382_ (_31128_, _31127_, _03790_);
  or _81383_ (_31129_, _31128_, _31123_);
  or _81384_ (_31130_, _31028_, _04192_);
  and _81385_ (_31131_, _31130_, _03152_);
  and _81386_ (_31132_, _31131_, _31129_);
  and _81387_ (_31133_, _31047_, _03151_);
  or _81388_ (_31134_, _31133_, _03520_);
  or _81389_ (_31135_, _31134_, _31132_);
  or _81390_ (_31136_, _31015_, _03521_);
  or _81391_ (_31137_, _31136_, _31025_);
  and _81392_ (_31138_, _31137_, _42963_);
  and _81393_ (_31139_, _31138_, _31135_);
  nor _81394_ (_31140_, \oc8051_golden_model_1.P2 [1], rst);
  nor _81395_ (_31141_, _31140_, _00000_);
  or _81396_ (_43346_, _31141_, _31139_);
  and _81397_ (_31142_, _10872_, \oc8051_golden_model_1.P2 [2]);
  and _81398_ (_31143_, _12401_, _05210_);
  or _81399_ (_31144_, _31143_, _31142_);
  and _81400_ (_31145_, _31144_, _03769_);
  nor _81401_ (_31148_, _10872_, _05026_);
  or _81402_ (_31149_, _31148_, _31142_);
  or _81403_ (_31150_, _31149_, _06039_);
  and _81404_ (_31151_, _31149_, _03568_);
  and _81405_ (_31152_, _10880_, \oc8051_golden_model_1.P2 [2]);
  and _81406_ (_31153_, _12278_, _05801_);
  or _81407_ (_31154_, _31153_, _31152_);
  or _81408_ (_31155_, _31154_, _03517_);
  nor _81409_ (_31156_, _12282_, _10872_);
  or _81410_ (_31157_, _31156_, _31142_);
  and _81411_ (_31159_, _31157_, _03570_);
  and _81412_ (_31160_, _04427_, \oc8051_golden_model_1.P2 [2]);
  and _81413_ (_31161_, _05210_, \oc8051_golden_model_1.ACC [2]);
  or _81414_ (_31162_, _31161_, _31142_);
  and _81415_ (_31163_, _31162_, _04426_);
  or _81416_ (_31164_, _31163_, _31160_);
  and _81417_ (_31165_, _31164_, _04444_);
  or _81418_ (_31166_, _31165_, _03516_);
  or _81419_ (_31167_, _31166_, _31159_);
  and _81420_ (_31168_, _31167_, _31155_);
  and _81421_ (_31170_, _31168_, _03983_);
  or _81422_ (_31171_, _31170_, _31151_);
  or _81423_ (_31172_, _31171_, _03575_);
  or _81424_ (_31173_, _31162_, _03583_);
  and _81425_ (_31174_, _31173_, _03513_);
  and _81426_ (_31175_, _31174_, _31172_);
  and _81427_ (_31176_, _12276_, _05801_);
  or _81428_ (_31177_, _31176_, _31152_);
  and _81429_ (_31178_, _31177_, _03512_);
  or _81430_ (_31179_, _31178_, _03505_);
  or _81431_ (_31181_, _31179_, _31175_);
  or _81432_ (_31182_, _31152_, _12309_);
  and _81433_ (_31183_, _31182_, _31154_);
  or _81434_ (_31184_, _31183_, _03506_);
  and _81435_ (_31185_, _31184_, _03500_);
  and _81436_ (_31186_, _31185_, _31181_);
  or _81437_ (_31187_, _12325_, _12276_);
  and _81438_ (_31188_, _31187_, _05801_);
  or _81439_ (_31189_, _31188_, _31152_);
  and _81440_ (_31190_, _31189_, _03499_);
  or _81441_ (_31192_, _31190_, _07314_);
  or _81442_ (_31193_, _31192_, _31186_);
  and _81443_ (_31194_, _31193_, _31150_);
  or _81444_ (_31195_, _31194_, _03479_);
  and _81445_ (_31196_, _06718_, _05210_);
  or _81446_ (_31197_, _31142_, _06044_);
  or _81447_ (_31198_, _31197_, _31196_);
  and _81448_ (_31199_, _31198_, _03474_);
  and _81449_ (_31200_, _31199_, _31195_);
  and _81450_ (_31201_, _06214_, \oc8051_golden_model_1.P2 [2]);
  and _81451_ (_31203_, _06242_, \oc8051_golden_model_1.P0 [2]);
  or _81452_ (_31204_, _31203_, _12344_);
  or _81453_ (_31205_, _31204_, _31201_);
  and _81454_ (_31206_, _06245_, \oc8051_golden_model_1.P1 [2]);
  and _81455_ (_31207_, _06249_, \oc8051_golden_model_1.P3 [2]);
  or _81456_ (_31208_, _31207_, _31206_);
  nor _81457_ (_31209_, _31208_, _12345_);
  nand _81458_ (_31210_, _31209_, _12353_);
  nor _81459_ (_31211_, _31210_, _31205_);
  and _81460_ (_31212_, _31211_, _12341_);
  nand _81461_ (_31214_, _31212_, _12381_);
  or _81462_ (_31215_, _31214_, _12338_);
  and _81463_ (_31216_, _31215_, _05210_);
  or _81464_ (_31217_, _31216_, _31142_);
  and _81465_ (_31218_, _31217_, _03221_);
  or _81466_ (_31219_, _31218_, _03437_);
  or _81467_ (_31220_, _31219_, _31200_);
  and _81468_ (_31221_, _05210_, _06261_);
  or _81469_ (_31222_, _31221_, _31142_);
  or _81470_ (_31223_, _31222_, _03438_);
  and _81471_ (_31225_, _31223_, _31220_);
  or _81472_ (_31226_, _31225_, _03636_);
  and _81473_ (_31227_, _12273_, _05210_);
  or _81474_ (_31228_, _31227_, _31142_);
  or _81475_ (_31229_, _31228_, _04499_);
  and _81476_ (_31230_, _31229_, _04501_);
  and _81477_ (_31231_, _31230_, _31226_);
  or _81478_ (_31232_, _31231_, _31145_);
  and _81479_ (_31233_, _31232_, _05769_);
  or _81480_ (_31234_, _31142_, _05665_);
  and _81481_ (_31236_, _31234_, _03754_);
  and _81482_ (_31237_, _31236_, _31222_);
  or _81483_ (_31238_, _31237_, _31233_);
  and _81484_ (_31239_, _31238_, _03753_);
  and _81485_ (_31240_, _31162_, _03752_);
  and _81486_ (_31241_, _31240_, _31234_);
  or _81487_ (_31242_, _31241_, _03758_);
  or _81488_ (_31243_, _31242_, _31239_);
  nor _81489_ (_31244_, _12272_, _10872_);
  or _81490_ (_31245_, _31142_, _03759_);
  or _81491_ (_31247_, _31245_, _31244_);
  and _81492_ (_31248_, _31247_, _04517_);
  and _81493_ (_31249_, _31248_, _31243_);
  nor _81494_ (_31250_, _12400_, _10872_);
  or _81495_ (_31251_, _31250_, _31142_);
  and _81496_ (_31252_, _31251_, _03760_);
  or _81497_ (_31253_, _31252_, _03790_);
  or _81498_ (_31254_, _31253_, _31249_);
  or _81499_ (_31255_, _31157_, _04192_);
  and _81500_ (_31256_, _31255_, _03152_);
  and _81501_ (_31258_, _31256_, _31254_);
  and _81502_ (_31259_, _31177_, _03151_);
  or _81503_ (_31260_, _31259_, _03520_);
  or _81504_ (_31261_, _31260_, _31258_);
  and _81505_ (_31262_, _12456_, _05210_);
  or _81506_ (_31263_, _31142_, _03521_);
  or _81507_ (_31264_, _31263_, _31262_);
  and _81508_ (_31265_, _31264_, _42963_);
  and _81509_ (_31266_, _31265_, _31261_);
  nor _81510_ (_31267_, \oc8051_golden_model_1.P2 [2], rst);
  nor _81511_ (_31269_, _31267_, _00000_);
  or _81512_ (_43347_, _31269_, _31266_);
  and _81513_ (_31270_, _10872_, \oc8051_golden_model_1.P2 [3]);
  and _81514_ (_31271_, _12604_, _05210_);
  or _81515_ (_31272_, _31271_, _31270_);
  and _81516_ (_31273_, _31272_, _03769_);
  nor _81517_ (_31274_, _10872_, _04843_);
  or _81518_ (_31275_, _31274_, _31270_);
  or _81519_ (_31276_, _31275_, _06039_);
  nor _81520_ (_31277_, _12486_, _10872_);
  or _81521_ (_31279_, _31277_, _31270_);
  or _81522_ (_31280_, _31279_, _04444_);
  and _81523_ (_31281_, _05210_, \oc8051_golden_model_1.ACC [3]);
  or _81524_ (_31282_, _31281_, _31270_);
  and _81525_ (_31283_, _31282_, _04426_);
  and _81526_ (_31284_, _04427_, \oc8051_golden_model_1.P2 [3]);
  or _81527_ (_31285_, _31284_, _03570_);
  or _81528_ (_31286_, _31285_, _31283_);
  and _81529_ (_31287_, _31286_, _03517_);
  and _81530_ (_31288_, _31287_, _31280_);
  and _81531_ (_31290_, _10880_, \oc8051_golden_model_1.P2 [3]);
  and _81532_ (_31291_, _12490_, _05801_);
  or _81533_ (_31292_, _31291_, _31290_);
  and _81534_ (_31293_, _31292_, _03516_);
  or _81535_ (_31294_, _31293_, _03568_);
  or _81536_ (_31295_, _31294_, _31288_);
  or _81537_ (_31296_, _31275_, _03983_);
  and _81538_ (_31297_, _31296_, _31295_);
  or _81539_ (_31298_, _31297_, _03575_);
  or _81540_ (_31299_, _31282_, _03583_);
  and _81541_ (_31301_, _31299_, _03513_);
  and _81542_ (_31302_, _31301_, _31298_);
  and _81543_ (_31303_, _12500_, _05801_);
  or _81544_ (_31304_, _31303_, _31290_);
  and _81545_ (_31305_, _31304_, _03512_);
  or _81546_ (_31306_, _31305_, _03505_);
  or _81547_ (_31307_, _31306_, _31302_);
  or _81548_ (_31308_, _31290_, _12507_);
  and _81549_ (_31309_, _31308_, _31292_);
  or _81550_ (_31310_, _31309_, _03506_);
  and _81551_ (_31312_, _31310_, _03500_);
  and _81552_ (_31313_, _31312_, _31307_);
  or _81553_ (_31314_, _12500_, _12523_);
  and _81554_ (_31315_, _31314_, _05801_);
  or _81555_ (_31316_, _31315_, _31290_);
  and _81556_ (_31317_, _31316_, _03499_);
  or _81557_ (_31318_, _31317_, _07314_);
  or _81558_ (_31319_, _31318_, _31313_);
  and _81559_ (_31320_, _31319_, _31276_);
  or _81560_ (_31321_, _31320_, _03479_);
  and _81561_ (_31323_, _06717_, _05210_);
  or _81562_ (_31324_, _31270_, _06044_);
  or _81563_ (_31325_, _31324_, _31323_);
  and _81564_ (_31326_, _31325_, _03474_);
  and _81565_ (_31327_, _31326_, _31321_);
  and _81566_ (_31328_, _06214_, \oc8051_golden_model_1.P2 [3]);
  and _81567_ (_31329_, _06242_, \oc8051_golden_model_1.P0 [3]);
  or _81568_ (_31330_, _31329_, _12543_);
  or _81569_ (_31331_, _31330_, _31328_);
  and _81570_ (_31332_, _06245_, \oc8051_golden_model_1.P1 [3]);
  and _81571_ (_31334_, _06249_, \oc8051_golden_model_1.P3 [3]);
  or _81572_ (_31335_, _31334_, _31332_);
  nor _81573_ (_31336_, _31335_, _12544_);
  nand _81574_ (_31337_, _31336_, _12552_);
  nor _81575_ (_31338_, _31337_, _31331_);
  and _81576_ (_31339_, _31338_, _12540_);
  nand _81577_ (_31340_, _31339_, _12580_);
  or _81578_ (_31341_, _31340_, _12537_);
  and _81579_ (_31342_, _31341_, _05210_);
  or _81580_ (_31343_, _31342_, _31270_);
  and _81581_ (_31345_, _31343_, _03221_);
  or _81582_ (_31346_, _31345_, _03437_);
  or _81583_ (_31347_, _31346_, _31327_);
  and _81584_ (_31348_, _05210_, _06217_);
  or _81585_ (_31349_, _31348_, _31270_);
  or _81586_ (_31350_, _31349_, _03438_);
  and _81587_ (_31351_, _31350_, _31347_);
  or _81588_ (_31352_, _31351_, _03636_);
  and _81589_ (_31353_, _12598_, _05210_);
  or _81590_ (_31354_, _31353_, _31270_);
  or _81591_ (_31356_, _31354_, _04499_);
  and _81592_ (_31357_, _31356_, _04501_);
  and _81593_ (_31358_, _31357_, _31352_);
  or _81594_ (_31359_, _31358_, _31273_);
  and _81595_ (_31360_, _31359_, _05769_);
  or _81596_ (_31361_, _31270_, _05521_);
  and _81597_ (_31362_, _31361_, _03754_);
  and _81598_ (_31363_, _31362_, _31349_);
  or _81599_ (_31364_, _31363_, _31360_);
  and _81600_ (_31365_, _31364_, _03753_);
  and _81601_ (_31367_, _31282_, _03752_);
  and _81602_ (_31368_, _31367_, _31361_);
  or _81603_ (_31369_, _31368_, _03758_);
  or _81604_ (_31370_, _31369_, _31365_);
  nor _81605_ (_31371_, _12597_, _10872_);
  or _81606_ (_31372_, _31270_, _03759_);
  or _81607_ (_31373_, _31372_, _31371_);
  and _81608_ (_31374_, _31373_, _04517_);
  and _81609_ (_31375_, _31374_, _31370_);
  nor _81610_ (_31376_, _12603_, _10872_);
  or _81611_ (_31378_, _31376_, _31270_);
  and _81612_ (_31379_, _31378_, _03760_);
  or _81613_ (_31380_, _31379_, _03790_);
  or _81614_ (_31381_, _31380_, _31375_);
  or _81615_ (_31382_, _31279_, _04192_);
  and _81616_ (_31383_, _31382_, _03152_);
  and _81617_ (_31384_, _31383_, _31381_);
  and _81618_ (_31385_, _31304_, _03151_);
  or _81619_ (_31386_, _31385_, _03520_);
  or _81620_ (_31387_, _31386_, _31384_);
  and _81621_ (_31389_, _12658_, _05210_);
  or _81622_ (_31390_, _31270_, _03521_);
  or _81623_ (_31391_, _31390_, _31389_);
  and _81624_ (_31392_, _31391_, _42963_);
  and _81625_ (_31393_, _31392_, _31387_);
  nor _81626_ (_31394_, \oc8051_golden_model_1.P2 [3], rst);
  nor _81627_ (_31395_, _31394_, _00000_);
  or _81628_ (_43350_, _31395_, _31393_);
  and _81629_ (_31396_, _10872_, \oc8051_golden_model_1.P2 [4]);
  and _81630_ (_31397_, _12844_, _05210_);
  or _81631_ (_31399_, _31397_, _31396_);
  and _81632_ (_31400_, _31399_, _03769_);
  nor _81633_ (_31401_, _05712_, _10872_);
  or _81634_ (_31402_, _31401_, _31396_);
  or _81635_ (_31403_, _31402_, _06039_);
  nor _81636_ (_31404_, _12733_, _10872_);
  or _81637_ (_31405_, _31404_, _31396_);
  or _81638_ (_31406_, _31405_, _04444_);
  and _81639_ (_31407_, _05210_, \oc8051_golden_model_1.ACC [4]);
  or _81640_ (_31408_, _31407_, _31396_);
  and _81641_ (_31410_, _31408_, _04426_);
  and _81642_ (_31411_, _04427_, \oc8051_golden_model_1.P2 [4]);
  or _81643_ (_31412_, _31411_, _03570_);
  or _81644_ (_31413_, _31412_, _31410_);
  and _81645_ (_31414_, _31413_, _03517_);
  and _81646_ (_31415_, _31414_, _31406_);
  and _81647_ (_31416_, _10880_, \oc8051_golden_model_1.P2 [4]);
  and _81648_ (_31417_, _12737_, _05801_);
  or _81649_ (_31418_, _31417_, _31416_);
  and _81650_ (_31419_, _31418_, _03516_);
  or _81651_ (_31421_, _31419_, _03568_);
  or _81652_ (_31422_, _31421_, _31415_);
  or _81653_ (_31423_, _31402_, _03983_);
  and _81654_ (_31424_, _31423_, _31422_);
  or _81655_ (_31425_, _31424_, _03575_);
  or _81656_ (_31426_, _31408_, _03583_);
  and _81657_ (_31427_, _31426_, _03513_);
  and _81658_ (_31428_, _31427_, _31425_);
  and _81659_ (_31429_, _12718_, _05801_);
  or _81660_ (_31430_, _31429_, _31416_);
  and _81661_ (_31431_, _31430_, _03512_);
  or _81662_ (_31432_, _31431_, _03505_);
  or _81663_ (_31433_, _31432_, _31428_);
  or _81664_ (_31434_, _31416_, _12752_);
  and _81665_ (_31435_, _31434_, _31418_);
  or _81666_ (_31436_, _31435_, _03506_);
  and _81667_ (_31437_, _31436_, _03500_);
  and _81668_ (_31438_, _31437_, _31433_);
  or _81669_ (_31439_, _12718_, _12715_);
  and _81670_ (_31440_, _31439_, _05801_);
  or _81671_ (_31442_, _31440_, _31416_);
  and _81672_ (_31443_, _31442_, _03499_);
  or _81673_ (_31444_, _31443_, _07314_);
  or _81674_ (_31445_, _31444_, _31438_);
  and _81675_ (_31446_, _31445_, _31403_);
  or _81676_ (_31447_, _31446_, _03479_);
  and _81677_ (_31448_, _06722_, _05210_);
  or _81678_ (_31449_, _31396_, _06044_);
  or _81679_ (_31450_, _31449_, _31448_);
  and _81680_ (_31451_, _31450_, _03474_);
  and _81681_ (_31453_, _31451_, _31447_);
  and _81682_ (_31454_, _06245_, \oc8051_golden_model_1.P1 [4]);
  and _81683_ (_31455_, _06249_, \oc8051_golden_model_1.P3 [4]);
  or _81684_ (_31456_, _31455_, _31454_);
  nor _81685_ (_31457_, _31456_, _12787_);
  nand _81686_ (_31458_, _31457_, _12786_);
  or _81687_ (_31459_, _31458_, _12779_);
  and _81688_ (_31460_, _06242_, \oc8051_golden_model_1.P0 [4]);
  and _81689_ (_31461_, _06214_, \oc8051_golden_model_1.P2 [4]);
  or _81690_ (_31462_, _31461_, _12798_);
  nor _81691_ (_31464_, _31462_, _31460_);
  nand _81692_ (_31465_, _31464_, _12797_);
  nor _81693_ (_31466_, _31465_, _31459_);
  nand _81694_ (_31467_, _31466_, _12824_);
  or _81695_ (_31468_, _31467_, _12778_);
  and _81696_ (_31469_, _31468_, _05210_);
  or _81697_ (_31470_, _31469_, _31396_);
  and _81698_ (_31471_, _31470_, _03221_);
  or _81699_ (_31472_, _31471_, _03437_);
  or _81700_ (_31473_, _31472_, _31453_);
  and _81701_ (_31475_, _06233_, _05210_);
  or _81702_ (_31476_, _31475_, _31396_);
  or _81703_ (_31477_, _31476_, _03438_);
  and _81704_ (_31478_, _31477_, _31473_);
  or _81705_ (_31479_, _31478_, _03636_);
  and _81706_ (_31480_, _12711_, _05210_);
  or _81707_ (_31481_, _31480_, _31396_);
  or _81708_ (_31482_, _31481_, _04499_);
  and _81709_ (_31483_, _31482_, _04501_);
  and _81710_ (_31484_, _31483_, _31479_);
  or _81711_ (_31486_, _31484_, _31400_);
  and _81712_ (_31487_, _31486_, _05769_);
  or _81713_ (_31488_, _31396_, _05761_);
  and _81714_ (_31489_, _31488_, _03754_);
  and _81715_ (_31490_, _31489_, _31476_);
  or _81716_ (_31491_, _31490_, _31487_);
  and _81717_ (_31492_, _31491_, _03753_);
  and _81718_ (_31493_, _31408_, _03752_);
  and _81719_ (_31494_, _31493_, _31488_);
  or _81720_ (_31495_, _31494_, _03758_);
  or _81721_ (_31497_, _31495_, _31492_);
  nor _81722_ (_31498_, _12710_, _10872_);
  or _81723_ (_31499_, _31396_, _03759_);
  or _81724_ (_31500_, _31499_, _31498_);
  and _81725_ (_31501_, _31500_, _04517_);
  and _81726_ (_31502_, _31501_, _31497_);
  nor _81727_ (_31503_, _12843_, _10872_);
  or _81728_ (_31504_, _31503_, _31396_);
  and _81729_ (_31505_, _31504_, _03760_);
  or _81730_ (_31506_, _31505_, _03790_);
  or _81731_ (_31508_, _31506_, _31502_);
  or _81732_ (_31509_, _31405_, _04192_);
  and _81733_ (_31510_, _31509_, _03152_);
  and _81734_ (_31511_, _31510_, _31508_);
  and _81735_ (_31512_, _31430_, _03151_);
  or _81736_ (_31513_, _31512_, _03520_);
  or _81737_ (_31514_, _31513_, _31511_);
  and _81738_ (_31515_, _12893_, _05210_);
  or _81739_ (_31516_, _31396_, _03521_);
  or _81740_ (_31517_, _31516_, _31515_);
  and _81741_ (_31519_, _31517_, _42963_);
  and _81742_ (_31520_, _31519_, _31514_);
  nor _81743_ (_31521_, \oc8051_golden_model_1.P2 [4], rst);
  nor _81744_ (_31522_, _31521_, _00000_);
  or _81745_ (_43351_, _31522_, _31520_);
  and _81746_ (_31523_, _10872_, \oc8051_golden_model_1.P2 [5]);
  and _81747_ (_31524_, _13042_, _05210_);
  or _81748_ (_31525_, _31524_, _31523_);
  and _81749_ (_31526_, _31525_, _03769_);
  nor _81750_ (_31527_, _05422_, _10872_);
  or _81751_ (_31529_, _31527_, _31523_);
  or _81752_ (_31530_, _31529_, _06039_);
  nor _81753_ (_31531_, _12930_, _10872_);
  or _81754_ (_31532_, _31531_, _31523_);
  or _81755_ (_31533_, _31532_, _04444_);
  and _81756_ (_31534_, _05210_, \oc8051_golden_model_1.ACC [5]);
  or _81757_ (_31535_, _31534_, _31523_);
  and _81758_ (_31536_, _31535_, _04426_);
  and _81759_ (_31537_, _04427_, \oc8051_golden_model_1.P2 [5]);
  or _81760_ (_31538_, _31537_, _03570_);
  or _81761_ (_31540_, _31538_, _31536_);
  and _81762_ (_31541_, _31540_, _03517_);
  and _81763_ (_31542_, _31541_, _31533_);
  and _81764_ (_31543_, _10880_, \oc8051_golden_model_1.P2 [5]);
  and _81765_ (_31544_, _12934_, _05801_);
  or _81766_ (_31545_, _31544_, _31543_);
  and _81767_ (_31546_, _31545_, _03516_);
  or _81768_ (_31547_, _31546_, _03568_);
  or _81769_ (_31548_, _31547_, _31542_);
  or _81770_ (_31549_, _31529_, _03983_);
  and _81771_ (_31551_, _31549_, _31548_);
  or _81772_ (_31552_, _31551_, _03575_);
  or _81773_ (_31553_, _31535_, _03583_);
  and _81774_ (_31554_, _31553_, _03513_);
  and _81775_ (_31555_, _31554_, _31552_);
  and _81776_ (_31556_, _12914_, _05801_);
  or _81777_ (_31557_, _31556_, _31543_);
  and _81778_ (_31558_, _31557_, _03512_);
  or _81779_ (_31559_, _31558_, _03505_);
  or _81780_ (_31560_, _31559_, _31555_);
  or _81781_ (_31562_, _31543_, _12949_);
  and _81782_ (_31563_, _31562_, _31545_);
  or _81783_ (_31564_, _31563_, _03506_);
  and _81784_ (_31565_, _31564_, _03500_);
  and _81785_ (_31566_, _31565_, _31560_);
  or _81786_ (_31567_, _12914_, _12911_);
  and _81787_ (_31568_, _31567_, _05801_);
  or _81788_ (_31569_, _31568_, _31543_);
  and _81789_ (_31570_, _31569_, _03499_);
  or _81790_ (_31571_, _31570_, _07314_);
  or _81791_ (_31573_, _31571_, _31566_);
  and _81792_ (_31574_, _31573_, _31530_);
  or _81793_ (_31575_, _31574_, _03479_);
  and _81794_ (_31576_, _06721_, _05210_);
  or _81795_ (_31577_, _31523_, _06044_);
  or _81796_ (_31578_, _31577_, _31576_);
  and _81797_ (_31579_, _31578_, _03474_);
  and _81798_ (_31580_, _31579_, _31575_);
  and _81799_ (_31581_, _06245_, \oc8051_golden_model_1.P1 [5]);
  and _81800_ (_31582_, _06249_, \oc8051_golden_model_1.P3 [5]);
  or _81801_ (_31584_, _31582_, _31581_);
  or _81802_ (_31585_, _31584_, _12983_);
  and _81803_ (_31586_, _06242_, \oc8051_golden_model_1.P0 [5]);
  and _81804_ (_31587_, _06214_, \oc8051_golden_model_1.P2 [5]);
  or _81805_ (_31588_, _31587_, _31586_);
  nor _81806_ (_31589_, _31588_, _31585_);
  and _81807_ (_31590_, _31589_, _13001_);
  and _81808_ (_31591_, _31590_, _12982_);
  nand _81809_ (_31592_, _31591_, _13018_);
  or _81810_ (_31593_, _31592_, _12975_);
  and _81811_ (_31595_, _31593_, _05210_);
  or _81812_ (_31596_, _31595_, _31523_);
  and _81813_ (_31597_, _31596_, _03221_);
  or _81814_ (_31598_, _31597_, _03437_);
  or _81815_ (_31599_, _31598_, _31580_);
  and _81816_ (_31600_, _06211_, _05210_);
  or _81817_ (_31601_, _31600_, _31523_);
  or _81818_ (_31602_, _31601_, _03438_);
  and _81819_ (_31603_, _31602_, _31599_);
  or _81820_ (_31604_, _31603_, _03636_);
  and _81821_ (_31606_, _13036_, _05210_);
  or _81822_ (_31607_, _31606_, _31523_);
  or _81823_ (_31608_, _31607_, _04499_);
  and _81824_ (_31609_, _31608_, _04501_);
  and _81825_ (_31610_, _31609_, _31604_);
  or _81826_ (_31611_, _31610_, _31526_);
  and _81827_ (_31612_, _31611_, _05769_);
  or _81828_ (_31613_, _31523_, _05472_);
  and _81829_ (_31614_, _31613_, _03754_);
  and _81830_ (_31615_, _31614_, _31601_);
  or _81831_ (_31617_, _31615_, _31612_);
  and _81832_ (_31618_, _31617_, _03753_);
  and _81833_ (_31619_, _31535_, _03752_);
  and _81834_ (_31620_, _31619_, _31613_);
  or _81835_ (_31621_, _31620_, _03758_);
  or _81836_ (_31622_, _31621_, _31618_);
  nor _81837_ (_31623_, _13035_, _10872_);
  or _81838_ (_31624_, _31523_, _03759_);
  or _81839_ (_31625_, _31624_, _31623_);
  and _81840_ (_31626_, _31625_, _04517_);
  and _81841_ (_31628_, _31626_, _31622_);
  nor _81842_ (_31629_, _13041_, _10872_);
  or _81843_ (_31630_, _31629_, _31523_);
  and _81844_ (_31631_, _31630_, _03760_);
  or _81845_ (_31632_, _31631_, _03790_);
  or _81846_ (_31633_, _31632_, _31628_);
  or _81847_ (_31634_, _31532_, _04192_);
  and _81848_ (_31635_, _31634_, _03152_);
  and _81849_ (_31636_, _31635_, _31633_);
  and _81850_ (_31637_, _31557_, _03151_);
  or _81851_ (_31639_, _31637_, _03520_);
  or _81852_ (_31640_, _31639_, _31636_);
  and _81853_ (_31641_, _13097_, _05210_);
  or _81854_ (_31642_, _31523_, _03521_);
  or _81855_ (_31643_, _31642_, _31641_);
  and _81856_ (_31644_, _31643_, _42963_);
  and _81857_ (_31645_, _31644_, _31640_);
  nor _81858_ (_31646_, \oc8051_golden_model_1.P2 [5], rst);
  nor _81859_ (_31647_, _31646_, _00000_);
  or _81860_ (_43352_, _31647_, _31645_);
  and _81861_ (_31649_, _10872_, \oc8051_golden_model_1.P2 [6]);
  and _81862_ (_31650_, _13259_, _05210_);
  or _81863_ (_31651_, _31650_, _31649_);
  and _81864_ (_31652_, _31651_, _03769_);
  nor _81865_ (_31653_, _05327_, _10872_);
  or _81866_ (_31654_, _31653_, _31649_);
  or _81867_ (_31655_, _31654_, _06039_);
  nor _81868_ (_31656_, _13122_, _10872_);
  or _81869_ (_31657_, _31656_, _31649_);
  or _81870_ (_31658_, _31657_, _04444_);
  and _81871_ (_31660_, _05210_, \oc8051_golden_model_1.ACC [6]);
  or _81872_ (_31661_, _31660_, _31649_);
  and _81873_ (_31662_, _31661_, _04426_);
  and _81874_ (_31663_, _04427_, \oc8051_golden_model_1.P2 [6]);
  or _81875_ (_31664_, _31663_, _03570_);
  or _81876_ (_31665_, _31664_, _31662_);
  and _81877_ (_31666_, _31665_, _03517_);
  and _81878_ (_31667_, _31666_, _31658_);
  and _81879_ (_31668_, _10880_, \oc8051_golden_model_1.P2 [6]);
  and _81880_ (_31669_, _13145_, _05801_);
  or _81881_ (_31671_, _31669_, _31668_);
  and _81882_ (_31672_, _31671_, _03516_);
  or _81883_ (_31673_, _31672_, _03568_);
  or _81884_ (_31674_, _31673_, _31667_);
  or _81885_ (_31675_, _31654_, _03983_);
  and _81886_ (_31676_, _31675_, _31674_);
  or _81887_ (_31677_, _31676_, _03575_);
  or _81888_ (_31678_, _31661_, _03583_);
  and _81889_ (_31679_, _31678_, _03513_);
  and _81890_ (_31680_, _31679_, _31677_);
  and _81891_ (_31682_, _13130_, _05801_);
  or _81892_ (_31683_, _31682_, _31668_);
  and _81893_ (_31684_, _31683_, _03512_);
  or _81894_ (_31685_, _31684_, _03505_);
  or _81895_ (_31686_, _31685_, _31680_);
  or _81896_ (_31687_, _31668_, _13160_);
  and _81897_ (_31688_, _31687_, _31671_);
  or _81898_ (_31689_, _31688_, _03506_);
  and _81899_ (_31690_, _31689_, _03500_);
  and _81900_ (_31691_, _31690_, _31686_);
  or _81901_ (_31693_, _13177_, _13130_);
  and _81902_ (_31694_, _31693_, _05801_);
  or _81903_ (_31695_, _31694_, _31668_);
  and _81904_ (_31696_, _31695_, _03499_);
  or _81905_ (_31697_, _31696_, _07314_);
  or _81906_ (_31698_, _31697_, _31691_);
  and _81907_ (_31699_, _31698_, _31655_);
  or _81908_ (_31700_, _31699_, _03479_);
  and _81909_ (_31701_, _06713_, _05210_);
  or _81910_ (_31702_, _31649_, _06044_);
  or _81911_ (_31704_, _31702_, _31701_);
  and _81912_ (_31705_, _31704_, _03474_);
  and _81913_ (_31706_, _31705_, _31700_);
  and _81914_ (_31707_, _06245_, \oc8051_golden_model_1.P1 [6]);
  and _81915_ (_31708_, _06249_, \oc8051_golden_model_1.P3 [6]);
  or _81916_ (_31709_, _31708_, _31707_);
  or _81917_ (_31710_, _31709_, _13199_);
  and _81918_ (_31711_, _06242_, \oc8051_golden_model_1.P0 [6]);
  and _81919_ (_31712_, _06214_, \oc8051_golden_model_1.P2 [6]);
  or _81920_ (_31713_, _31712_, _31711_);
  nor _81921_ (_31714_, _31713_, _31710_);
  and _81922_ (_31715_, _31714_, _13217_);
  and _81923_ (_31716_, _31715_, _13198_);
  nand _81924_ (_31717_, _31716_, _13234_);
  or _81925_ (_31718_, _31717_, _13191_);
  and _81926_ (_31719_, _31718_, _05210_);
  or _81927_ (_31720_, _31719_, _31649_);
  and _81928_ (_31721_, _31720_, _03221_);
  or _81929_ (_31722_, _31721_, _03437_);
  or _81930_ (_31723_, _31722_, _31706_);
  and _81931_ (_31726_, _13244_, _05210_);
  or _81932_ (_31727_, _31726_, _31649_);
  or _81933_ (_31728_, _31727_, _03438_);
  and _81934_ (_31729_, _31728_, _31723_);
  or _81935_ (_31730_, _31729_, _03636_);
  and _81936_ (_31731_, _13253_, _05210_);
  or _81937_ (_31732_, _31731_, _31649_);
  or _81938_ (_31733_, _31732_, _04499_);
  and _81939_ (_31734_, _31733_, _04501_);
  and _81940_ (_31735_, _31734_, _31730_);
  or _81941_ (_31737_, _31735_, _31652_);
  and _81942_ (_31738_, _31737_, _05769_);
  or _81943_ (_31739_, _31649_, _05377_);
  and _81944_ (_31740_, _31739_, _03754_);
  and _81945_ (_31741_, _31740_, _31727_);
  or _81946_ (_31742_, _31741_, _31738_);
  and _81947_ (_31743_, _31742_, _03753_);
  and _81948_ (_31744_, _31661_, _03752_);
  and _81949_ (_31745_, _31744_, _31739_);
  or _81950_ (_31746_, _31745_, _03758_);
  or _81951_ (_31748_, _31746_, _31743_);
  nor _81952_ (_31749_, _13251_, _10872_);
  or _81953_ (_31750_, _31649_, _03759_);
  or _81954_ (_31751_, _31750_, _31749_);
  and _81955_ (_31752_, _31751_, _04517_);
  and _81956_ (_31753_, _31752_, _31748_);
  nor _81957_ (_31754_, _13258_, _10872_);
  or _81958_ (_31755_, _31754_, _31649_);
  and _81959_ (_31756_, _31755_, _03760_);
  or _81960_ (_31757_, _31756_, _03790_);
  or _81961_ (_31759_, _31757_, _31753_);
  or _81962_ (_31760_, _31657_, _04192_);
  and _81963_ (_31761_, _31760_, _03152_);
  and _81964_ (_31762_, _31761_, _31759_);
  and _81965_ (_31763_, _31683_, _03151_);
  or _81966_ (_31764_, _31763_, _03520_);
  or _81967_ (_31765_, _31764_, _31762_);
  and _81968_ (_31766_, _13312_, _05210_);
  or _81969_ (_31767_, _31649_, _03521_);
  or _81970_ (_31768_, _31767_, _31766_);
  and _81971_ (_31770_, _31768_, _42963_);
  and _81972_ (_31771_, _31770_, _31765_);
  nor _81973_ (_31772_, \oc8051_golden_model_1.P2 [6], rst);
  nor _81974_ (_31773_, _31772_, _00000_);
  or _81975_ (_43353_, _31773_, _31771_);
  and _81976_ (_31774_, _10989_, \oc8051_golden_model_1.P3 [0]);
  and _81977_ (_31775_, _11995_, _05200_);
  or _81978_ (_31776_, _31775_, _31774_);
  and _81979_ (_31777_, _31776_, _03769_);
  and _81980_ (_31778_, _05941_, _05200_);
  or _81981_ (_31780_, _31778_, _31774_);
  and _81982_ (_31781_, _31780_, _03570_);
  and _81983_ (_31782_, _04427_, \oc8051_golden_model_1.P3 [0]);
  and _81984_ (_31783_, _05200_, \oc8051_golden_model_1.ACC [0]);
  or _81985_ (_31784_, _31783_, _31774_);
  and _81986_ (_31785_, _31784_, _04426_);
  or _81987_ (_31786_, _31785_, _31782_);
  and _81988_ (_31787_, _31786_, _04444_);
  or _81989_ (_31788_, _31787_, _03516_);
  or _81990_ (_31789_, _31788_, _31781_);
  and _81991_ (_31791_, _11887_, _05796_);
  and _81992_ (_31792_, _10997_, \oc8051_golden_model_1.P3 [0]);
  or _81993_ (_31793_, _31792_, _03517_);
  or _81994_ (_31794_, _31793_, _31791_);
  and _81995_ (_31795_, _31794_, _03983_);
  and _81996_ (_31796_, _31795_, _31789_);
  and _81997_ (_31797_, _05200_, _04419_);
  or _81998_ (_31798_, _31797_, _31774_);
  and _81999_ (_31799_, _31798_, _03568_);
  or _82000_ (_31800_, _31799_, _03575_);
  or _82001_ (_31802_, _31800_, _31796_);
  or _82002_ (_31803_, _31784_, _03583_);
  and _82003_ (_31804_, _31803_, _03513_);
  and _82004_ (_31805_, _31804_, _31802_);
  and _82005_ (_31806_, _31774_, _03512_);
  or _82006_ (_31807_, _31806_, _03505_);
  or _82007_ (_31808_, _31807_, _31805_);
  or _82008_ (_31809_, _31780_, _03506_);
  and _82009_ (_31810_, _31809_, _03500_);
  and _82010_ (_31811_, _31810_, _31808_);
  and _82011_ (_31813_, _30938_, _05796_);
  or _82012_ (_31814_, _31813_, _31792_);
  and _82013_ (_31815_, _31814_, _03499_);
  or _82014_ (_31816_, _31815_, _07314_);
  or _82015_ (_31817_, _31816_, _31811_);
  or _82016_ (_31818_, _31798_, _06039_);
  and _82017_ (_31819_, _31818_, _31817_);
  or _82018_ (_31820_, _31819_, _03479_);
  and _82019_ (_31821_, _06715_, _05200_);
  or _82020_ (_31822_, _31774_, _06044_);
  or _82021_ (_31824_, _31822_, _31821_);
  and _82022_ (_31825_, _31824_, _03474_);
  and _82023_ (_31826_, _31825_, _31820_);
  and _82024_ (_31827_, _30965_, _05200_);
  or _82025_ (_31828_, _31827_, _31774_);
  and _82026_ (_31829_, _31828_, _03221_);
  or _82027_ (_31830_, _31829_, _03437_);
  or _82028_ (_31831_, _31830_, _31826_);
  and _82029_ (_31832_, _05200_, _06202_);
  or _82030_ (_31833_, _31832_, _31774_);
  or _82031_ (_31835_, _31833_, _03438_);
  and _82032_ (_31836_, _31835_, _31831_);
  or _82033_ (_31837_, _31836_, _03636_);
  and _82034_ (_31838_, _11990_, _05200_);
  or _82035_ (_31839_, _31838_, _31774_);
  or _82036_ (_31840_, _31839_, _04499_);
  and _82037_ (_31841_, _31840_, _04501_);
  and _82038_ (_31842_, _31841_, _31837_);
  or _82039_ (_31843_, _31842_, _31777_);
  and _82040_ (_31844_, _31843_, _05769_);
  nand _82041_ (_31846_, _31833_, _03754_);
  nor _82042_ (_31847_, _31846_, _31778_);
  or _82043_ (_31848_, _31847_, _31844_);
  and _82044_ (_31849_, _31848_, _03753_);
  or _82045_ (_31850_, _31774_, _05617_);
  and _82046_ (_31851_, _31784_, _03752_);
  and _82047_ (_31852_, _31851_, _31850_);
  or _82048_ (_31853_, _31852_, _03758_);
  or _82049_ (_31854_, _31853_, _31849_);
  nor _82050_ (_31855_, _11988_, _10989_);
  or _82051_ (_31857_, _31774_, _03759_);
  or _82052_ (_31858_, _31857_, _31855_);
  and _82053_ (_31859_, _31858_, _04517_);
  and _82054_ (_31860_, _31859_, _31854_);
  nor _82055_ (_31861_, _11870_, _10989_);
  or _82056_ (_31862_, _31861_, _31774_);
  and _82057_ (_31863_, _31862_, _03760_);
  or _82058_ (_31864_, _31863_, _03790_);
  or _82059_ (_31865_, _31864_, _31860_);
  or _82060_ (_31866_, _31780_, _04192_);
  and _82061_ (_31868_, _31866_, _03152_);
  and _82062_ (_31869_, _31868_, _31865_);
  and _82063_ (_31870_, _31774_, _03151_);
  or _82064_ (_31871_, _31870_, _03520_);
  or _82065_ (_31872_, _31871_, _31869_);
  or _82066_ (_31873_, _31780_, _03521_);
  and _82067_ (_31874_, _31873_, _42963_);
  and _82068_ (_31875_, _31874_, _31872_);
  nor _82069_ (_31876_, \oc8051_golden_model_1.P3 [0], rst);
  nor _82070_ (_31877_, _31876_, _00000_);
  or _82071_ (_43355_, _31877_, _31875_);
  or _82072_ (_31879_, _05200_, \oc8051_golden_model_1.P3 [1]);
  and _82073_ (_31880_, _12252_, _05200_);
  not _82074_ (_31881_, _31880_);
  and _82075_ (_31882_, _31881_, _31879_);
  or _82076_ (_31883_, _31882_, _04444_);
  nand _82077_ (_31884_, _05200_, _03233_);
  and _82078_ (_31885_, _31884_, _31879_);
  and _82079_ (_31886_, _31885_, _04426_);
  and _82080_ (_31887_, _04427_, \oc8051_golden_model_1.P3 [1]);
  or _82081_ (_31889_, _31887_, _03570_);
  or _82082_ (_31890_, _31889_, _31886_);
  and _82083_ (_31891_, _31890_, _03517_);
  and _82084_ (_31892_, _31891_, _31883_);
  and _82085_ (_31893_, _12083_, _05796_);
  and _82086_ (_31894_, _10997_, \oc8051_golden_model_1.P3 [1]);
  or _82087_ (_31895_, _31894_, _03568_);
  or _82088_ (_31896_, _31895_, _31893_);
  and _82089_ (_31897_, _31896_, _14165_);
  or _82090_ (_31898_, _31897_, _31892_);
  and _82091_ (_31900_, _10989_, \oc8051_golden_model_1.P3 [1]);
  nor _82092_ (_31901_, _10989_, _04603_);
  or _82093_ (_31902_, _31901_, _31900_);
  or _82094_ (_31903_, _31902_, _03983_);
  and _82095_ (_31904_, _31903_, _31898_);
  or _82096_ (_31905_, _31904_, _03575_);
  or _82097_ (_31906_, _31885_, _03583_);
  and _82098_ (_31907_, _31906_, _03513_);
  and _82099_ (_31908_, _31907_, _31905_);
  and _82100_ (_31909_, _12069_, _05796_);
  or _82101_ (_31911_, _31909_, _31894_);
  and _82102_ (_31912_, _31911_, _03512_);
  or _82103_ (_31913_, _31912_, _03505_);
  or _82104_ (_31914_, _31913_, _31908_);
  and _82105_ (_31915_, _31893_, _12098_);
  or _82106_ (_31916_, _31894_, _03506_);
  or _82107_ (_31917_, _31916_, _31915_);
  and _82108_ (_31918_, _31917_, _31914_);
  and _82109_ (_31919_, _31918_, _03500_);
  and _82110_ (_31920_, _31057_, _05796_);
  or _82111_ (_31922_, _31894_, _31920_);
  and _82112_ (_31923_, _31922_, _03499_);
  or _82113_ (_31924_, _31923_, _07314_);
  or _82114_ (_31925_, _31924_, _31919_);
  or _82115_ (_31926_, _31902_, _06039_);
  and _82116_ (_31927_, _31926_, _31925_);
  or _82117_ (_31928_, _31927_, _03479_);
  and _82118_ (_31929_, _06714_, _05200_);
  or _82119_ (_31930_, _31900_, _06044_);
  or _82120_ (_31931_, _31930_, _31929_);
  and _82121_ (_31933_, _31931_, _03474_);
  and _82122_ (_31934_, _31933_, _31928_);
  and _82123_ (_31935_, _31085_, _05200_);
  or _82124_ (_31936_, _31935_, _31900_);
  and _82125_ (_31937_, _31936_, _03221_);
  or _82126_ (_31938_, _31937_, _31934_);
  and _82127_ (_31939_, _31938_, _03438_);
  nand _82128_ (_31940_, _05200_, _04317_);
  and _82129_ (_31941_, _31879_, _03437_);
  and _82130_ (_31942_, _31941_, _31940_);
  or _82131_ (_31944_, _31942_, _31939_);
  and _82132_ (_31945_, _31944_, _04499_);
  or _82133_ (_31946_, _12191_, _10989_);
  and _82134_ (_31947_, _31879_, _03636_);
  and _82135_ (_31948_, _31947_, _31946_);
  or _82136_ (_31949_, _31948_, _31945_);
  and _82137_ (_31950_, _31949_, _04501_);
  or _82138_ (_31951_, _12197_, _10989_);
  and _82139_ (_31952_, _31879_, _03769_);
  and _82140_ (_31953_, _31952_, _31951_);
  or _82141_ (_31955_, _31953_, _31950_);
  and _82142_ (_31956_, _31955_, _05769_);
  or _82143_ (_31957_, _12190_, _10989_);
  and _82144_ (_31958_, _31957_, _03754_);
  and _82145_ (_31959_, _31958_, _31879_);
  or _82146_ (_31960_, _31959_, _31956_);
  and _82147_ (_31961_, _31960_, _03753_);
  or _82148_ (_31962_, _31900_, _05569_);
  and _82149_ (_31963_, _31885_, _03752_);
  and _82150_ (_31964_, _31963_, _31962_);
  or _82151_ (_31966_, _31964_, _31961_);
  and _82152_ (_31967_, _31966_, _03759_);
  or _82153_ (_31968_, _31940_, _05569_);
  and _82154_ (_31969_, _31879_, _03758_);
  and _82155_ (_31970_, _31969_, _31968_);
  or _82156_ (_31971_, _31970_, _31967_);
  and _82157_ (_31972_, _31971_, _04517_);
  or _82158_ (_31973_, _31884_, _05569_);
  and _82159_ (_31974_, _31879_, _03760_);
  and _82160_ (_31975_, _31974_, _31973_);
  or _82161_ (_31977_, _31975_, _03790_);
  or _82162_ (_31978_, _31977_, _31972_);
  or _82163_ (_31979_, _31882_, _04192_);
  and _82164_ (_31980_, _31979_, _03152_);
  and _82165_ (_31981_, _31980_, _31978_);
  and _82166_ (_31982_, _31911_, _03151_);
  or _82167_ (_31983_, _31982_, _03520_);
  or _82168_ (_31984_, _31983_, _31981_);
  or _82169_ (_31985_, _31900_, _03521_);
  or _82170_ (_31986_, _31985_, _31880_);
  and _82171_ (_31988_, _31986_, _42963_);
  and _82172_ (_31989_, _31988_, _31984_);
  nor _82173_ (_31990_, \oc8051_golden_model_1.P3 [1], rst);
  nor _82174_ (_31991_, _31990_, _00000_);
  or _82175_ (_43356_, _31991_, _31989_);
  and _82176_ (_31992_, _10989_, \oc8051_golden_model_1.P3 [2]);
  and _82177_ (_31993_, _12401_, _05200_);
  or _82178_ (_31994_, _31993_, _31992_);
  and _82179_ (_31995_, _31994_, _03769_);
  nor _82180_ (_31996_, _10989_, _05026_);
  or _82181_ (_31998_, _31996_, _31992_);
  or _82182_ (_31999_, _31998_, _06039_);
  and _82183_ (_32000_, _31998_, _03568_);
  and _82184_ (_32001_, _10997_, \oc8051_golden_model_1.P3 [2]);
  and _82185_ (_32002_, _12278_, _05796_);
  or _82186_ (_32003_, _32002_, _32001_);
  or _82187_ (_32004_, _32003_, _03517_);
  nor _82188_ (_32005_, _12282_, _10989_);
  or _82189_ (_32006_, _32005_, _31992_);
  and _82190_ (_32007_, _32006_, _03570_);
  and _82191_ (_32009_, _04427_, \oc8051_golden_model_1.P3 [2]);
  and _82192_ (_32010_, _05200_, \oc8051_golden_model_1.ACC [2]);
  or _82193_ (_32011_, _32010_, _31992_);
  and _82194_ (_32012_, _32011_, _04426_);
  or _82195_ (_32013_, _32012_, _32009_);
  and _82196_ (_32014_, _32013_, _04444_);
  or _82197_ (_32015_, _32014_, _03516_);
  or _82198_ (_32016_, _32015_, _32007_);
  and _82199_ (_32017_, _32016_, _32004_);
  and _82200_ (_32018_, _32017_, _03983_);
  or _82201_ (_32020_, _32018_, _32000_);
  or _82202_ (_32021_, _32020_, _03575_);
  or _82203_ (_32022_, _32011_, _03583_);
  and _82204_ (_32023_, _32022_, _03513_);
  and _82205_ (_32024_, _32023_, _32021_);
  and _82206_ (_32025_, _12276_, _05796_);
  or _82207_ (_32026_, _32025_, _32001_);
  and _82208_ (_32027_, _32026_, _03512_);
  or _82209_ (_32028_, _32027_, _03505_);
  or _82210_ (_32029_, _32028_, _32024_);
  or _82211_ (_32031_, _32001_, _12309_);
  and _82212_ (_32032_, _32031_, _32003_);
  or _82213_ (_32033_, _32032_, _03506_);
  and _82214_ (_32034_, _32033_, _03500_);
  and _82215_ (_32035_, _32034_, _32029_);
  and _82216_ (_32036_, _31187_, _05796_);
  or _82217_ (_32037_, _32036_, _32001_);
  and _82218_ (_32038_, _32037_, _03499_);
  or _82219_ (_32039_, _32038_, _07314_);
  or _82220_ (_32040_, _32039_, _32035_);
  and _82221_ (_32042_, _32040_, _31999_);
  or _82222_ (_32043_, _32042_, _03479_);
  and _82223_ (_32044_, _06718_, _05200_);
  or _82224_ (_32045_, _31992_, _06044_);
  or _82225_ (_32046_, _32045_, _32044_);
  and _82226_ (_32047_, _32046_, _03474_);
  and _82227_ (_32048_, _32047_, _32043_);
  and _82228_ (_32049_, _31215_, _05200_);
  or _82229_ (_32050_, _32049_, _31992_);
  and _82230_ (_32051_, _32050_, _03221_);
  or _82231_ (_32053_, _32051_, _03437_);
  or _82232_ (_32054_, _32053_, _32048_);
  and _82233_ (_32055_, _05200_, _06261_);
  or _82234_ (_32056_, _32055_, _31992_);
  or _82235_ (_32057_, _32056_, _03438_);
  and _82236_ (_32058_, _32057_, _32054_);
  or _82237_ (_32059_, _32058_, _03636_);
  and _82238_ (_32060_, _12273_, _05200_);
  or _82239_ (_32061_, _32060_, _31992_);
  or _82240_ (_32062_, _32061_, _04499_);
  and _82241_ (_32064_, _32062_, _04501_);
  and _82242_ (_32065_, _32064_, _32059_);
  or _82243_ (_32066_, _32065_, _31995_);
  and _82244_ (_32067_, _32066_, _05769_);
  or _82245_ (_32068_, _31992_, _05665_);
  and _82246_ (_32069_, _32068_, _03754_);
  and _82247_ (_32070_, _32069_, _32056_);
  or _82248_ (_32071_, _32070_, _32067_);
  and _82249_ (_32072_, _32071_, _03753_);
  and _82250_ (_32073_, _32011_, _03752_);
  and _82251_ (_32075_, _32073_, _32068_);
  or _82252_ (_32076_, _32075_, _03758_);
  or _82253_ (_32077_, _32076_, _32072_);
  nor _82254_ (_32078_, _12272_, _10989_);
  or _82255_ (_32079_, _31992_, _03759_);
  or _82256_ (_32080_, _32079_, _32078_);
  and _82257_ (_32081_, _32080_, _04517_);
  and _82258_ (_32082_, _32081_, _32077_);
  nor _82259_ (_32083_, _12400_, _10989_);
  or _82260_ (_32084_, _32083_, _31992_);
  and _82261_ (_32086_, _32084_, _03760_);
  or _82262_ (_32087_, _32086_, _03790_);
  or _82263_ (_32088_, _32087_, _32082_);
  or _82264_ (_32089_, _32006_, _04192_);
  and _82265_ (_32090_, _32089_, _03152_);
  and _82266_ (_32091_, _32090_, _32088_);
  and _82267_ (_32092_, _32026_, _03151_);
  or _82268_ (_32093_, _32092_, _03520_);
  or _82269_ (_32094_, _32093_, _32091_);
  and _82270_ (_32095_, _12456_, _05200_);
  or _82271_ (_32097_, _31992_, _03521_);
  or _82272_ (_32098_, _32097_, _32095_);
  and _82273_ (_32099_, _32098_, _42963_);
  and _82274_ (_32100_, _32099_, _32094_);
  nor _82275_ (_32101_, \oc8051_golden_model_1.P3 [2], rst);
  nor _82276_ (_32102_, _32101_, _00000_);
  or _82277_ (_43357_, _32102_, _32100_);
  and _82278_ (_32103_, _10989_, \oc8051_golden_model_1.P3 [3]);
  and _82279_ (_32104_, _12604_, _05200_);
  or _82280_ (_32105_, _32104_, _32103_);
  and _82281_ (_32107_, _32105_, _03769_);
  nor _82282_ (_32108_, _10989_, _04843_);
  or _82283_ (_32109_, _32108_, _32103_);
  or _82284_ (_32110_, _32109_, _06039_);
  nor _82285_ (_32111_, _12486_, _10989_);
  or _82286_ (_32112_, _32111_, _32103_);
  or _82287_ (_32113_, _32112_, _04444_);
  and _82288_ (_32114_, _05200_, \oc8051_golden_model_1.ACC [3]);
  or _82289_ (_32115_, _32114_, _32103_);
  and _82290_ (_32116_, _32115_, _04426_);
  and _82291_ (_32118_, _04427_, \oc8051_golden_model_1.P3 [3]);
  or _82292_ (_32119_, _32118_, _03570_);
  or _82293_ (_32120_, _32119_, _32116_);
  and _82294_ (_32121_, _32120_, _03517_);
  and _82295_ (_32122_, _32121_, _32113_);
  and _82296_ (_32123_, _10997_, \oc8051_golden_model_1.P3 [3]);
  and _82297_ (_32124_, _12490_, _05796_);
  or _82298_ (_32125_, _32124_, _32123_);
  and _82299_ (_32126_, _32125_, _03516_);
  or _82300_ (_32127_, _32126_, _03568_);
  or _82301_ (_32129_, _32127_, _32122_);
  or _82302_ (_32130_, _32109_, _03983_);
  and _82303_ (_32131_, _32130_, _32129_);
  or _82304_ (_32132_, _32131_, _03575_);
  or _82305_ (_32133_, _32115_, _03583_);
  and _82306_ (_32134_, _32133_, _03513_);
  and _82307_ (_32135_, _32134_, _32132_);
  and _82308_ (_32136_, _12500_, _05796_);
  or _82309_ (_32137_, _32136_, _32123_);
  and _82310_ (_32138_, _32137_, _03512_);
  or _82311_ (_32140_, _32138_, _03505_);
  or _82312_ (_32141_, _32140_, _32135_);
  or _82313_ (_32142_, _32123_, _12507_);
  and _82314_ (_32143_, _32142_, _32125_);
  or _82315_ (_32144_, _32143_, _03506_);
  and _82316_ (_32145_, _32144_, _03500_);
  and _82317_ (_32146_, _32145_, _32141_);
  and _82318_ (_32147_, _31314_, _05796_);
  or _82319_ (_32148_, _32147_, _32123_);
  and _82320_ (_32149_, _32148_, _03499_);
  or _82321_ (_32151_, _32149_, _07314_);
  or _82322_ (_32152_, _32151_, _32146_);
  and _82323_ (_32153_, _32152_, _32110_);
  or _82324_ (_32154_, _32153_, _03479_);
  and _82325_ (_32155_, _06717_, _05200_);
  or _82326_ (_32156_, _32103_, _06044_);
  or _82327_ (_32157_, _32156_, _32155_);
  and _82328_ (_32158_, _32157_, _03474_);
  and _82329_ (_32159_, _32158_, _32154_);
  and _82330_ (_32160_, _31341_, _05200_);
  or _82331_ (_32162_, _32160_, _32103_);
  and _82332_ (_32163_, _32162_, _03221_);
  or _82333_ (_32164_, _32163_, _03437_);
  or _82334_ (_32165_, _32164_, _32159_);
  and _82335_ (_32166_, _05200_, _06217_);
  or _82336_ (_32167_, _32166_, _32103_);
  or _82337_ (_32168_, _32167_, _03438_);
  and _82338_ (_32169_, _32168_, _32165_);
  or _82339_ (_32170_, _32169_, _03636_);
  and _82340_ (_32171_, _12598_, _05200_);
  or _82341_ (_32173_, _32171_, _32103_);
  or _82342_ (_32174_, _32173_, _04499_);
  and _82343_ (_32175_, _32174_, _04501_);
  and _82344_ (_32176_, _32175_, _32170_);
  or _82345_ (_32177_, _32176_, _32107_);
  and _82346_ (_32178_, _32177_, _05769_);
  or _82347_ (_32179_, _32103_, _05521_);
  and _82348_ (_32180_, _32179_, _03754_);
  and _82349_ (_32181_, _32180_, _32167_);
  or _82350_ (_32182_, _32181_, _32178_);
  and _82351_ (_32184_, _32182_, _03753_);
  and _82352_ (_32185_, _32115_, _03752_);
  and _82353_ (_32186_, _32185_, _32179_);
  or _82354_ (_32187_, _32186_, _03758_);
  or _82355_ (_32188_, _32187_, _32184_);
  nor _82356_ (_32189_, _12597_, _10989_);
  or _82357_ (_32190_, _32103_, _03759_);
  or _82358_ (_32191_, _32190_, _32189_);
  and _82359_ (_32192_, _32191_, _04517_);
  and _82360_ (_32193_, _32192_, _32188_);
  nor _82361_ (_32195_, _12603_, _10989_);
  or _82362_ (_32196_, _32195_, _32103_);
  and _82363_ (_32197_, _32196_, _03760_);
  or _82364_ (_32198_, _32197_, _03790_);
  or _82365_ (_32199_, _32198_, _32193_);
  or _82366_ (_32200_, _32112_, _04192_);
  and _82367_ (_32201_, _32200_, _03152_);
  and _82368_ (_32202_, _32201_, _32199_);
  and _82369_ (_32203_, _32137_, _03151_);
  or _82370_ (_32204_, _32203_, _03520_);
  or _82371_ (_32206_, _32204_, _32202_);
  and _82372_ (_32207_, _12658_, _05200_);
  or _82373_ (_32208_, _32103_, _03521_);
  or _82374_ (_32209_, _32208_, _32207_);
  and _82375_ (_32210_, _32209_, _42963_);
  and _82376_ (_32211_, _32210_, _32206_);
  nor _82377_ (_32212_, \oc8051_golden_model_1.P3 [3], rst);
  nor _82378_ (_32213_, _32212_, _00000_);
  or _82379_ (_43358_, _32213_, _32211_);
  and _82380_ (_32214_, _10989_, \oc8051_golden_model_1.P3 [4]);
  and _82381_ (_32216_, _12844_, _05200_);
  or _82382_ (_32217_, _32216_, _32214_);
  and _82383_ (_32218_, _32217_, _03769_);
  nor _82384_ (_32219_, _05712_, _10989_);
  or _82385_ (_32220_, _32219_, _32214_);
  or _82386_ (_32221_, _32220_, _06039_);
  nor _82387_ (_32222_, _12733_, _10989_);
  or _82388_ (_32223_, _32222_, _32214_);
  or _82389_ (_32224_, _32223_, _04444_);
  and _82390_ (_32225_, _05200_, \oc8051_golden_model_1.ACC [4]);
  or _82391_ (_32227_, _32225_, _32214_);
  and _82392_ (_32228_, _32227_, _04426_);
  and _82393_ (_32229_, _04427_, \oc8051_golden_model_1.P3 [4]);
  or _82394_ (_32230_, _32229_, _03570_);
  or _82395_ (_32231_, _32230_, _32228_);
  and _82396_ (_32232_, _32231_, _03517_);
  and _82397_ (_32233_, _32232_, _32224_);
  and _82398_ (_32234_, _10997_, \oc8051_golden_model_1.P3 [4]);
  and _82399_ (_32235_, _12737_, _05796_);
  or _82400_ (_32236_, _32235_, _32234_);
  and _82401_ (_32237_, _32236_, _03516_);
  or _82402_ (_32238_, _32237_, _03568_);
  or _82403_ (_32239_, _32238_, _32233_);
  or _82404_ (_32240_, _32220_, _03983_);
  and _82405_ (_32241_, _32240_, _32239_);
  or _82406_ (_32242_, _32241_, _03575_);
  or _82407_ (_32243_, _32227_, _03583_);
  and _82408_ (_32244_, _32243_, _03513_);
  and _82409_ (_32245_, _32244_, _32242_);
  and _82410_ (_32246_, _12718_, _05796_);
  or _82411_ (_32248_, _32246_, _32234_);
  and _82412_ (_32249_, _32248_, _03512_);
  or _82413_ (_32250_, _32249_, _03505_);
  or _82414_ (_32251_, _32250_, _32245_);
  or _82415_ (_32252_, _32234_, _12752_);
  and _82416_ (_32253_, _32252_, _32236_);
  or _82417_ (_32254_, _32253_, _03506_);
  and _82418_ (_32255_, _32254_, _03500_);
  and _82419_ (_32256_, _32255_, _32251_);
  and _82420_ (_32257_, _31439_, _05796_);
  or _82421_ (_32259_, _32257_, _32234_);
  and _82422_ (_32260_, _32259_, _03499_);
  or _82423_ (_32261_, _32260_, _07314_);
  or _82424_ (_32262_, _32261_, _32256_);
  and _82425_ (_32263_, _32262_, _32221_);
  or _82426_ (_32264_, _32263_, _03479_);
  and _82427_ (_32265_, _06722_, _05200_);
  or _82428_ (_32266_, _32214_, _06044_);
  or _82429_ (_32267_, _32266_, _32265_);
  and _82430_ (_32268_, _32267_, _03474_);
  and _82431_ (_32270_, _32268_, _32264_);
  and _82432_ (_32271_, _31468_, _05200_);
  or _82433_ (_32272_, _32271_, _32214_);
  and _82434_ (_32273_, _32272_, _03221_);
  or _82435_ (_32274_, _32273_, _03437_);
  or _82436_ (_32275_, _32274_, _32270_);
  and _82437_ (_32276_, _06233_, _05200_);
  or _82438_ (_32277_, _32276_, _32214_);
  or _82439_ (_32278_, _32277_, _03438_);
  and _82440_ (_32279_, _32278_, _32275_);
  or _82441_ (_32281_, _32279_, _03636_);
  and _82442_ (_32282_, _12711_, _05200_);
  or _82443_ (_32283_, _32282_, _32214_);
  or _82444_ (_32284_, _32283_, _04499_);
  and _82445_ (_32285_, _32284_, _04501_);
  and _82446_ (_32286_, _32285_, _32281_);
  or _82447_ (_32287_, _32286_, _32218_);
  and _82448_ (_32288_, _32287_, _05769_);
  or _82449_ (_32289_, _32214_, _05761_);
  and _82450_ (_32290_, _32289_, _03754_);
  and _82451_ (_32292_, _32290_, _32277_);
  or _82452_ (_32293_, _32292_, _32288_);
  and _82453_ (_32294_, _32293_, _03753_);
  and _82454_ (_32295_, _32227_, _03752_);
  and _82455_ (_32296_, _32295_, _32289_);
  or _82456_ (_32297_, _32296_, _03758_);
  or _82457_ (_32298_, _32297_, _32294_);
  nor _82458_ (_32299_, _12710_, _10989_);
  or _82459_ (_32300_, _32214_, _03759_);
  or _82460_ (_32301_, _32300_, _32299_);
  and _82461_ (_32303_, _32301_, _04517_);
  and _82462_ (_32304_, _32303_, _32298_);
  nor _82463_ (_32305_, _12843_, _10989_);
  or _82464_ (_32306_, _32305_, _32214_);
  and _82465_ (_32307_, _32306_, _03760_);
  or _82466_ (_32308_, _32307_, _03790_);
  or _82467_ (_32309_, _32308_, _32304_);
  or _82468_ (_32310_, _32223_, _04192_);
  and _82469_ (_32311_, _32310_, _03152_);
  and _82470_ (_32312_, _32311_, _32309_);
  and _82471_ (_32314_, _32248_, _03151_);
  or _82472_ (_32315_, _32314_, _03520_);
  or _82473_ (_32316_, _32315_, _32312_);
  and _82474_ (_32317_, _12893_, _05200_);
  or _82475_ (_32318_, _32214_, _03521_);
  or _82476_ (_32319_, _32318_, _32317_);
  and _82477_ (_32320_, _32319_, _42963_);
  and _82478_ (_32321_, _32320_, _32316_);
  nor _82479_ (_32322_, \oc8051_golden_model_1.P3 [4], rst);
  nor _82480_ (_32323_, _32322_, _00000_);
  or _82481_ (_43359_, _32323_, _32321_);
  and _82482_ (_32325_, _10989_, \oc8051_golden_model_1.P3 [5]);
  and _82483_ (_32326_, _13042_, _05200_);
  or _82484_ (_32327_, _32326_, _32325_);
  and _82485_ (_32328_, _32327_, _03769_);
  nor _82486_ (_32329_, _05422_, _10989_);
  or _82487_ (_32330_, _32329_, _32325_);
  or _82488_ (_32331_, _32330_, _06039_);
  nor _82489_ (_32332_, _12930_, _10989_);
  or _82490_ (_32333_, _32332_, _32325_);
  or _82491_ (_32335_, _32333_, _04444_);
  and _82492_ (_32336_, _05200_, \oc8051_golden_model_1.ACC [5]);
  or _82493_ (_32337_, _32336_, _32325_);
  and _82494_ (_32338_, _32337_, _04426_);
  and _82495_ (_32339_, _04427_, \oc8051_golden_model_1.P3 [5]);
  or _82496_ (_32340_, _32339_, _03570_);
  or _82497_ (_32341_, _32340_, _32338_);
  and _82498_ (_32342_, _32341_, _03517_);
  and _82499_ (_32343_, _32342_, _32335_);
  and _82500_ (_32344_, _10997_, \oc8051_golden_model_1.P3 [5]);
  and _82501_ (_32345_, _12934_, _05796_);
  or _82502_ (_32346_, _32345_, _32344_);
  and _82503_ (_32347_, _32346_, _03516_);
  or _82504_ (_32348_, _32347_, _03568_);
  or _82505_ (_32349_, _32348_, _32343_);
  or _82506_ (_32350_, _32330_, _03983_);
  and _82507_ (_32351_, _32350_, _32349_);
  or _82508_ (_32352_, _32351_, _03575_);
  or _82509_ (_32353_, _32337_, _03583_);
  and _82510_ (_32354_, _32353_, _03513_);
  and _82511_ (_32357_, _32354_, _32352_);
  and _82512_ (_32358_, _12914_, _05796_);
  or _82513_ (_32359_, _32358_, _32344_);
  and _82514_ (_32360_, _32359_, _03512_);
  or _82515_ (_32361_, _32360_, _03505_);
  or _82516_ (_32362_, _32361_, _32357_);
  or _82517_ (_32363_, _32344_, _12949_);
  and _82518_ (_32364_, _32363_, _32346_);
  or _82519_ (_32365_, _32364_, _03506_);
  and _82520_ (_32366_, _32365_, _03500_);
  and _82521_ (_32368_, _32366_, _32362_);
  and _82522_ (_32369_, _31567_, _05796_);
  or _82523_ (_32370_, _32369_, _32344_);
  and _82524_ (_32371_, _32370_, _03499_);
  or _82525_ (_32372_, _32371_, _07314_);
  or _82526_ (_32373_, _32372_, _32368_);
  and _82527_ (_32374_, _32373_, _32331_);
  or _82528_ (_32375_, _32374_, _03479_);
  and _82529_ (_32376_, _06721_, _05200_);
  or _82530_ (_32377_, _32325_, _06044_);
  or _82531_ (_32379_, _32377_, _32376_);
  and _82532_ (_32380_, _32379_, _03474_);
  and _82533_ (_32381_, _32380_, _32375_);
  and _82534_ (_32382_, _31593_, _05200_);
  or _82535_ (_32383_, _32382_, _32325_);
  and _82536_ (_32384_, _32383_, _03221_);
  or _82537_ (_32385_, _32384_, _03437_);
  or _82538_ (_32386_, _32385_, _32381_);
  and _82539_ (_32387_, _06211_, _05200_);
  or _82540_ (_32388_, _32387_, _32325_);
  or _82541_ (_32390_, _32388_, _03438_);
  and _82542_ (_32391_, _32390_, _32386_);
  or _82543_ (_32392_, _32391_, _03636_);
  and _82544_ (_32393_, _13036_, _05200_);
  or _82545_ (_32394_, _32393_, _32325_);
  or _82546_ (_32395_, _32394_, _04499_);
  and _82547_ (_32396_, _32395_, _04501_);
  and _82548_ (_32397_, _32396_, _32392_);
  or _82549_ (_32398_, _32397_, _32328_);
  and _82550_ (_32399_, _32398_, _05769_);
  or _82551_ (_32401_, _32325_, _05472_);
  and _82552_ (_32402_, _32401_, _03754_);
  and _82553_ (_32403_, _32402_, _32388_);
  or _82554_ (_32404_, _32403_, _32399_);
  and _82555_ (_32405_, _32404_, _03753_);
  and _82556_ (_32406_, _32337_, _03752_);
  and _82557_ (_32407_, _32406_, _32401_);
  or _82558_ (_32408_, _32407_, _03758_);
  or _82559_ (_32409_, _32408_, _32405_);
  nor _82560_ (_32410_, _13035_, _10989_);
  or _82561_ (_32412_, _32325_, _03759_);
  or _82562_ (_32413_, _32412_, _32410_);
  and _82563_ (_32414_, _32413_, _04517_);
  and _82564_ (_32415_, _32414_, _32409_);
  nor _82565_ (_32416_, _13041_, _10989_);
  or _82566_ (_32417_, _32416_, _32325_);
  and _82567_ (_32418_, _32417_, _03760_);
  or _82568_ (_32419_, _32418_, _03790_);
  or _82569_ (_32420_, _32419_, _32415_);
  or _82570_ (_32421_, _32333_, _04192_);
  and _82571_ (_32423_, _32421_, _03152_);
  and _82572_ (_32424_, _32423_, _32420_);
  and _82573_ (_32425_, _32359_, _03151_);
  or _82574_ (_32426_, _32425_, _03520_);
  or _82575_ (_32427_, _32426_, _32424_);
  and _82576_ (_32428_, _13097_, _05200_);
  or _82577_ (_32429_, _32325_, _03521_);
  or _82578_ (_32430_, _32429_, _32428_);
  and _82579_ (_32431_, _32430_, _42963_);
  and _82580_ (_32432_, _32431_, _32427_);
  nor _82581_ (_32434_, \oc8051_golden_model_1.P3 [5], rst);
  nor _82582_ (_32435_, _32434_, _00000_);
  or _82583_ (_43360_, _32435_, _32432_);
  and _82584_ (_32436_, _10989_, \oc8051_golden_model_1.P3 [6]);
  and _82585_ (_32437_, _13259_, _05200_);
  or _82586_ (_32438_, _32437_, _32436_);
  and _82587_ (_32439_, _32438_, _03769_);
  nor _82588_ (_32440_, _05327_, _10989_);
  or _82589_ (_32441_, _32440_, _32436_);
  or _82590_ (_32442_, _32441_, _06039_);
  nor _82591_ (_32444_, _13122_, _10989_);
  or _82592_ (_32445_, _32444_, _32436_);
  or _82593_ (_32446_, _32445_, _04444_);
  and _82594_ (_32447_, _05200_, \oc8051_golden_model_1.ACC [6]);
  or _82595_ (_32448_, _32447_, _32436_);
  and _82596_ (_32449_, _32448_, _04426_);
  and _82597_ (_32450_, _04427_, \oc8051_golden_model_1.P3 [6]);
  or _82598_ (_32451_, _32450_, _03570_);
  or _82599_ (_32452_, _32451_, _32449_);
  and _82600_ (_32453_, _32452_, _03517_);
  and _82601_ (_32455_, _32453_, _32446_);
  and _82602_ (_32456_, _10997_, \oc8051_golden_model_1.P3 [6]);
  and _82603_ (_32457_, _13145_, _05796_);
  or _82604_ (_32458_, _32457_, _32456_);
  and _82605_ (_32459_, _32458_, _03516_);
  or _82606_ (_32460_, _32459_, _03568_);
  or _82607_ (_32461_, _32460_, _32455_);
  or _82608_ (_32462_, _32441_, _03983_);
  and _82609_ (_32463_, _32462_, _32461_);
  or _82610_ (_32464_, _32463_, _03575_);
  or _82611_ (_32466_, _32448_, _03583_);
  and _82612_ (_32467_, _32466_, _03513_);
  and _82613_ (_32468_, _32467_, _32464_);
  and _82614_ (_32469_, _13130_, _05796_);
  or _82615_ (_32470_, _32469_, _32456_);
  and _82616_ (_32471_, _32470_, _03512_);
  or _82617_ (_32472_, _32471_, _03505_);
  or _82618_ (_32473_, _32472_, _32468_);
  or _82619_ (_32474_, _32456_, _13160_);
  and _82620_ (_32475_, _32474_, _32458_);
  or _82621_ (_32477_, _32475_, _03506_);
  and _82622_ (_32478_, _32477_, _03500_);
  and _82623_ (_32479_, _32478_, _32473_);
  and _82624_ (_32480_, _31693_, _05796_);
  or _82625_ (_32481_, _32480_, _32456_);
  and _82626_ (_32482_, _32481_, _03499_);
  or _82627_ (_32483_, _32482_, _07314_);
  or _82628_ (_32484_, _32483_, _32479_);
  and _82629_ (_32485_, _32484_, _32442_);
  or _82630_ (_32486_, _32485_, _03479_);
  and _82631_ (_32488_, _06713_, _05200_);
  or _82632_ (_32489_, _32436_, _06044_);
  or _82633_ (_32490_, _32489_, _32488_);
  and _82634_ (_32491_, _32490_, _03474_);
  and _82635_ (_32492_, _32491_, _32486_);
  and _82636_ (_32493_, _31718_, _05200_);
  or _82637_ (_32494_, _32493_, _32436_);
  and _82638_ (_32495_, _32494_, _03221_);
  or _82639_ (_32496_, _32495_, _03437_);
  or _82640_ (_32497_, _32496_, _32492_);
  and _82641_ (_32499_, _13244_, _05200_);
  or _82642_ (_32500_, _32499_, _32436_);
  or _82643_ (_32501_, _32500_, _03438_);
  and _82644_ (_32502_, _32501_, _32497_);
  or _82645_ (_32503_, _32502_, _03636_);
  and _82646_ (_32504_, _13253_, _05200_);
  or _82647_ (_32505_, _32504_, _32436_);
  or _82648_ (_32506_, _32505_, _04499_);
  and _82649_ (_32507_, _32506_, _04501_);
  and _82650_ (_32508_, _32507_, _32503_);
  or _82651_ (_32510_, _32508_, _32439_);
  and _82652_ (_32511_, _32510_, _05769_);
  or _82653_ (_32512_, _32436_, _05377_);
  and _82654_ (_32513_, _32512_, _03754_);
  and _82655_ (_32514_, _32513_, _32500_);
  or _82656_ (_32515_, _32514_, _32511_);
  and _82657_ (_32516_, _32515_, _03753_);
  and _82658_ (_32517_, _32448_, _03752_);
  and _82659_ (_32518_, _32517_, _32512_);
  or _82660_ (_32519_, _32518_, _03758_);
  or _82661_ (_32521_, _32519_, _32516_);
  nor _82662_ (_32522_, _13251_, _10989_);
  or _82663_ (_32523_, _32436_, _03759_);
  or _82664_ (_32524_, _32523_, _32522_);
  and _82665_ (_32525_, _32524_, _04517_);
  and _82666_ (_32526_, _32525_, _32521_);
  nor _82667_ (_32527_, _13258_, _10989_);
  or _82668_ (_32528_, _32527_, _32436_);
  and _82669_ (_32529_, _32528_, _03760_);
  or _82670_ (_32530_, _32529_, _03790_);
  or _82671_ (_32532_, _32530_, _32526_);
  or _82672_ (_32533_, _32445_, _04192_);
  and _82673_ (_32534_, _32533_, _03152_);
  and _82674_ (_32535_, _32534_, _32532_);
  and _82675_ (_32536_, _32470_, _03151_);
  or _82676_ (_32537_, _32536_, _03520_);
  or _82677_ (_32538_, _32537_, _32535_);
  and _82678_ (_32539_, _13312_, _05200_);
  or _82679_ (_32540_, _32436_, _03521_);
  or _82680_ (_32541_, _32540_, _32539_);
  and _82681_ (_32543_, _32541_, _42963_);
  and _82682_ (_32544_, _32543_, _32538_);
  nor _82683_ (_32545_, \oc8051_golden_model_1.P3 [6], rst);
  nor _82684_ (_32546_, _32545_, _00000_);
  or _82685_ (_43361_, _32546_, _32544_);
  and _82686_ (_32547_, _11092_, \oc8051_golden_model_1.P0 [0]);
  and _82687_ (_32548_, _11995_, _05276_);
  or _82688_ (_32549_, _32548_, _32547_);
  and _82689_ (_32550_, _32549_, _03769_);
  and _82690_ (_32551_, _05276_, _04419_);
  or _82691_ (_32553_, _32551_, _32547_);
  or _82692_ (_32554_, _32553_, _06039_);
  and _82693_ (_32555_, _05941_, _05276_);
  or _82694_ (_32556_, _32555_, _32547_);
  or _82695_ (_32557_, _32556_, _04444_);
  and _82696_ (_32558_, _05276_, \oc8051_golden_model_1.ACC [0]);
  or _82697_ (_32559_, _32558_, _32547_);
  and _82698_ (_32560_, _32559_, _04426_);
  and _82699_ (_32561_, _04427_, \oc8051_golden_model_1.P0 [0]);
  or _82700_ (_32562_, _32561_, _03570_);
  or _82701_ (_32564_, _32562_, _32560_);
  and _82702_ (_32565_, _32564_, _03517_);
  and _82703_ (_32566_, _32565_, _32557_);
  and _82704_ (_32567_, _11100_, \oc8051_golden_model_1.P0 [0]);
  and _82705_ (_32568_, _11887_, _05205_);
  or _82706_ (_32569_, _32568_, _32567_);
  and _82707_ (_32570_, _32569_, _03516_);
  or _82708_ (_32571_, _32570_, _32566_);
  and _82709_ (_32572_, _32571_, _03983_);
  and _82710_ (_32573_, _32553_, _03568_);
  or _82711_ (_32575_, _32573_, _03575_);
  or _82712_ (_32576_, _32575_, _32572_);
  or _82713_ (_32577_, _32559_, _03583_);
  and _82714_ (_32578_, _32577_, _03513_);
  and _82715_ (_32579_, _32578_, _32576_);
  and _82716_ (_32580_, _32547_, _03512_);
  or _82717_ (_32581_, _32580_, _03505_);
  or _82718_ (_32582_, _32581_, _32579_);
  or _82719_ (_32583_, _32556_, _03506_);
  and _82720_ (_32584_, _32583_, _03500_);
  and _82721_ (_32586_, _32584_, _32582_);
  and _82722_ (_32587_, _30938_, _05205_);
  or _82723_ (_32588_, _32587_, _32567_);
  and _82724_ (_32589_, _32588_, _03499_);
  or _82725_ (_32590_, _32589_, _07314_);
  or _82726_ (_32591_, _32590_, _32586_);
  and _82727_ (_32592_, _32591_, _32554_);
  or _82728_ (_32593_, _32592_, _03479_);
  and _82729_ (_32594_, _06715_, _05276_);
  or _82730_ (_32595_, _32547_, _06044_);
  or _82731_ (_32597_, _32595_, _32594_);
  and _82732_ (_32598_, _32597_, _03474_);
  and _82733_ (_32599_, _32598_, _32593_);
  and _82734_ (_32600_, _30965_, _05276_);
  or _82735_ (_32601_, _32600_, _32547_);
  and _82736_ (_32602_, _32601_, _03221_);
  or _82737_ (_32603_, _32602_, _03437_);
  or _82738_ (_32604_, _32603_, _32599_);
  and _82739_ (_32605_, _05276_, _06202_);
  or _82740_ (_32606_, _32605_, _32547_);
  or _82741_ (_32608_, _32606_, _03438_);
  and _82742_ (_32609_, _32608_, _32604_);
  or _82743_ (_32610_, _32609_, _03636_);
  and _82744_ (_32611_, _11990_, _05276_);
  or _82745_ (_32612_, _32611_, _32547_);
  or _82746_ (_32613_, _32612_, _04499_);
  and _82747_ (_32614_, _32613_, _04501_);
  and _82748_ (_32615_, _32614_, _32610_);
  or _82749_ (_32616_, _32615_, _32550_);
  and _82750_ (_32617_, _32616_, _05769_);
  nand _82751_ (_32619_, _32606_, _03754_);
  nor _82752_ (_32620_, _32619_, _32555_);
  or _82753_ (_32621_, _32620_, _32617_);
  and _82754_ (_32622_, _32621_, _03753_);
  or _82755_ (_32623_, _32547_, _05617_);
  and _82756_ (_32624_, _32559_, _03752_);
  and _82757_ (_32625_, _32624_, _32623_);
  or _82758_ (_32626_, _32625_, _03758_);
  or _82759_ (_32627_, _32626_, _32622_);
  nor _82760_ (_32628_, _11988_, _11092_);
  or _82761_ (_32630_, _32547_, _03759_);
  or _82762_ (_32631_, _32630_, _32628_);
  and _82763_ (_32632_, _32631_, _04517_);
  and _82764_ (_32633_, _32632_, _32627_);
  nor _82765_ (_32634_, _11870_, _11092_);
  or _82766_ (_32635_, _32634_, _32547_);
  and _82767_ (_32636_, _32635_, _03760_);
  or _82768_ (_32637_, _32636_, _03790_);
  or _82769_ (_32638_, _32637_, _32633_);
  or _82770_ (_32639_, _32556_, _04192_);
  and _82771_ (_32641_, _32639_, _03152_);
  and _82772_ (_32642_, _32641_, _32638_);
  and _82773_ (_32643_, _32547_, _03151_);
  or _82774_ (_32644_, _32643_, _03520_);
  or _82775_ (_32645_, _32644_, _32642_);
  or _82776_ (_32646_, _32556_, _03521_);
  and _82777_ (_32647_, _32646_, _42963_);
  and _82778_ (_32648_, _32647_, _32645_);
  nor _82779_ (_32649_, \oc8051_golden_model_1.P0 [0], rst);
  nor _82780_ (_32650_, _32649_, _00000_);
  or _82781_ (_43363_, _32650_, _32648_);
  and _82782_ (_32651_, _11092_, \oc8051_golden_model_1.P0 [1]);
  nor _82783_ (_32652_, _11092_, _04603_);
  or _82784_ (_32653_, _32652_, _32651_);
  and _82785_ (_32654_, _32653_, _03568_);
  and _82786_ (_32655_, _11100_, \oc8051_golden_model_1.P0 [1]);
  and _82787_ (_32656_, _12083_, _05205_);
  or _82788_ (_32657_, _32656_, _32655_);
  or _82789_ (_32658_, _32657_, _03517_);
  or _82790_ (_32659_, _05276_, \oc8051_golden_model_1.P0 [1]);
  and _82791_ (_32662_, _12252_, _05276_);
  not _82792_ (_32663_, _32662_);
  and _82793_ (_32664_, _32663_, _32659_);
  and _82794_ (_32665_, _32664_, _03570_);
  nand _82795_ (_32666_, _05276_, _03233_);
  and _82796_ (_32667_, _32666_, _32659_);
  and _82797_ (_32668_, _32667_, _04426_);
  and _82798_ (_32669_, _04427_, \oc8051_golden_model_1.P0 [1]);
  or _82799_ (_32670_, _32669_, _32668_);
  and _82800_ (_32671_, _32670_, _04444_);
  or _82801_ (_32673_, _32671_, _03516_);
  or _82802_ (_32674_, _32673_, _32665_);
  and _82803_ (_32675_, _32674_, _32658_);
  and _82804_ (_32676_, _32675_, _03983_);
  or _82805_ (_32677_, _32676_, _32654_);
  or _82806_ (_32678_, _32677_, _03575_);
  or _82807_ (_32679_, _32667_, _03583_);
  and _82808_ (_32680_, _32679_, _03513_);
  and _82809_ (_32681_, _32680_, _32678_);
  and _82810_ (_32682_, _12069_, _05205_);
  or _82811_ (_32684_, _32682_, _32655_);
  and _82812_ (_32685_, _32684_, _03512_);
  or _82813_ (_32686_, _32685_, _03505_);
  or _82814_ (_32687_, _32686_, _32681_);
  or _82815_ (_32688_, _32655_, _12098_);
  and _82816_ (_32689_, _32688_, _32657_);
  or _82817_ (_32690_, _32689_, _03506_);
  and _82818_ (_32691_, _32690_, _03500_);
  and _82819_ (_32692_, _32691_, _32687_);
  and _82820_ (_32693_, _31057_, _05205_);
  or _82821_ (_32695_, _32693_, _32655_);
  and _82822_ (_32696_, _32695_, _03499_);
  or _82823_ (_32697_, _32696_, _07314_);
  or _82824_ (_32698_, _32697_, _32692_);
  or _82825_ (_32699_, _32653_, _06039_);
  and _82826_ (_32700_, _32699_, _32698_);
  or _82827_ (_32701_, _32700_, _03479_);
  and _82828_ (_32702_, _06714_, _05276_);
  or _82829_ (_32703_, _32651_, _06044_);
  or _82830_ (_32704_, _32703_, _32702_);
  and _82831_ (_32706_, _32704_, _03474_);
  and _82832_ (_32707_, _32706_, _32701_);
  and _82833_ (_32708_, _31085_, _05276_);
  or _82834_ (_32709_, _32708_, _32651_);
  and _82835_ (_32710_, _32709_, _03221_);
  or _82836_ (_32711_, _32710_, _32707_);
  and _82837_ (_32712_, _32711_, _03438_);
  nand _82838_ (_32713_, _05276_, _04317_);
  and _82839_ (_32714_, _32659_, _03437_);
  and _82840_ (_32715_, _32714_, _32713_);
  or _82841_ (_32717_, _32715_, _32712_);
  and _82842_ (_32718_, _32717_, _04499_);
  or _82843_ (_32719_, _12191_, _11092_);
  and _82844_ (_32720_, _32659_, _03636_);
  and _82845_ (_32721_, _32720_, _32719_);
  or _82846_ (_32722_, _32721_, _32718_);
  and _82847_ (_32723_, _32722_, _04501_);
  or _82848_ (_32724_, _12197_, _11092_);
  and _82849_ (_32725_, _32659_, _03769_);
  and _82850_ (_32726_, _32725_, _32724_);
  or _82851_ (_32728_, _32726_, _32723_);
  and _82852_ (_32729_, _32728_, _05769_);
  or _82853_ (_32730_, _12190_, _11092_);
  and _82854_ (_32731_, _32730_, _03754_);
  and _82855_ (_32732_, _32731_, _32659_);
  or _82856_ (_32733_, _32732_, _32729_);
  and _82857_ (_32734_, _32733_, _03753_);
  or _82858_ (_32735_, _32651_, _05569_);
  and _82859_ (_32736_, _32667_, _03752_);
  and _82860_ (_32737_, _32736_, _32735_);
  or _82861_ (_32739_, _32737_, _32734_);
  and _82862_ (_32740_, _32739_, _03759_);
  or _82863_ (_32741_, _32713_, _05569_);
  and _82864_ (_32742_, _32659_, _03758_);
  and _82865_ (_32743_, _32742_, _32741_);
  or _82866_ (_32744_, _32743_, _32740_);
  and _82867_ (_32745_, _32744_, _04517_);
  nand _82868_ (_32746_, _12196_, _05276_);
  and _82869_ (_32747_, _32746_, _03760_);
  and _82870_ (_32748_, _32747_, _32659_);
  or _82871_ (_32750_, _32748_, _03790_);
  or _82872_ (_32751_, _32750_, _32745_);
  or _82873_ (_32752_, _32664_, _04192_);
  and _82874_ (_32753_, _32752_, _03152_);
  and _82875_ (_32754_, _32753_, _32751_);
  and _82876_ (_32755_, _32684_, _03151_);
  or _82877_ (_32756_, _32755_, _03520_);
  or _82878_ (_32757_, _32756_, _32754_);
  or _82879_ (_32758_, _32651_, _03521_);
  or _82880_ (_32759_, _32758_, _32662_);
  and _82881_ (_32761_, _32759_, _42963_);
  and _82882_ (_32762_, _32761_, _32757_);
  nor _82883_ (_32763_, \oc8051_golden_model_1.P0 [1], rst);
  nor _82884_ (_32764_, _32763_, _00000_);
  or _82885_ (_43364_, _32764_, _32762_);
  and _82886_ (_32765_, _11092_, \oc8051_golden_model_1.P0 [2]);
  and _82887_ (_32766_, _12401_, _05276_);
  or _82888_ (_32767_, _32766_, _32765_);
  and _82889_ (_32768_, _32767_, _03769_);
  nor _82890_ (_32769_, _11092_, _05026_);
  or _82891_ (_32771_, _32769_, _32765_);
  or _82892_ (_32772_, _32771_, _06039_);
  and _82893_ (_32773_, _32771_, _03568_);
  and _82894_ (_32774_, _11100_, \oc8051_golden_model_1.P0 [2]);
  and _82895_ (_32775_, _12278_, _05205_);
  or _82896_ (_32776_, _32775_, _32774_);
  or _82897_ (_32777_, _32776_, _03517_);
  nor _82898_ (_32778_, _12282_, _11092_);
  or _82899_ (_32779_, _32778_, _32765_);
  and _82900_ (_32780_, _32779_, _03570_);
  and _82901_ (_32782_, _04427_, \oc8051_golden_model_1.P0 [2]);
  and _82902_ (_32783_, _05276_, \oc8051_golden_model_1.ACC [2]);
  or _82903_ (_32784_, _32783_, _32765_);
  and _82904_ (_32785_, _32784_, _04426_);
  or _82905_ (_32786_, _32785_, _32782_);
  and _82906_ (_32787_, _32786_, _04444_);
  or _82907_ (_32788_, _32787_, _03516_);
  or _82908_ (_32789_, _32788_, _32780_);
  and _82909_ (_32790_, _32789_, _32777_);
  and _82910_ (_32791_, _32790_, _03983_);
  or _82911_ (_32793_, _32791_, _32773_);
  or _82912_ (_32794_, _32793_, _03575_);
  or _82913_ (_32795_, _32784_, _03583_);
  and _82914_ (_32796_, _32795_, _03513_);
  and _82915_ (_32797_, _32796_, _32794_);
  and _82916_ (_32798_, _12276_, _05205_);
  or _82917_ (_32799_, _32798_, _32774_);
  and _82918_ (_32800_, _32799_, _03512_);
  or _82919_ (_32801_, _32800_, _03505_);
  or _82920_ (_32802_, _32801_, _32797_);
  or _82921_ (_32804_, _32774_, _12309_);
  and _82922_ (_32805_, _32804_, _32776_);
  or _82923_ (_32806_, _32805_, _03506_);
  and _82924_ (_32807_, _32806_, _03500_);
  and _82925_ (_32808_, _32807_, _32802_);
  and _82926_ (_32809_, _31187_, _05205_);
  or _82927_ (_32810_, _32809_, _32774_);
  and _82928_ (_32811_, _32810_, _03499_);
  or _82929_ (_32812_, _32811_, _07314_);
  or _82930_ (_32813_, _32812_, _32808_);
  and _82931_ (_32815_, _32813_, _32772_);
  or _82932_ (_32816_, _32815_, _03479_);
  and _82933_ (_32817_, _06718_, _05276_);
  or _82934_ (_32818_, _32765_, _06044_);
  or _82935_ (_32819_, _32818_, _32817_);
  and _82936_ (_32820_, _32819_, _03474_);
  and _82937_ (_32821_, _32820_, _32816_);
  and _82938_ (_32822_, _31215_, _05276_);
  or _82939_ (_32823_, _32822_, _32765_);
  and _82940_ (_32824_, _32823_, _03221_);
  or _82941_ (_32826_, _32824_, _03437_);
  or _82942_ (_32827_, _32826_, _32821_);
  and _82943_ (_32828_, _05276_, _06261_);
  or _82944_ (_32829_, _32828_, _32765_);
  or _82945_ (_32830_, _32829_, _03438_);
  and _82946_ (_32831_, _32830_, _32827_);
  or _82947_ (_32832_, _32831_, _03636_);
  and _82948_ (_32833_, _12273_, _05276_);
  or _82949_ (_32834_, _32833_, _32765_);
  or _82950_ (_32835_, _32834_, _04499_);
  and _82951_ (_32837_, _32835_, _04501_);
  and _82952_ (_32838_, _32837_, _32832_);
  or _82953_ (_32839_, _32838_, _32768_);
  and _82954_ (_32840_, _32839_, _05769_);
  or _82955_ (_32841_, _32765_, _05665_);
  and _82956_ (_32842_, _32841_, _03754_);
  and _82957_ (_32843_, _32842_, _32829_);
  or _82958_ (_32844_, _32843_, _32840_);
  and _82959_ (_32845_, _32844_, _03753_);
  and _82960_ (_32846_, _32784_, _03752_);
  and _82961_ (_32848_, _32846_, _32841_);
  or _82962_ (_32849_, _32848_, _03758_);
  or _82963_ (_32850_, _32849_, _32845_);
  nor _82964_ (_32851_, _12272_, _11092_);
  or _82965_ (_32852_, _32765_, _03759_);
  or _82966_ (_32853_, _32852_, _32851_);
  and _82967_ (_32854_, _32853_, _04517_);
  and _82968_ (_32855_, _32854_, _32850_);
  nor _82969_ (_32856_, _12400_, _11092_);
  or _82970_ (_32857_, _32856_, _32765_);
  and _82971_ (_32859_, _32857_, _03760_);
  or _82972_ (_32860_, _32859_, _03790_);
  or _82973_ (_32861_, _32860_, _32855_);
  or _82974_ (_32862_, _32779_, _04192_);
  and _82975_ (_32863_, _32862_, _03152_);
  and _82976_ (_32864_, _32863_, _32861_);
  and _82977_ (_32865_, _32799_, _03151_);
  or _82978_ (_32866_, _32865_, _03520_);
  or _82979_ (_32867_, _32866_, _32864_);
  and _82980_ (_32868_, _12456_, _05276_);
  or _82981_ (_32870_, _32765_, _03521_);
  or _82982_ (_32871_, _32870_, _32868_);
  and _82983_ (_32872_, _32871_, _42963_);
  and _82984_ (_32873_, _32872_, _32867_);
  nor _82985_ (_32874_, \oc8051_golden_model_1.P0 [2], rst);
  nor _82986_ (_32875_, _32874_, _00000_);
  or _82987_ (_43365_, _32875_, _32873_);
  and _82988_ (_32876_, _11092_, \oc8051_golden_model_1.P0 [3]);
  and _82989_ (_32877_, _12604_, _05276_);
  or _82990_ (_32878_, _32877_, _32876_);
  and _82991_ (_32880_, _32878_, _03769_);
  nor _82992_ (_32881_, _11092_, _04843_);
  or _82993_ (_32882_, _32881_, _32876_);
  or _82994_ (_32883_, _32882_, _06039_);
  nor _82995_ (_32884_, _12486_, _11092_);
  or _82996_ (_32885_, _32884_, _32876_);
  or _82997_ (_32886_, _32885_, _04444_);
  and _82998_ (_32887_, _05276_, \oc8051_golden_model_1.ACC [3]);
  or _82999_ (_32888_, _32887_, _32876_);
  and _83000_ (_32889_, _32888_, _04426_);
  and _83001_ (_32891_, _04427_, \oc8051_golden_model_1.P0 [3]);
  or _83002_ (_32892_, _32891_, _03570_);
  or _83003_ (_32893_, _32892_, _32889_);
  and _83004_ (_32894_, _32893_, _03517_);
  and _83005_ (_32895_, _32894_, _32886_);
  and _83006_ (_32896_, _11100_, \oc8051_golden_model_1.P0 [3]);
  and _83007_ (_32897_, _12490_, _05205_);
  or _83008_ (_32898_, _32897_, _32896_);
  and _83009_ (_32899_, _32898_, _03516_);
  or _83010_ (_32900_, _32899_, _03568_);
  or _83011_ (_32902_, _32900_, _32895_);
  or _83012_ (_32903_, _32882_, _03983_);
  and _83013_ (_32904_, _32903_, _32902_);
  or _83014_ (_32905_, _32904_, _03575_);
  or _83015_ (_32906_, _32888_, _03583_);
  and _83016_ (_32907_, _32906_, _03513_);
  and _83017_ (_32908_, _32907_, _32905_);
  and _83018_ (_32909_, _12500_, _05205_);
  or _83019_ (_32910_, _32909_, _32896_);
  and _83020_ (_32911_, _32910_, _03512_);
  or _83021_ (_32913_, _32911_, _03505_);
  or _83022_ (_32914_, _32913_, _32908_);
  or _83023_ (_32915_, _32896_, _12507_);
  and _83024_ (_32916_, _32915_, _32898_);
  or _83025_ (_32917_, _32916_, _03506_);
  and _83026_ (_32918_, _32917_, _03500_);
  and _83027_ (_32919_, _32918_, _32914_);
  and _83028_ (_32920_, _31314_, _05205_);
  or _83029_ (_32921_, _32920_, _32896_);
  and _83030_ (_32922_, _32921_, _03499_);
  or _83031_ (_32924_, _32922_, _07314_);
  or _83032_ (_32925_, _32924_, _32919_);
  and _83033_ (_32926_, _32925_, _32883_);
  or _83034_ (_32927_, _32926_, _03479_);
  and _83035_ (_32928_, _06717_, _05276_);
  or _83036_ (_32929_, _32876_, _06044_);
  or _83037_ (_32930_, _32929_, _32928_);
  and _83038_ (_32931_, _32930_, _03474_);
  and _83039_ (_32932_, _32931_, _32927_);
  and _83040_ (_32933_, _31341_, _05276_);
  or _83041_ (_32935_, _32933_, _32876_);
  and _83042_ (_32936_, _32935_, _03221_);
  or _83043_ (_32937_, _32936_, _03437_);
  or _83044_ (_32938_, _32937_, _32932_);
  and _83045_ (_32939_, _05276_, _06217_);
  or _83046_ (_32940_, _32939_, _32876_);
  or _83047_ (_32941_, _32940_, _03438_);
  and _83048_ (_32942_, _32941_, _32938_);
  or _83049_ (_32943_, _32942_, _03636_);
  and _83050_ (_32944_, _12598_, _05276_);
  or _83051_ (_32946_, _32944_, _32876_);
  or _83052_ (_32947_, _32946_, _04499_);
  and _83053_ (_32948_, _32947_, _04501_);
  and _83054_ (_32949_, _32948_, _32943_);
  or _83055_ (_32950_, _32949_, _32880_);
  and _83056_ (_32951_, _32950_, _05769_);
  or _83057_ (_32952_, _32876_, _05521_);
  and _83058_ (_32953_, _32952_, _03754_);
  and _83059_ (_32954_, _32953_, _32940_);
  or _83060_ (_32955_, _32954_, _32951_);
  and _83061_ (_32957_, _32955_, _03753_);
  and _83062_ (_32958_, _32888_, _03752_);
  and _83063_ (_32959_, _32958_, _32952_);
  or _83064_ (_32960_, _32959_, _03758_);
  or _83065_ (_32961_, _32960_, _32957_);
  nor _83066_ (_32962_, _12597_, _11092_);
  or _83067_ (_32963_, _32876_, _03759_);
  or _83068_ (_32964_, _32963_, _32962_);
  and _83069_ (_32965_, _32964_, _04517_);
  and _83070_ (_32966_, _32965_, _32961_);
  nor _83071_ (_32968_, _12603_, _11092_);
  or _83072_ (_32969_, _32968_, _32876_);
  and _83073_ (_32970_, _32969_, _03760_);
  or _83074_ (_32971_, _32970_, _03790_);
  or _83075_ (_32972_, _32971_, _32966_);
  or _83076_ (_32973_, _32885_, _04192_);
  and _83077_ (_32974_, _32973_, _03152_);
  and _83078_ (_32975_, _32974_, _32972_);
  and _83079_ (_32976_, _32910_, _03151_);
  or _83080_ (_32977_, _32976_, _03520_);
  or _83081_ (_32979_, _32977_, _32975_);
  and _83082_ (_32980_, _12658_, _05276_);
  or _83083_ (_32981_, _32876_, _03521_);
  or _83084_ (_32982_, _32981_, _32980_);
  and _83085_ (_32983_, _32982_, _42963_);
  and _83086_ (_32984_, _32983_, _32979_);
  nor _83087_ (_32985_, \oc8051_golden_model_1.P0 [3], rst);
  nor _83088_ (_32986_, _32985_, _00000_);
  or _83089_ (_43366_, _32986_, _32984_);
  and _83090_ (_32987_, _11092_, \oc8051_golden_model_1.P0 [4]);
  and _83091_ (_32988_, _12844_, _05276_);
  or _83092_ (_32989_, _32988_, _32987_);
  and _83093_ (_32990_, _32989_, _03769_);
  nor _83094_ (_32991_, _05712_, _11092_);
  or _83095_ (_32992_, _32991_, _32987_);
  or _83096_ (_32993_, _32992_, _06039_);
  nor _83097_ (_32994_, _12733_, _11092_);
  or _83098_ (_32995_, _32994_, _32987_);
  or _83099_ (_32996_, _32995_, _04444_);
  and _83100_ (_32997_, _05276_, \oc8051_golden_model_1.ACC [4]);
  or _83101_ (_32998_, _32997_, _32987_);
  and _83102_ (_32999_, _32998_, _04426_);
  and _83103_ (_33000_, _04427_, \oc8051_golden_model_1.P0 [4]);
  or _83104_ (_33001_, _33000_, _03570_);
  or _83105_ (_33002_, _33001_, _32999_);
  and _83106_ (_33003_, _33002_, _03517_);
  and _83107_ (_33004_, _33003_, _32996_);
  and _83108_ (_33005_, _11100_, \oc8051_golden_model_1.P0 [4]);
  and _83109_ (_33006_, _12737_, _05205_);
  or _83110_ (_33007_, _33006_, _33005_);
  and _83111_ (_33010_, _33007_, _03516_);
  or _83112_ (_33011_, _33010_, _03568_);
  or _83113_ (_33012_, _33011_, _33004_);
  or _83114_ (_33013_, _32992_, _03983_);
  and _83115_ (_33014_, _33013_, _33012_);
  or _83116_ (_33015_, _33014_, _03575_);
  or _83117_ (_33016_, _32998_, _03583_);
  and _83118_ (_33017_, _33016_, _03513_);
  and _83119_ (_33018_, _33017_, _33015_);
  and _83120_ (_33019_, _12718_, _05205_);
  or _83121_ (_33021_, _33019_, _33005_);
  and _83122_ (_33022_, _33021_, _03512_);
  or _83123_ (_33023_, _33022_, _03505_);
  or _83124_ (_33024_, _33023_, _33018_);
  or _83125_ (_33025_, _33005_, _12752_);
  and _83126_ (_33026_, _33025_, _33007_);
  or _83127_ (_33027_, _33026_, _03506_);
  and _83128_ (_33028_, _33027_, _03500_);
  and _83129_ (_33029_, _33028_, _33024_);
  and _83130_ (_33030_, _31439_, _05205_);
  or _83131_ (_33032_, _33030_, _33005_);
  and _83132_ (_33033_, _33032_, _03499_);
  or _83133_ (_33034_, _33033_, _07314_);
  or _83134_ (_33035_, _33034_, _33029_);
  and _83135_ (_33036_, _33035_, _32993_);
  or _83136_ (_33037_, _33036_, _03479_);
  and _83137_ (_33038_, _06722_, _05276_);
  or _83138_ (_33039_, _32987_, _06044_);
  or _83139_ (_33040_, _33039_, _33038_);
  and _83140_ (_33041_, _33040_, _03474_);
  and _83141_ (_33043_, _33041_, _33037_);
  and _83142_ (_33044_, _31468_, _05276_);
  or _83143_ (_33045_, _33044_, _32987_);
  and _83144_ (_33046_, _33045_, _03221_);
  or _83145_ (_33047_, _33046_, _03437_);
  or _83146_ (_33048_, _33047_, _33043_);
  and _83147_ (_33049_, _06233_, _05276_);
  or _83148_ (_33050_, _33049_, _32987_);
  or _83149_ (_33051_, _33050_, _03438_);
  and _83150_ (_33052_, _33051_, _33048_);
  or _83151_ (_33054_, _33052_, _03636_);
  and _83152_ (_33055_, _12711_, _05276_);
  or _83153_ (_33056_, _33055_, _32987_);
  or _83154_ (_33057_, _33056_, _04499_);
  and _83155_ (_33058_, _33057_, _04501_);
  and _83156_ (_33059_, _33058_, _33054_);
  or _83157_ (_33060_, _33059_, _32990_);
  and _83158_ (_33061_, _33060_, _05769_);
  or _83159_ (_33062_, _32987_, _05761_);
  and _83160_ (_33063_, _33062_, _03754_);
  and _83161_ (_33065_, _33063_, _33050_);
  or _83162_ (_33066_, _33065_, _33061_);
  and _83163_ (_33067_, _33066_, _03753_);
  and _83164_ (_33068_, _32998_, _03752_);
  and _83165_ (_33069_, _33068_, _33062_);
  or _83166_ (_33070_, _33069_, _03758_);
  or _83167_ (_33071_, _33070_, _33067_);
  nor _83168_ (_33072_, _12710_, _11092_);
  or _83169_ (_33073_, _32987_, _03759_);
  or _83170_ (_33074_, _33073_, _33072_);
  and _83171_ (_33076_, _33074_, _04517_);
  and _83172_ (_33077_, _33076_, _33071_);
  nor _83173_ (_33078_, _12843_, _11092_);
  or _83174_ (_33079_, _33078_, _32987_);
  and _83175_ (_33080_, _33079_, _03760_);
  or _83176_ (_33081_, _33080_, _03790_);
  or _83177_ (_33082_, _33081_, _33077_);
  or _83178_ (_33083_, _32995_, _04192_);
  and _83179_ (_33084_, _33083_, _03152_);
  and _83180_ (_33085_, _33084_, _33082_);
  and _83181_ (_33087_, _33021_, _03151_);
  or _83182_ (_33088_, _33087_, _03520_);
  or _83183_ (_33089_, _33088_, _33085_);
  and _83184_ (_33090_, _12893_, _05276_);
  or _83185_ (_33091_, _32987_, _03521_);
  or _83186_ (_33092_, _33091_, _33090_);
  and _83187_ (_33093_, _33092_, _42963_);
  and _83188_ (_33094_, _33093_, _33089_);
  nor _83189_ (_33095_, \oc8051_golden_model_1.P0 [4], rst);
  nor _83190_ (_33096_, _33095_, _00000_);
  or _83191_ (_43367_, _33096_, _33094_);
  not _83192_ (_33098_, \oc8051_golden_model_1.P0 [5]);
  nor _83193_ (_33099_, _42963_, _33098_);
  or _83194_ (_33100_, _33099_, rst);
  nor _83195_ (_33101_, _05276_, _33098_);
  and _83196_ (_33102_, _13042_, _05276_);
  or _83197_ (_33103_, _33102_, _33101_);
  and _83198_ (_33104_, _33103_, _03769_);
  nor _83199_ (_33105_, _05422_, _11092_);
  or _83200_ (_33106_, _33105_, _33101_);
  or _83201_ (_33108_, _33106_, _06039_);
  nor _83202_ (_33109_, _12930_, _11092_);
  or _83203_ (_33110_, _33109_, _33101_);
  or _83204_ (_33111_, _33110_, _04444_);
  and _83205_ (_33112_, _05276_, \oc8051_golden_model_1.ACC [5]);
  or _83206_ (_33113_, _33112_, _33101_);
  and _83207_ (_33114_, _33113_, _04426_);
  nor _83208_ (_33115_, _04426_, _33098_);
  or _83209_ (_33116_, _33115_, _03570_);
  or _83210_ (_33117_, _33116_, _33114_);
  and _83211_ (_33119_, _33117_, _03517_);
  and _83212_ (_33120_, _33119_, _33111_);
  nor _83213_ (_33121_, _05205_, _33098_);
  and _83214_ (_33122_, _12934_, _05205_);
  or _83215_ (_33123_, _33122_, _33121_);
  and _83216_ (_33124_, _33123_, _03516_);
  or _83217_ (_33125_, _33124_, _03568_);
  or _83218_ (_33126_, _33125_, _33120_);
  or _83219_ (_33127_, _33106_, _03983_);
  and _83220_ (_33128_, _33127_, _33126_);
  or _83221_ (_33130_, _33128_, _03575_);
  or _83222_ (_33131_, _33113_, _03583_);
  and _83223_ (_33132_, _33131_, _03513_);
  and _83224_ (_33133_, _33132_, _33130_);
  and _83225_ (_33134_, _12914_, _05205_);
  or _83226_ (_33135_, _33134_, _33121_);
  and _83227_ (_33136_, _33135_, _03512_);
  or _83228_ (_33137_, _33136_, _03505_);
  or _83229_ (_33138_, _33137_, _33133_);
  or _83230_ (_33139_, _33121_, _12949_);
  and _83231_ (_33141_, _33139_, _33123_);
  or _83232_ (_33142_, _33141_, _03506_);
  and _83233_ (_33143_, _33142_, _03500_);
  and _83234_ (_33144_, _33143_, _33138_);
  and _83235_ (_33145_, _31567_, _05205_);
  or _83236_ (_33146_, _33145_, _33121_);
  and _83237_ (_33147_, _33146_, _03499_);
  or _83238_ (_33148_, _33147_, _07314_);
  or _83239_ (_33149_, _33148_, _33144_);
  and _83240_ (_33150_, _33149_, _33108_);
  or _83241_ (_33152_, _33150_, _03479_);
  and _83242_ (_33153_, _06721_, _05276_);
  or _83243_ (_33154_, _33101_, _06044_);
  or _83244_ (_33155_, _33154_, _33153_);
  and _83245_ (_33156_, _33155_, _03474_);
  and _83246_ (_33157_, _33156_, _33152_);
  and _83247_ (_33158_, _31593_, _05276_);
  or _83248_ (_33159_, _33158_, _33101_);
  and _83249_ (_33160_, _33159_, _03221_);
  or _83250_ (_33161_, _33160_, _03437_);
  or _83251_ (_33163_, _33161_, _33157_);
  and _83252_ (_33164_, _06211_, _05276_);
  or _83253_ (_33165_, _33164_, _33101_);
  or _83254_ (_33166_, _33165_, _03438_);
  and _83255_ (_33167_, _33166_, _33163_);
  or _83256_ (_33168_, _33167_, _03636_);
  and _83257_ (_33169_, _13036_, _05276_);
  or _83258_ (_33170_, _33169_, _33101_);
  or _83259_ (_33171_, _33170_, _04499_);
  and _83260_ (_33172_, _33171_, _04501_);
  and _83261_ (_33174_, _33172_, _33168_);
  or _83262_ (_33175_, _33174_, _33104_);
  and _83263_ (_33176_, _33175_, _05769_);
  or _83264_ (_33177_, _33101_, _05472_);
  and _83265_ (_33178_, _33177_, _03754_);
  and _83266_ (_33179_, _33178_, _33165_);
  or _83267_ (_33180_, _33179_, _33176_);
  and _83268_ (_33181_, _33180_, _03753_);
  and _83269_ (_33182_, _33113_, _03752_);
  and _83270_ (_33183_, _33182_, _33177_);
  or _83271_ (_33185_, _33183_, _03758_);
  or _83272_ (_33186_, _33185_, _33181_);
  nor _83273_ (_33187_, _13035_, _11092_);
  or _83274_ (_33188_, _33101_, _03759_);
  or _83275_ (_33189_, _33188_, _33187_);
  and _83276_ (_33190_, _33189_, _04517_);
  and _83277_ (_33191_, _33190_, _33186_);
  nor _83278_ (_33192_, _13041_, _11092_);
  or _83279_ (_33193_, _33192_, _33101_);
  and _83280_ (_33194_, _33193_, _03760_);
  or _83281_ (_33196_, _33194_, _03790_);
  or _83282_ (_33197_, _33196_, _33191_);
  or _83283_ (_33198_, _33110_, _04192_);
  and _83284_ (_33199_, _33198_, _03152_);
  and _83285_ (_33200_, _33199_, _33197_);
  and _83286_ (_33201_, _33135_, _03151_);
  or _83287_ (_33202_, _33201_, _03520_);
  or _83288_ (_33203_, _33202_, _33200_);
  and _83289_ (_33204_, _13097_, _05276_);
  or _83290_ (_33205_, _33101_, _03521_);
  or _83291_ (_33207_, _33205_, _33204_);
  and _83292_ (_33208_, _33207_, _42963_);
  and _83293_ (_33209_, _33208_, _33203_);
  or _83294_ (_43369_, _33209_, _33100_);
  and _83295_ (_33210_, _11092_, \oc8051_golden_model_1.P0 [6]);
  and _83296_ (_33211_, _13259_, _05276_);
  or _83297_ (_33212_, _33211_, _33210_);
  and _83298_ (_33213_, _33212_, _03769_);
  nor _83299_ (_33214_, _05327_, _11092_);
  or _83300_ (_33215_, _33214_, _33210_);
  or _83301_ (_33217_, _33215_, _06039_);
  nor _83302_ (_33218_, _13122_, _11092_);
  or _83303_ (_33219_, _33218_, _33210_);
  or _83304_ (_33220_, _33219_, _04444_);
  and _83305_ (_33221_, _05276_, \oc8051_golden_model_1.ACC [6]);
  or _83306_ (_33222_, _33221_, _33210_);
  and _83307_ (_33223_, _33222_, _04426_);
  and _83308_ (_33224_, _04427_, \oc8051_golden_model_1.P0 [6]);
  or _83309_ (_33225_, _33224_, _03570_);
  or _83310_ (_33226_, _33225_, _33223_);
  and _83311_ (_33228_, _33226_, _03517_);
  and _83312_ (_33229_, _33228_, _33220_);
  and _83313_ (_33230_, _11100_, \oc8051_golden_model_1.P0 [6]);
  and _83314_ (_33231_, _13145_, _05205_);
  or _83315_ (_33232_, _33231_, _33230_);
  and _83316_ (_33233_, _33232_, _03516_);
  or _83317_ (_33234_, _33233_, _03568_);
  or _83318_ (_33235_, _33234_, _33229_);
  or _83319_ (_33236_, _33215_, _03983_);
  and _83320_ (_33237_, _33236_, _33235_);
  or _83321_ (_33239_, _33237_, _03575_);
  or _83322_ (_33240_, _33222_, _03583_);
  and _83323_ (_33241_, _33240_, _03513_);
  and _83324_ (_33242_, _33241_, _33239_);
  and _83325_ (_33243_, _13130_, _05205_);
  or _83326_ (_33244_, _33243_, _33230_);
  and _83327_ (_33245_, _33244_, _03512_);
  or _83328_ (_33246_, _33245_, _03505_);
  or _83329_ (_33247_, _33246_, _33242_);
  or _83330_ (_33248_, _33230_, _13160_);
  and _83331_ (_33250_, _33248_, _33232_);
  or _83332_ (_33251_, _33250_, _03506_);
  and _83333_ (_33252_, _33251_, _03500_);
  and _83334_ (_33253_, _33252_, _33247_);
  and _83335_ (_33254_, _31693_, _05205_);
  or _83336_ (_33255_, _33254_, _33230_);
  and _83337_ (_33256_, _33255_, _03499_);
  or _83338_ (_33257_, _33256_, _07314_);
  or _83339_ (_33258_, _33257_, _33253_);
  and _83340_ (_33259_, _33258_, _33217_);
  or _83341_ (_33261_, _33259_, _03479_);
  and _83342_ (_33262_, _06713_, _05276_);
  or _83343_ (_33263_, _33210_, _06044_);
  or _83344_ (_33264_, _33263_, _33262_);
  and _83345_ (_33265_, _33264_, _03474_);
  and _83346_ (_33266_, _33265_, _33261_);
  and _83347_ (_33267_, _31718_, _05276_);
  or _83348_ (_33268_, _33267_, _33210_);
  and _83349_ (_33269_, _33268_, _03221_);
  or _83350_ (_33270_, _33269_, _03437_);
  or _83351_ (_33272_, _33270_, _33266_);
  and _83352_ (_33273_, _13244_, _05276_);
  or _83353_ (_33274_, _33273_, _33210_);
  or _83354_ (_33275_, _33274_, _03438_);
  and _83355_ (_33276_, _33275_, _33272_);
  or _83356_ (_33277_, _33276_, _03636_);
  and _83357_ (_33278_, _13253_, _05276_);
  or _83358_ (_33279_, _33278_, _33210_);
  or _83359_ (_33280_, _33279_, _04499_);
  and _83360_ (_33281_, _33280_, _04501_);
  and _83361_ (_33283_, _33281_, _33277_);
  or _83362_ (_33284_, _33283_, _33213_);
  and _83363_ (_33285_, _33284_, _05769_);
  or _83364_ (_33286_, _33210_, _05377_);
  and _83365_ (_33287_, _33286_, _03754_);
  and _83366_ (_33288_, _33287_, _33274_);
  or _83367_ (_33289_, _33288_, _33285_);
  and _83368_ (_33290_, _33289_, _03753_);
  and _83369_ (_33291_, _33222_, _03752_);
  and _83370_ (_33292_, _33291_, _33286_);
  or _83371_ (_33294_, _33292_, _03758_);
  or _83372_ (_33295_, _33294_, _33290_);
  nor _83373_ (_33296_, _13251_, _11092_);
  or _83374_ (_33297_, _33210_, _03759_);
  or _83375_ (_33298_, _33297_, _33296_);
  and _83376_ (_33299_, _33298_, _04517_);
  and _83377_ (_33300_, _33299_, _33295_);
  nor _83378_ (_33301_, _13258_, _11092_);
  or _83379_ (_33302_, _33301_, _33210_);
  and _83380_ (_33303_, _33302_, _03760_);
  or _83381_ (_33305_, _33303_, _03790_);
  or _83382_ (_33306_, _33305_, _33300_);
  or _83383_ (_33307_, _33219_, _04192_);
  and _83384_ (_33308_, _33307_, _03152_);
  and _83385_ (_33309_, _33308_, _33306_);
  and _83386_ (_33310_, _33244_, _03151_);
  or _83387_ (_33311_, _33310_, _03520_);
  or _83388_ (_33312_, _33311_, _33309_);
  and _83389_ (_33313_, _13312_, _05276_);
  or _83390_ (_33314_, _33210_, _03521_);
  or _83391_ (_33316_, _33314_, _33313_);
  and _83392_ (_33317_, _33316_, _42963_);
  and _83393_ (_33318_, _33317_, _33312_);
  nor _83394_ (_33319_, \oc8051_golden_model_1.P0 [6], rst);
  nor _83395_ (_33320_, _33319_, _00000_);
  or _83396_ (_43370_, _33320_, _33318_);
  nor _83397_ (_33321_, \oc8051_golden_model_1.P1 [0], rst);
  nor _83398_ (_33322_, _33321_, _00000_);
  and _83399_ (_33323_, _11197_, \oc8051_golden_model_1.P1 [0]);
  and _83400_ (_33324_, _11995_, _05244_);
  or _83401_ (_33326_, _33324_, _33323_);
  and _83402_ (_33327_, _33326_, _03769_);
  and _83403_ (_33328_, _05941_, _05244_);
  or _83404_ (_33329_, _33328_, _33323_);
  and _83405_ (_33330_, _33329_, _03570_);
  and _83406_ (_33331_, _04427_, \oc8051_golden_model_1.P1 [0]);
  and _83407_ (_33332_, _05244_, \oc8051_golden_model_1.ACC [0]);
  or _83408_ (_33333_, _33332_, _33323_);
  and _83409_ (_33334_, _33333_, _04426_);
  or _83410_ (_33335_, _33334_, _33331_);
  and _83411_ (_33337_, _33335_, _04444_);
  or _83412_ (_33338_, _33337_, _03516_);
  or _83413_ (_33339_, _33338_, _33330_);
  and _83414_ (_33340_, _11887_, _05811_);
  and _83415_ (_33341_, _11205_, \oc8051_golden_model_1.P1 [0]);
  or _83416_ (_33342_, _33341_, _03517_);
  or _83417_ (_33343_, _33342_, _33340_);
  and _83418_ (_33344_, _33343_, _03983_);
  and _83419_ (_33345_, _33344_, _33339_);
  and _83420_ (_33346_, _05244_, _04419_);
  or _83421_ (_33348_, _33346_, _33323_);
  and _83422_ (_33349_, _33348_, _03568_);
  or _83423_ (_33350_, _33349_, _03575_);
  or _83424_ (_33351_, _33350_, _33345_);
  or _83425_ (_33352_, _33333_, _03583_);
  and _83426_ (_33353_, _33352_, _03513_);
  and _83427_ (_33354_, _33353_, _33351_);
  and _83428_ (_33355_, _33323_, _03512_);
  or _83429_ (_33356_, _33355_, _03505_);
  or _83430_ (_33357_, _33356_, _33354_);
  or _83431_ (_33359_, _33329_, _03506_);
  and _83432_ (_33360_, _33359_, _03500_);
  and _83433_ (_33361_, _33360_, _33357_);
  and _83434_ (_33362_, _30938_, _05811_);
  or _83435_ (_33363_, _33362_, _33341_);
  and _83436_ (_33364_, _33363_, _03499_);
  or _83437_ (_33365_, _33364_, _07314_);
  or _83438_ (_33366_, _33365_, _33361_);
  or _83439_ (_33367_, _33348_, _06039_);
  and _83440_ (_33368_, _33367_, _33366_);
  or _83441_ (_33369_, _33368_, _03479_);
  and _83442_ (_33370_, _06715_, _05244_);
  or _83443_ (_33371_, _33323_, _06044_);
  or _83444_ (_33372_, _33371_, _33370_);
  and _83445_ (_33373_, _33372_, _03474_);
  and _83446_ (_33374_, _33373_, _33369_);
  and _83447_ (_33375_, _30965_, _05244_);
  or _83448_ (_33376_, _33375_, _33323_);
  and _83449_ (_33377_, _33376_, _03221_);
  or _83450_ (_33378_, _33377_, _03437_);
  or _83451_ (_33381_, _33378_, _33374_);
  and _83452_ (_33382_, _05244_, _06202_);
  or _83453_ (_33383_, _33382_, _33323_);
  or _83454_ (_33384_, _33383_, _03438_);
  and _83455_ (_33385_, _33384_, _33381_);
  or _83456_ (_33386_, _33385_, _03636_);
  and _83457_ (_33387_, _11990_, _05244_);
  or _83458_ (_33388_, _33387_, _33323_);
  or _83459_ (_33389_, _33388_, _04499_);
  and _83460_ (_33390_, _33389_, _04501_);
  and _83461_ (_33392_, _33390_, _33386_);
  or _83462_ (_33393_, _33392_, _33327_);
  and _83463_ (_33394_, _33393_, _05769_);
  nand _83464_ (_33395_, _33383_, _03754_);
  nor _83465_ (_33396_, _33395_, _33328_);
  or _83466_ (_33397_, _33396_, _33394_);
  and _83467_ (_33398_, _33397_, _03753_);
  or _83468_ (_33399_, _33323_, _05617_);
  and _83469_ (_33400_, _33333_, _03752_);
  and _83470_ (_33401_, _33400_, _33399_);
  or _83471_ (_33403_, _33401_, _03758_);
  or _83472_ (_33404_, _33403_, _33398_);
  nor _83473_ (_33405_, _11988_, _11197_);
  or _83474_ (_33406_, _33323_, _03759_);
  or _83475_ (_33407_, _33406_, _33405_);
  and _83476_ (_33408_, _33407_, _04517_);
  and _83477_ (_33409_, _33408_, _33404_);
  nor _83478_ (_33410_, _11870_, _11197_);
  or _83479_ (_33411_, _33410_, _33323_);
  and _83480_ (_33412_, _33411_, _03760_);
  or _83481_ (_33414_, _33412_, _03790_);
  or _83482_ (_33415_, _33414_, _33409_);
  or _83483_ (_33416_, _33329_, _04192_);
  and _83484_ (_33417_, _33416_, _03152_);
  and _83485_ (_33418_, _33417_, _33415_);
  and _83486_ (_33419_, _33323_, _03151_);
  or _83487_ (_33420_, _33419_, _03520_);
  or _83488_ (_33421_, _33420_, _33418_);
  or _83489_ (_33422_, _33329_, _03521_);
  and _83490_ (_33423_, _33422_, _42963_);
  and _83491_ (_33425_, _33423_, _33421_);
  or _83492_ (_43371_, _33425_, _33322_);
  or _83493_ (_33426_, _05244_, \oc8051_golden_model_1.P1 [1]);
  and _83494_ (_33427_, _12252_, _05244_);
  not _83495_ (_33428_, _33427_);
  and _83496_ (_33429_, _33428_, _33426_);
  or _83497_ (_33430_, _33429_, _04444_);
  nand _83498_ (_33431_, _05244_, _03233_);
  and _83499_ (_33432_, _33431_, _33426_);
  and _83500_ (_33433_, _33432_, _04426_);
  and _83501_ (_33435_, _04427_, \oc8051_golden_model_1.P1 [1]);
  or _83502_ (_33436_, _33435_, _03570_);
  or _83503_ (_33437_, _33436_, _33433_);
  and _83504_ (_33438_, _33437_, _03517_);
  and _83505_ (_33439_, _33438_, _33430_);
  and _83506_ (_33440_, _12083_, _05811_);
  and _83507_ (_33441_, _11205_, \oc8051_golden_model_1.P1 [1]);
  or _83508_ (_33442_, _33441_, _03568_);
  or _83509_ (_33443_, _33442_, _33440_);
  and _83510_ (_33444_, _33443_, _14165_);
  or _83511_ (_33446_, _33444_, _33439_);
  and _83512_ (_33447_, _11197_, \oc8051_golden_model_1.P1 [1]);
  nor _83513_ (_33448_, _11197_, _04603_);
  or _83514_ (_33449_, _33448_, _33447_);
  or _83515_ (_33450_, _33449_, _03983_);
  and _83516_ (_33451_, _33450_, _33446_);
  or _83517_ (_33452_, _33451_, _03575_);
  or _83518_ (_33453_, _33432_, _03583_);
  and _83519_ (_33454_, _33453_, _03513_);
  and _83520_ (_33455_, _33454_, _33452_);
  and _83521_ (_33457_, _12069_, _05811_);
  or _83522_ (_33458_, _33457_, _33441_);
  and _83523_ (_33459_, _33458_, _03512_);
  or _83524_ (_33460_, _33459_, _03505_);
  or _83525_ (_33461_, _33460_, _33455_);
  and _83526_ (_33462_, _33440_, _12098_);
  or _83527_ (_33463_, _33441_, _03506_);
  or _83528_ (_33464_, _33463_, _33462_);
  and _83529_ (_33465_, _33464_, _33461_);
  and _83530_ (_33466_, _33465_, _03500_);
  and _83531_ (_33468_, _31057_, _05811_);
  or _83532_ (_33469_, _33441_, _33468_);
  and _83533_ (_33470_, _33469_, _03499_);
  or _83534_ (_33471_, _33470_, _07314_);
  or _83535_ (_33472_, _33471_, _33466_);
  or _83536_ (_33473_, _33449_, _06039_);
  and _83537_ (_33474_, _33473_, _33472_);
  or _83538_ (_33475_, _33474_, _03479_);
  and _83539_ (_33476_, _06714_, _05244_);
  or _83540_ (_33477_, _33447_, _06044_);
  or _83541_ (_33479_, _33477_, _33476_);
  and _83542_ (_33480_, _33479_, _03474_);
  and _83543_ (_33481_, _33480_, _33475_);
  and _83544_ (_33482_, _31085_, _05244_);
  or _83545_ (_33483_, _33482_, _33447_);
  and _83546_ (_33484_, _33483_, _03221_);
  or _83547_ (_33485_, _33484_, _33481_);
  and _83548_ (_33486_, _33485_, _03438_);
  nand _83549_ (_33487_, _05244_, _04317_);
  and _83550_ (_33488_, _33426_, _03437_);
  and _83551_ (_33490_, _33488_, _33487_);
  or _83552_ (_33491_, _33490_, _33486_);
  and _83553_ (_33492_, _33491_, _04499_);
  or _83554_ (_33493_, _12191_, _11197_);
  and _83555_ (_33494_, _33426_, _03636_);
  and _83556_ (_33495_, _33494_, _33493_);
  or _83557_ (_33496_, _33495_, _33492_);
  and _83558_ (_33497_, _33496_, _04501_);
  or _83559_ (_33498_, _12197_, _11197_);
  and _83560_ (_33499_, _33426_, _03769_);
  and _83561_ (_33501_, _33499_, _33498_);
  or _83562_ (_33502_, _33501_, _33497_);
  and _83563_ (_33503_, _33502_, _05769_);
  or _83564_ (_33504_, _12190_, _11197_);
  and _83565_ (_33505_, _33504_, _03754_);
  and _83566_ (_33506_, _33505_, _33426_);
  or _83567_ (_33507_, _33506_, _33503_);
  and _83568_ (_33508_, _33507_, _03753_);
  or _83569_ (_33509_, _33447_, _05569_);
  and _83570_ (_33510_, _33432_, _03752_);
  and _83571_ (_33512_, _33510_, _33509_);
  or _83572_ (_33513_, _33512_, _33508_);
  and _83573_ (_33514_, _33513_, _03759_);
  or _83574_ (_33515_, _33487_, _05569_);
  and _83575_ (_33516_, _33426_, _03758_);
  and _83576_ (_33517_, _33516_, _33515_);
  or _83577_ (_33518_, _33517_, _33514_);
  and _83578_ (_33519_, _33518_, _04517_);
  nand _83579_ (_33520_, _12196_, _05244_);
  and _83580_ (_33521_, _33520_, _03760_);
  and _83581_ (_33523_, _33521_, _33426_);
  or _83582_ (_33524_, _33523_, _03790_);
  or _83583_ (_33525_, _33524_, _33519_);
  or _83584_ (_33526_, _33429_, _04192_);
  and _83585_ (_33527_, _33526_, _03152_);
  and _83586_ (_33528_, _33527_, _33525_);
  and _83587_ (_33529_, _33458_, _03151_);
  or _83588_ (_33530_, _33529_, _03520_);
  or _83589_ (_33531_, _33530_, _33528_);
  or _83590_ (_33532_, _33447_, _03521_);
  or _83591_ (_33534_, _33532_, _33427_);
  and _83592_ (_33535_, _33534_, _42963_);
  and _83593_ (_33536_, _33535_, _33531_);
  nor _83594_ (_33537_, \oc8051_golden_model_1.P1 [1], rst);
  nor _83595_ (_33538_, _33537_, _00000_);
  or _83596_ (_43373_, _33538_, _33536_);
  and _83597_ (_33539_, _11197_, \oc8051_golden_model_1.P1 [2]);
  and _83598_ (_33540_, _12401_, _05244_);
  or _83599_ (_33541_, _33540_, _33539_);
  and _83600_ (_33542_, _33541_, _03769_);
  nor _83601_ (_33544_, _11197_, _05026_);
  or _83602_ (_33545_, _33544_, _33539_);
  or _83603_ (_33546_, _33545_, _06039_);
  or _83604_ (_33547_, _33545_, _03983_);
  nor _83605_ (_33548_, _12282_, _11197_);
  or _83606_ (_33549_, _33548_, _33539_);
  or _83607_ (_33550_, _33549_, _04444_);
  and _83608_ (_33551_, _05244_, \oc8051_golden_model_1.ACC [2]);
  or _83609_ (_33552_, _33551_, _33539_);
  and _83610_ (_33553_, _33552_, _04426_);
  and _83611_ (_33555_, _04427_, \oc8051_golden_model_1.P1 [2]);
  or _83612_ (_33556_, _33555_, _03570_);
  or _83613_ (_33557_, _33556_, _33553_);
  and _83614_ (_33558_, _33557_, _03517_);
  and _83615_ (_33559_, _33558_, _33550_);
  and _83616_ (_33560_, _11205_, \oc8051_golden_model_1.P1 [2]);
  and _83617_ (_33561_, _12278_, _05811_);
  or _83618_ (_33562_, _33561_, _33560_);
  and _83619_ (_33563_, _33562_, _03516_);
  or _83620_ (_33564_, _33563_, _03568_);
  or _83621_ (_33566_, _33564_, _33559_);
  and _83622_ (_33567_, _33566_, _33547_);
  or _83623_ (_33568_, _33567_, _03575_);
  or _83624_ (_33569_, _33552_, _03583_);
  and _83625_ (_33570_, _33569_, _03513_);
  and _83626_ (_33571_, _33570_, _33568_);
  and _83627_ (_33572_, _12276_, _05811_);
  or _83628_ (_33573_, _33572_, _33560_);
  and _83629_ (_33574_, _33573_, _03512_);
  or _83630_ (_33575_, _33574_, _03505_);
  or _83631_ (_33577_, _33575_, _33571_);
  and _83632_ (_33578_, _33561_, _12309_);
  or _83633_ (_33579_, _33560_, _03506_);
  or _83634_ (_33580_, _33579_, _33578_);
  and _83635_ (_33581_, _33580_, _03500_);
  and _83636_ (_33582_, _33581_, _33577_);
  and _83637_ (_33583_, _31187_, _05811_);
  or _83638_ (_33584_, _33583_, _33560_);
  and _83639_ (_33585_, _33584_, _03499_);
  or _83640_ (_33586_, _33585_, _07314_);
  or _83641_ (_33588_, _33586_, _33582_);
  and _83642_ (_33589_, _33588_, _33546_);
  or _83643_ (_33590_, _33589_, _03479_);
  and _83644_ (_33591_, _06718_, _05244_);
  or _83645_ (_33592_, _33539_, _06044_);
  or _83646_ (_33593_, _33592_, _33591_);
  and _83647_ (_33594_, _33593_, _03474_);
  and _83648_ (_33595_, _33594_, _33590_);
  and _83649_ (_33596_, _31215_, _05244_);
  or _83650_ (_33597_, _33596_, _33539_);
  and _83651_ (_33599_, _33597_, _03221_);
  or _83652_ (_33600_, _33599_, _03437_);
  or _83653_ (_33601_, _33600_, _33595_);
  and _83654_ (_33602_, _05244_, _06261_);
  or _83655_ (_33603_, _33602_, _33539_);
  or _83656_ (_33604_, _33603_, _03438_);
  and _83657_ (_33605_, _33604_, _33601_);
  or _83658_ (_33606_, _33605_, _03636_);
  and _83659_ (_33607_, _12273_, _05244_);
  or _83660_ (_33608_, _33607_, _33539_);
  or _83661_ (_33610_, _33608_, _04499_);
  and _83662_ (_33611_, _33610_, _04501_);
  and _83663_ (_33612_, _33611_, _33606_);
  or _83664_ (_33613_, _33612_, _33542_);
  and _83665_ (_33614_, _33613_, _05769_);
  or _83666_ (_33615_, _33539_, _05665_);
  and _83667_ (_33616_, _33615_, _03754_);
  and _83668_ (_33617_, _33616_, _33603_);
  or _83669_ (_33618_, _33617_, _33614_);
  and _83670_ (_33619_, _33618_, _03753_);
  and _83671_ (_33621_, _33552_, _03752_);
  and _83672_ (_33622_, _33621_, _33615_);
  or _83673_ (_33623_, _33622_, _03758_);
  or _83674_ (_33624_, _33623_, _33619_);
  nor _83675_ (_33625_, _12272_, _11197_);
  or _83676_ (_33626_, _33539_, _03759_);
  or _83677_ (_33627_, _33626_, _33625_);
  and _83678_ (_33628_, _33627_, _04517_);
  and _83679_ (_33629_, _33628_, _33624_);
  nor _83680_ (_33630_, _12400_, _11197_);
  or _83681_ (_33632_, _33630_, _33539_);
  and _83682_ (_33633_, _33632_, _03760_);
  or _83683_ (_33634_, _33633_, _03790_);
  or _83684_ (_33635_, _33634_, _33629_);
  or _83685_ (_33636_, _33549_, _04192_);
  and _83686_ (_33637_, _33636_, _03152_);
  and _83687_ (_33638_, _33637_, _33635_);
  and _83688_ (_33639_, _33573_, _03151_);
  or _83689_ (_33640_, _33639_, _03520_);
  or _83690_ (_33641_, _33640_, _33638_);
  and _83691_ (_33643_, _12456_, _05244_);
  or _83692_ (_33644_, _33539_, _03521_);
  or _83693_ (_33645_, _33644_, _33643_);
  and _83694_ (_33646_, _33645_, _42963_);
  and _83695_ (_33647_, _33646_, _33641_);
  nor _83696_ (_33648_, \oc8051_golden_model_1.P1 [2], rst);
  nor _83697_ (_33649_, _33648_, _00000_);
  or _83698_ (_43374_, _33649_, _33647_);
  and _83699_ (_33650_, _11197_, \oc8051_golden_model_1.P1 [3]);
  and _83700_ (_33651_, _12604_, _05244_);
  or _83701_ (_33653_, _33651_, _33650_);
  and _83702_ (_33654_, _33653_, _03769_);
  nor _83703_ (_33655_, _11197_, _04843_);
  or _83704_ (_33656_, _33655_, _33650_);
  or _83705_ (_33657_, _33656_, _06039_);
  nor _83706_ (_33658_, _12486_, _11197_);
  or _83707_ (_33659_, _33658_, _33650_);
  or _83708_ (_33660_, _33659_, _04444_);
  and _83709_ (_33661_, _05244_, \oc8051_golden_model_1.ACC [3]);
  or _83710_ (_33662_, _33661_, _33650_);
  and _83711_ (_33664_, _33662_, _04426_);
  and _83712_ (_33665_, _04427_, \oc8051_golden_model_1.P1 [3]);
  or _83713_ (_33666_, _33665_, _03570_);
  or _83714_ (_33667_, _33666_, _33664_);
  and _83715_ (_33668_, _33667_, _03517_);
  and _83716_ (_33669_, _33668_, _33660_);
  and _83717_ (_33670_, _11205_, \oc8051_golden_model_1.P1 [3]);
  and _83718_ (_33671_, _12490_, _05811_);
  or _83719_ (_33672_, _33671_, _33670_);
  and _83720_ (_33673_, _33672_, _03516_);
  or _83721_ (_33675_, _33673_, _03568_);
  or _83722_ (_33676_, _33675_, _33669_);
  or _83723_ (_33677_, _33656_, _03983_);
  and _83724_ (_33678_, _33677_, _33676_);
  or _83725_ (_33679_, _33678_, _03575_);
  or _83726_ (_33680_, _33662_, _03583_);
  and _83727_ (_33681_, _33680_, _03513_);
  and _83728_ (_33682_, _33681_, _33679_);
  and _83729_ (_33683_, _12500_, _05811_);
  or _83730_ (_33684_, _33683_, _33670_);
  and _83731_ (_33686_, _33684_, _03512_);
  or _83732_ (_33687_, _33686_, _03505_);
  or _83733_ (_33688_, _33687_, _33682_);
  or _83734_ (_33689_, _33670_, _12507_);
  and _83735_ (_33690_, _33689_, _33672_);
  or _83736_ (_33691_, _33690_, _03506_);
  and _83737_ (_33692_, _33691_, _03500_);
  and _83738_ (_33693_, _33692_, _33688_);
  and _83739_ (_33694_, _31314_, _05811_);
  or _83740_ (_33695_, _33694_, _33670_);
  and _83741_ (_33697_, _33695_, _03499_);
  or _83742_ (_33698_, _33697_, _07314_);
  or _83743_ (_33699_, _33698_, _33693_);
  and _83744_ (_33700_, _33699_, _33657_);
  or _83745_ (_33701_, _33700_, _03479_);
  and _83746_ (_33702_, _06717_, _05244_);
  or _83747_ (_33703_, _33650_, _06044_);
  or _83748_ (_33704_, _33703_, _33702_);
  and _83749_ (_33705_, _33704_, _03474_);
  and _83750_ (_33706_, _33705_, _33701_);
  and _83751_ (_33708_, _31341_, _05244_);
  or _83752_ (_33709_, _33708_, _33650_);
  and _83753_ (_33710_, _33709_, _03221_);
  or _83754_ (_33711_, _33710_, _03437_);
  or _83755_ (_33712_, _33711_, _33706_);
  and _83756_ (_33713_, _05244_, _06217_);
  or _83757_ (_33714_, _33713_, _33650_);
  or _83758_ (_33715_, _33714_, _03438_);
  and _83759_ (_33716_, _33715_, _33712_);
  or _83760_ (_33717_, _33716_, _03636_);
  and _83761_ (_33718_, _12598_, _05244_);
  or _83762_ (_33719_, _33718_, _33650_);
  or _83763_ (_33720_, _33719_, _04499_);
  and _83764_ (_33721_, _33720_, _04501_);
  and _83765_ (_33722_, _33721_, _33717_);
  or _83766_ (_33723_, _33722_, _33654_);
  and _83767_ (_33724_, _33723_, _05769_);
  or _83768_ (_33725_, _33650_, _05521_);
  and _83769_ (_33726_, _33725_, _03754_);
  and _83770_ (_33727_, _33726_, _33714_);
  or _83771_ (_33729_, _33727_, _33724_);
  and _83772_ (_33730_, _33729_, _03753_);
  and _83773_ (_33731_, _33662_, _03752_);
  and _83774_ (_33732_, _33731_, _33725_);
  or _83775_ (_33733_, _33732_, _03758_);
  or _83776_ (_33734_, _33733_, _33730_);
  nor _83777_ (_33735_, _12597_, _11197_);
  or _83778_ (_33736_, _33650_, _03759_);
  or _83779_ (_33737_, _33736_, _33735_);
  and _83780_ (_33738_, _33737_, _04517_);
  and _83781_ (_33740_, _33738_, _33734_);
  nor _83782_ (_33741_, _12603_, _11197_);
  or _83783_ (_33742_, _33741_, _33650_);
  and _83784_ (_33743_, _33742_, _03760_);
  or _83785_ (_33744_, _33743_, _03790_);
  or _83786_ (_33745_, _33744_, _33740_);
  or _83787_ (_33746_, _33659_, _04192_);
  and _83788_ (_33747_, _33746_, _03152_);
  and _83789_ (_33748_, _33747_, _33745_);
  and _83790_ (_33749_, _33684_, _03151_);
  or _83791_ (_33751_, _33749_, _03520_);
  or _83792_ (_33752_, _33751_, _33748_);
  and _83793_ (_33753_, _12658_, _05244_);
  or _83794_ (_33754_, _33650_, _03521_);
  or _83795_ (_33755_, _33754_, _33753_);
  and _83796_ (_33756_, _33755_, _42963_);
  and _83797_ (_33757_, _33756_, _33752_);
  nor _83798_ (_33758_, \oc8051_golden_model_1.P1 [3], rst);
  nor _83799_ (_33759_, _33758_, _00000_);
  or _83800_ (_43375_, _33759_, _33757_);
  and _83801_ (_33761_, _11197_, \oc8051_golden_model_1.P1 [4]);
  and _83802_ (_33762_, _12844_, _05244_);
  or _83803_ (_33763_, _33762_, _33761_);
  and _83804_ (_33764_, _33763_, _03769_);
  nor _83805_ (_33765_, _05712_, _11197_);
  or _83806_ (_33766_, _33765_, _33761_);
  or _83807_ (_33767_, _33766_, _06039_);
  nor _83808_ (_33768_, _12733_, _11197_);
  or _83809_ (_33769_, _33768_, _33761_);
  or _83810_ (_33770_, _33769_, _04444_);
  and _83811_ (_33772_, _05244_, \oc8051_golden_model_1.ACC [4]);
  or _83812_ (_33773_, _33772_, _33761_);
  and _83813_ (_33774_, _33773_, _04426_);
  and _83814_ (_33775_, _04427_, \oc8051_golden_model_1.P1 [4]);
  or _83815_ (_33776_, _33775_, _03570_);
  or _83816_ (_33777_, _33776_, _33774_);
  and _83817_ (_33778_, _33777_, _03517_);
  and _83818_ (_33779_, _33778_, _33770_);
  and _83819_ (_33780_, _11205_, \oc8051_golden_model_1.P1 [4]);
  and _83820_ (_33781_, _12737_, _05811_);
  or _83821_ (_33783_, _33781_, _33780_);
  and _83822_ (_33784_, _33783_, _03516_);
  or _83823_ (_33785_, _33784_, _03568_);
  or _83824_ (_33786_, _33785_, _33779_);
  or _83825_ (_33787_, _33766_, _03983_);
  and _83826_ (_33788_, _33787_, _33786_);
  or _83827_ (_33789_, _33788_, _03575_);
  or _83828_ (_33790_, _33773_, _03583_);
  and _83829_ (_33791_, _33790_, _03513_);
  and _83830_ (_33792_, _33791_, _33789_);
  and _83831_ (_33794_, _12718_, _05811_);
  or _83832_ (_33795_, _33794_, _33780_);
  and _83833_ (_33796_, _33795_, _03512_);
  or _83834_ (_33797_, _33796_, _03505_);
  or _83835_ (_33798_, _33797_, _33792_);
  or _83836_ (_33799_, _33780_, _12752_);
  and _83837_ (_33800_, _33799_, _33783_);
  or _83838_ (_33801_, _33800_, _03506_);
  and _83839_ (_33802_, _33801_, _03500_);
  and _83840_ (_33803_, _33802_, _33798_);
  and _83841_ (_33805_, _31439_, _05811_);
  or _83842_ (_33806_, _33805_, _33780_);
  and _83843_ (_33807_, _33806_, _03499_);
  or _83844_ (_33808_, _33807_, _07314_);
  or _83845_ (_33809_, _33808_, _33803_);
  and _83846_ (_33810_, _33809_, _33767_);
  or _83847_ (_33811_, _33810_, _03479_);
  and _83848_ (_33812_, _06722_, _05244_);
  or _83849_ (_33813_, _33761_, _06044_);
  or _83850_ (_33814_, _33813_, _33812_);
  and _83851_ (_33816_, _33814_, _03474_);
  and _83852_ (_33817_, _33816_, _33811_);
  and _83853_ (_33818_, _31468_, _05244_);
  or _83854_ (_33819_, _33818_, _33761_);
  and _83855_ (_33820_, _33819_, _03221_);
  or _83856_ (_33821_, _33820_, _03437_);
  or _83857_ (_33822_, _33821_, _33817_);
  and _83858_ (_33823_, _06233_, _05244_);
  or _83859_ (_33824_, _33823_, _33761_);
  or _83860_ (_33825_, _33824_, _03438_);
  and _83861_ (_33827_, _33825_, _33822_);
  or _83862_ (_33828_, _33827_, _03636_);
  and _83863_ (_33829_, _12711_, _05244_);
  or _83864_ (_33830_, _33829_, _33761_);
  or _83865_ (_33831_, _33830_, _04499_);
  and _83866_ (_33832_, _33831_, _04501_);
  and _83867_ (_33833_, _33832_, _33828_);
  or _83868_ (_33834_, _33833_, _33764_);
  and _83869_ (_33835_, _33834_, _05769_);
  or _83870_ (_33836_, _33761_, _05761_);
  and _83871_ (_33838_, _33836_, _03754_);
  and _83872_ (_33839_, _33838_, _33824_);
  or _83873_ (_33840_, _33839_, _33835_);
  and _83874_ (_33841_, _33840_, _03753_);
  and _83875_ (_33842_, _33773_, _03752_);
  and _83876_ (_33843_, _33842_, _33836_);
  or _83877_ (_33844_, _33843_, _03758_);
  or _83878_ (_33845_, _33844_, _33841_);
  nor _83879_ (_33846_, _12710_, _11197_);
  or _83880_ (_33847_, _33761_, _03759_);
  or _83881_ (_33849_, _33847_, _33846_);
  and _83882_ (_33850_, _33849_, _04517_);
  and _83883_ (_33851_, _33850_, _33845_);
  nor _83884_ (_33852_, _12843_, _11197_);
  or _83885_ (_33853_, _33852_, _33761_);
  and _83886_ (_33854_, _33853_, _03760_);
  or _83887_ (_33855_, _33854_, _03790_);
  or _83888_ (_33856_, _33855_, _33851_);
  or _83889_ (_33857_, _33769_, _04192_);
  and _83890_ (_33858_, _33857_, _03152_);
  and _83891_ (_33860_, _33858_, _33856_);
  and _83892_ (_33861_, _33795_, _03151_);
  or _83893_ (_33862_, _33861_, _03520_);
  or _83894_ (_33863_, _33862_, _33860_);
  and _83895_ (_33864_, _12893_, _05244_);
  or _83896_ (_33865_, _33761_, _03521_);
  or _83897_ (_33866_, _33865_, _33864_);
  and _83898_ (_33867_, _33866_, _42963_);
  and _83899_ (_33868_, _33867_, _33863_);
  nor _83900_ (_33869_, \oc8051_golden_model_1.P1 [4], rst);
  nor _83901_ (_33871_, _33869_, _00000_);
  or _83902_ (_43376_, _33871_, _33868_);
  and _83903_ (_33872_, _11197_, \oc8051_golden_model_1.P1 [5]);
  and _83904_ (_33873_, _13042_, _05244_);
  or _83905_ (_33874_, _33873_, _33872_);
  and _83906_ (_33875_, _33874_, _03769_);
  nor _83907_ (_33876_, _05422_, _11197_);
  or _83908_ (_33877_, _33876_, _33872_);
  or _83909_ (_33878_, _33877_, _06039_);
  nor _83910_ (_33879_, _12930_, _11197_);
  or _83911_ (_33881_, _33879_, _33872_);
  or _83912_ (_33882_, _33881_, _04444_);
  and _83913_ (_33883_, _05244_, \oc8051_golden_model_1.ACC [5]);
  or _83914_ (_33884_, _33883_, _33872_);
  and _83915_ (_33885_, _33884_, _04426_);
  and _83916_ (_33886_, _04427_, \oc8051_golden_model_1.P1 [5]);
  or _83917_ (_33887_, _33886_, _03570_);
  or _83918_ (_33888_, _33887_, _33885_);
  and _83919_ (_33889_, _33888_, _03517_);
  and _83920_ (_33890_, _33889_, _33882_);
  and _83921_ (_33891_, _11205_, \oc8051_golden_model_1.P1 [5]);
  and _83922_ (_33892_, _12934_, _05811_);
  or _83923_ (_33893_, _33892_, _33891_);
  and _83924_ (_33894_, _33893_, _03516_);
  or _83925_ (_33895_, _33894_, _03568_);
  or _83926_ (_33896_, _33895_, _33890_);
  or _83927_ (_33897_, _33877_, _03983_);
  and _83928_ (_33898_, _33897_, _33896_);
  or _83929_ (_33899_, _33898_, _03575_);
  or _83930_ (_33900_, _33884_, _03583_);
  and _83931_ (_33903_, _33900_, _03513_);
  and _83932_ (_33904_, _33903_, _33899_);
  and _83933_ (_33905_, _12914_, _05811_);
  or _83934_ (_33906_, _33905_, _33891_);
  and _83935_ (_33907_, _33906_, _03512_);
  or _83936_ (_33908_, _33907_, _03505_);
  or _83937_ (_33909_, _33908_, _33904_);
  or _83938_ (_33910_, _33891_, _12949_);
  and _83939_ (_33911_, _33910_, _33893_);
  or _83940_ (_33912_, _33911_, _03506_);
  and _83941_ (_33914_, _33912_, _03500_);
  and _83942_ (_33915_, _33914_, _33909_);
  and _83943_ (_33916_, _31567_, _05811_);
  or _83944_ (_33917_, _33916_, _33891_);
  and _83945_ (_33918_, _33917_, _03499_);
  or _83946_ (_33919_, _33918_, _07314_);
  or _83947_ (_33920_, _33919_, _33915_);
  and _83948_ (_33921_, _33920_, _33878_);
  or _83949_ (_33922_, _33921_, _03479_);
  and _83950_ (_33923_, _06721_, _05244_);
  or _83951_ (_33925_, _33872_, _06044_);
  or _83952_ (_33926_, _33925_, _33923_);
  and _83953_ (_33927_, _33926_, _03474_);
  and _83954_ (_33928_, _33927_, _33922_);
  and _83955_ (_33929_, _31593_, _05244_);
  or _83956_ (_33930_, _33929_, _33872_);
  and _83957_ (_33931_, _33930_, _03221_);
  or _83958_ (_33932_, _33931_, _03437_);
  or _83959_ (_33933_, _33932_, _33928_);
  and _83960_ (_33934_, _06211_, _05244_);
  or _83961_ (_33936_, _33934_, _33872_);
  or _83962_ (_33937_, _33936_, _03438_);
  and _83963_ (_33938_, _33937_, _33933_);
  or _83964_ (_33939_, _33938_, _03636_);
  and _83965_ (_33940_, _13036_, _05244_);
  or _83966_ (_33941_, _33940_, _33872_);
  or _83967_ (_33942_, _33941_, _04499_);
  and _83968_ (_33943_, _33942_, _04501_);
  and _83969_ (_33944_, _33943_, _33939_);
  or _83970_ (_33945_, _33944_, _33875_);
  and _83971_ (_33947_, _33945_, _05769_);
  or _83972_ (_33948_, _33872_, _05472_);
  and _83973_ (_33949_, _33948_, _03754_);
  and _83974_ (_33950_, _33949_, _33936_);
  or _83975_ (_33951_, _33950_, _33947_);
  and _83976_ (_33952_, _33951_, _03753_);
  and _83977_ (_33953_, _33884_, _03752_);
  and _83978_ (_33954_, _33953_, _33948_);
  or _83979_ (_33955_, _33954_, _03758_);
  or _83980_ (_33956_, _33955_, _33952_);
  nor _83981_ (_33958_, _13035_, _11197_);
  or _83982_ (_33959_, _33872_, _03759_);
  or _83983_ (_33960_, _33959_, _33958_);
  and _83984_ (_33961_, _33960_, _04517_);
  and _83985_ (_33962_, _33961_, _33956_);
  nor _83986_ (_33963_, _13041_, _11197_);
  or _83987_ (_33964_, _33963_, _33872_);
  and _83988_ (_33965_, _33964_, _03760_);
  or _83989_ (_33966_, _33965_, _03790_);
  or _83990_ (_33967_, _33966_, _33962_);
  or _83991_ (_33969_, _33881_, _04192_);
  and _83992_ (_33970_, _33969_, _03152_);
  and _83993_ (_33971_, _33970_, _33967_);
  and _83994_ (_33972_, _33906_, _03151_);
  or _83995_ (_33973_, _33972_, _03520_);
  or _83996_ (_33974_, _33973_, _33971_);
  and _83997_ (_33975_, _13097_, _05244_);
  or _83998_ (_33976_, _33872_, _03521_);
  or _83999_ (_33977_, _33976_, _33975_);
  and _84000_ (_33978_, _33977_, _42963_);
  and _84001_ (_33980_, _33978_, _33974_);
  nor _84002_ (_33981_, \oc8051_golden_model_1.P1 [5], rst);
  nor _84003_ (_33982_, _33981_, _00000_);
  or _84004_ (_43377_, _33982_, _33980_);
  and _84005_ (_33983_, _11197_, \oc8051_golden_model_1.P1 [6]);
  and _84006_ (_33984_, _13259_, _05244_);
  or _84007_ (_33985_, _33984_, _33983_);
  and _84008_ (_33986_, _33985_, _03769_);
  nor _84009_ (_33987_, _05327_, _11197_);
  or _84010_ (_33988_, _33987_, _33983_);
  or _84011_ (_33990_, _33988_, _06039_);
  nor _84012_ (_33991_, _13122_, _11197_);
  or _84013_ (_33992_, _33991_, _33983_);
  or _84014_ (_33993_, _33992_, _04444_);
  and _84015_ (_33994_, _05244_, \oc8051_golden_model_1.ACC [6]);
  or _84016_ (_33995_, _33994_, _33983_);
  and _84017_ (_33996_, _33995_, _04426_);
  and _84018_ (_33997_, _04427_, \oc8051_golden_model_1.P1 [6]);
  or _84019_ (_33998_, _33997_, _03570_);
  or _84020_ (_33999_, _33998_, _33996_);
  and _84021_ (_34001_, _33999_, _03517_);
  and _84022_ (_34002_, _34001_, _33993_);
  and _84023_ (_34003_, _11205_, \oc8051_golden_model_1.P1 [6]);
  and _84024_ (_34004_, _13145_, _05811_);
  or _84025_ (_34005_, _34004_, _34003_);
  and _84026_ (_34006_, _34005_, _03516_);
  or _84027_ (_34007_, _34006_, _03568_);
  or _84028_ (_34008_, _34007_, _34002_);
  or _84029_ (_34009_, _33988_, _03983_);
  and _84030_ (_34010_, _34009_, _34008_);
  or _84031_ (_34012_, _34010_, _03575_);
  or _84032_ (_34013_, _33995_, _03583_);
  and _84033_ (_34014_, _34013_, _03513_);
  and _84034_ (_34015_, _34014_, _34012_);
  and _84035_ (_34016_, _13130_, _05811_);
  or _84036_ (_34017_, _34016_, _34003_);
  and _84037_ (_34018_, _34017_, _03512_);
  or _84038_ (_34019_, _34018_, _03505_);
  or _84039_ (_34020_, _34019_, _34015_);
  or _84040_ (_34021_, _34003_, _13160_);
  and _84041_ (_34023_, _34021_, _34005_);
  or _84042_ (_34024_, _34023_, _03506_);
  and _84043_ (_34025_, _34024_, _03500_);
  and _84044_ (_34026_, _34025_, _34020_);
  and _84045_ (_34027_, _31693_, _05811_);
  or _84046_ (_34028_, _34027_, _34003_);
  and _84047_ (_34029_, _34028_, _03499_);
  or _84048_ (_34030_, _34029_, _07314_);
  or _84049_ (_34031_, _34030_, _34026_);
  and _84050_ (_34032_, _34031_, _33990_);
  or _84051_ (_34034_, _34032_, _03479_);
  and _84052_ (_34035_, _06713_, _05244_);
  or _84053_ (_34036_, _33983_, _06044_);
  or _84054_ (_34037_, _34036_, _34035_);
  and _84055_ (_34038_, _34037_, _03474_);
  and _84056_ (_34039_, _34038_, _34034_);
  and _84057_ (_34040_, _31718_, _05244_);
  or _84058_ (_34041_, _34040_, _33983_);
  and _84059_ (_34042_, _34041_, _03221_);
  or _84060_ (_34043_, _34042_, _03437_);
  or _84061_ (_34045_, _34043_, _34039_);
  and _84062_ (_34046_, _13244_, _05244_);
  or _84063_ (_34047_, _34046_, _33983_);
  or _84064_ (_34048_, _34047_, _03438_);
  and _84065_ (_34049_, _34048_, _34045_);
  or _84066_ (_34050_, _34049_, _03636_);
  and _84067_ (_34051_, _13253_, _05244_);
  or _84068_ (_34052_, _34051_, _33983_);
  or _84069_ (_34053_, _34052_, _04499_);
  and _84070_ (_34054_, _34053_, _04501_);
  and _84071_ (_34056_, _34054_, _34050_);
  or _84072_ (_34057_, _34056_, _33986_);
  and _84073_ (_34058_, _34057_, _05769_);
  or _84074_ (_34059_, _33983_, _05377_);
  and _84075_ (_34060_, _34059_, _03754_);
  and _84076_ (_34061_, _34060_, _34047_);
  or _84077_ (_34062_, _34061_, _34058_);
  and _84078_ (_34063_, _34062_, _03753_);
  and _84079_ (_34064_, _33995_, _03752_);
  and _84080_ (_34065_, _34064_, _34059_);
  or _84081_ (_34067_, _34065_, _03758_);
  or _84082_ (_34068_, _34067_, _34063_);
  nor _84083_ (_34069_, _13251_, _11197_);
  or _84084_ (_34070_, _33983_, _03759_);
  or _84085_ (_34071_, _34070_, _34069_);
  and _84086_ (_34072_, _34071_, _04517_);
  and _84087_ (_34073_, _34072_, _34068_);
  nor _84088_ (_34074_, _13258_, _11197_);
  or _84089_ (_34075_, _34074_, _33983_);
  and _84090_ (_34076_, _34075_, _03760_);
  or _84091_ (_34078_, _34076_, _03790_);
  or _84092_ (_34079_, _34078_, _34073_);
  or _84093_ (_34080_, _33992_, _04192_);
  and _84094_ (_34081_, _34080_, _03152_);
  and _84095_ (_34082_, _34081_, _34079_);
  and _84096_ (_34083_, _34017_, _03151_);
  or _84097_ (_34084_, _34083_, _03520_);
  or _84098_ (_34085_, _34084_, _34082_);
  and _84099_ (_34086_, _13312_, _05244_);
  or _84100_ (_34087_, _33983_, _03521_);
  or _84101_ (_34089_, _34087_, _34086_);
  and _84102_ (_34090_, _34089_, _42963_);
  and _84103_ (_34091_, _34090_, _34085_);
  nor _84104_ (_34092_, \oc8051_golden_model_1.P1 [6], rst);
  nor _84105_ (_34093_, _34092_, _00000_);
  or _84106_ (_43378_, _34093_, _34091_);
  nor _84107_ (_34094_, \oc8051_golden_model_1.SP [0], rst);
  nor _84108_ (_34095_, _34094_, _00000_);
  and _84109_ (_34096_, _05269_, _04419_);
  nor _84110_ (_34097_, _05269_, _03502_);
  or _84111_ (_34099_, _34097_, _06039_);
  or _84112_ (_34100_, _34099_, _34096_);
  and _84113_ (_34101_, _05941_, _05269_);
  or _84114_ (_34102_, _34101_, _34097_);
  or _84115_ (_34103_, _34102_, _04444_);
  and _84116_ (_34104_, _05269_, \oc8051_golden_model_1.ACC [0]);
  or _84117_ (_34105_, _34104_, _34097_);
  and _84118_ (_34106_, _34105_, _04426_);
  nor _84119_ (_34107_, _04426_, _03502_);
  or _84120_ (_34108_, _34107_, _03570_);
  or _84121_ (_34110_, _34108_, _34106_);
  and _84122_ (_34111_, _34110_, _03983_);
  and _84123_ (_34112_, _34111_, _34103_);
  or _84124_ (_34113_, _04031_, _03575_);
  or _84125_ (_34114_, _34113_, _34112_);
  or _84126_ (_34115_, _34105_, _03583_);
  and _84127_ (_34116_, _34115_, _04887_);
  and _84128_ (_34117_, _34116_, _34114_);
  nand _84129_ (_34118_, _06039_, _04469_);
  or _84130_ (_34119_, _34118_, _34117_);
  and _84131_ (_34121_, _34119_, _34100_);
  or _84132_ (_34122_, _34121_, _03479_);
  and _84133_ (_34123_, _06715_, _05269_);
  or _84134_ (_34124_, _34097_, _06044_);
  or _84135_ (_34125_, _34124_, _34123_);
  and _84136_ (_34126_, _34125_, _34122_);
  or _84137_ (_34127_, _34126_, _03221_);
  nor _84138_ (_34128_, _11975_, _11355_);
  or _84139_ (_34129_, _34128_, _34097_);
  or _84140_ (_34130_, _34129_, _03474_);
  and _84141_ (_34132_, _34130_, _03438_);
  and _84142_ (_34133_, _34132_, _34127_);
  and _84143_ (_34134_, _05269_, _06202_);
  or _84144_ (_34135_, _34134_, _34097_);
  and _84145_ (_34136_, _34135_, _03437_);
  or _84146_ (_34137_, _34136_, _03636_);
  or _84147_ (_34138_, _34137_, _34133_);
  and _84148_ (_34139_, _11990_, _05269_);
  or _84149_ (_34140_, _34139_, _34097_);
  or _84150_ (_34141_, _34140_, _04499_);
  and _84151_ (_34143_, _34141_, _34138_);
  or _84152_ (_34144_, _34143_, _03769_);
  and _84153_ (_34145_, _11995_, _05269_);
  or _84154_ (_34146_, _34145_, _34097_);
  or _84155_ (_34147_, _34146_, _04501_);
  and _84156_ (_34148_, _34147_, _05769_);
  and _84157_ (_34149_, _34148_, _34144_);
  nand _84158_ (_34150_, _34135_, _04504_);
  nor _84159_ (_34151_, _34150_, _34101_);
  or _84160_ (_34152_, _34151_, _34149_);
  and _84161_ (_34154_, _34152_, _03753_);
  or _84162_ (_34155_, _34097_, _05617_);
  and _84163_ (_34156_, _34105_, _03752_);
  and _84164_ (_34157_, _34156_, _34155_);
  or _84165_ (_34158_, _34157_, _03758_);
  or _84166_ (_34159_, _34158_, _34154_);
  nor _84167_ (_34160_, _11988_, _11355_);
  or _84168_ (_34161_, _34097_, _03759_);
  or _84169_ (_34162_, _34161_, _34160_);
  and _84170_ (_34163_, _34162_, _04517_);
  and _84171_ (_34164_, _34163_, _34159_);
  nor _84172_ (_34165_, _11870_, _11355_);
  or _84173_ (_34166_, _34165_, _34097_);
  and _84174_ (_34167_, _34166_, _03760_);
  or _84175_ (_34168_, _34167_, _17076_);
  or _84176_ (_34169_, _34168_, _34164_);
  or _84177_ (_34170_, _34102_, _03882_);
  and _84178_ (_34171_, _34170_, _42963_);
  and _84179_ (_34172_, _34171_, _34169_);
  or _84180_ (_43379_, _34172_, _34095_);
  nor _84181_ (_34175_, _05269_, _04333_);
  and _84182_ (_34176_, _12252_, _05269_);
  or _84183_ (_34177_, _34176_, _34175_);
  and _84184_ (_34178_, _34177_, _03520_);
  nand _84185_ (_34179_, _03775_, \oc8051_golden_model_1.SP [1]);
  not _84186_ (_34180_, _34176_);
  or _84187_ (_34181_, _05269_, \oc8051_golden_model_1.SP [1]);
  and _84188_ (_34182_, _34181_, _34180_);
  or _84189_ (_34183_, _34182_, _04444_);
  nand _84190_ (_34184_, _03923_, \oc8051_golden_model_1.SP [1]);
  nand _84191_ (_34186_, _05269_, _03233_);
  and _84192_ (_34187_, _34186_, _34181_);
  and _84193_ (_34188_, _34187_, _04426_);
  nor _84194_ (_34189_, _04426_, _04333_);
  or _84195_ (_34190_, _34189_, _03923_);
  or _84196_ (_34191_, _34190_, _34188_);
  and _84197_ (_34192_, _34191_, _34184_);
  or _84198_ (_34193_, _34192_, _03570_);
  and _84199_ (_34194_, _34193_, _03203_);
  and _84200_ (_34195_, _34194_, _34183_);
  nor _84201_ (_34197_, _03203_, \oc8051_golden_model_1.SP [1]);
  or _84202_ (_34198_, _34197_, _03568_);
  or _84203_ (_34199_, _34198_, _34195_);
  nand _84204_ (_34200_, _04553_, _03568_);
  and _84205_ (_34201_, _34200_, _34199_);
  or _84206_ (_34202_, _34201_, _03575_);
  or _84207_ (_34203_, _34187_, _03583_);
  and _84208_ (_34204_, _34203_, _04887_);
  and _84209_ (_34205_, _34204_, _34202_);
  or _84210_ (_34206_, _04744_, _04640_);
  or _84211_ (_34208_, _34206_, _34205_);
  nand _84212_ (_34209_, _04744_, \oc8051_golden_model_1.SP [1]);
  and _84213_ (_34210_, _34209_, _06039_);
  and _84214_ (_34211_, _34210_, _34208_);
  nand _84215_ (_34212_, _05269_, _04603_);
  and _84216_ (_34213_, _34181_, _07314_);
  and _84217_ (_34214_, _34213_, _34212_);
  or _84218_ (_34215_, _34214_, _03479_);
  or _84219_ (_34216_, _34215_, _34211_);
  and _84220_ (_34217_, _06714_, _05269_);
  or _84221_ (_34219_, _34175_, _06044_);
  or _84222_ (_34220_, _34219_, _34217_);
  and _84223_ (_34221_, _34220_, _03474_);
  and _84224_ (_34222_, _34221_, _34216_);
  nand _84225_ (_34223_, _12176_, _05269_);
  and _84226_ (_34224_, _34181_, _03221_);
  and _84227_ (_34225_, _34224_, _34223_);
  or _84228_ (_34226_, _34225_, _34222_);
  and _84229_ (_34227_, _34226_, _03438_);
  nand _84230_ (_34228_, _05269_, _04317_);
  and _84231_ (_34230_, _34181_, _03437_);
  and _84232_ (_34231_, _34230_, _34228_);
  or _84233_ (_34232_, _34231_, _03189_);
  or _84234_ (_34233_, _34232_, _34227_);
  and _84235_ (_34234_, _03189_, \oc8051_golden_model_1.SP [1]);
  nor _84236_ (_34235_, _34234_, _03636_);
  and _84237_ (_34236_, _34235_, _34233_);
  or _84238_ (_34237_, _12191_, _11355_);
  and _84239_ (_34238_, _34181_, _03636_);
  and _84240_ (_34239_, _34238_, _34237_);
  or _84241_ (_34241_, _34239_, _34236_);
  and _84242_ (_34242_, _34241_, _04501_);
  or _84243_ (_34243_, _12197_, _11355_);
  and _84244_ (_34244_, _34181_, _03769_);
  and _84245_ (_34245_, _34244_, _34243_);
  or _84246_ (_34246_, _34245_, _34242_);
  and _84247_ (_34247_, _34246_, _05769_);
  or _84248_ (_34248_, _12190_, _11355_);
  and _84249_ (_34249_, _34248_, _03754_);
  and _84250_ (_34250_, _34249_, _34181_);
  or _84251_ (_34252_, _34250_, _34247_);
  and _84252_ (_34253_, _34252_, _09960_);
  and _84253_ (_34254_, _03192_, _04333_);
  or _84254_ (_34255_, _34175_, _05569_);
  and _84255_ (_34256_, _34187_, _03752_);
  and _84256_ (_34257_, _34256_, _34255_);
  or _84257_ (_34258_, _34257_, _34254_);
  or _84258_ (_34259_, _34258_, _34253_);
  and _84259_ (_34260_, _34259_, _03759_);
  or _84260_ (_34261_, _34228_, _05569_);
  and _84261_ (_34263_, _34181_, _03758_);
  and _84262_ (_34264_, _34263_, _34261_);
  or _84263_ (_34265_, _34264_, _34260_);
  and _84264_ (_34266_, _34265_, _04517_);
  or _84265_ (_34267_, _34186_, _05569_);
  and _84266_ (_34268_, _34181_, _03760_);
  and _84267_ (_34269_, _34268_, _34267_);
  or _84268_ (_34270_, _34269_, _03775_);
  or _84269_ (_34271_, _34270_, _34266_);
  nand _84270_ (_34272_, _34271_, _34179_);
  nor _84271_ (_34274_, _03522_, _03179_);
  nand _84272_ (_34275_, _34274_, _34272_);
  or _84273_ (_34276_, _34274_, _04333_);
  and _84274_ (_34277_, _34276_, _04192_);
  and _84275_ (_34278_, _34277_, _34275_);
  and _84276_ (_34279_, _34182_, _03790_);
  or _84277_ (_34280_, _34279_, _04947_);
  or _84278_ (_34281_, _34280_, _34278_);
  or _84279_ (_34282_, _04533_, _04333_);
  and _84280_ (_34283_, _34282_, _03521_);
  and _84281_ (_34285_, _34283_, _34281_);
  or _84282_ (_34286_, _34285_, _34178_);
  and _84283_ (_34287_, _34286_, _42963_);
  nor _84284_ (_34288_, \oc8051_golden_model_1.SP [1], rst);
  nor _84285_ (_34289_, _34288_, _00000_);
  or _84286_ (_43380_, _34289_, _34287_);
  nor _84287_ (_34290_, _42963_, _03982_);
  or _84288_ (_34291_, _34290_, rst);
  nor _84289_ (_34292_, _05269_, _03982_);
  and _84290_ (_34293_, _12401_, _05269_);
  or _84291_ (_34295_, _34293_, _34292_);
  and _84292_ (_34296_, _34295_, _03769_);
  nor _84293_ (_34297_, _11355_, _05026_);
  or _84294_ (_34298_, _34292_, _06039_);
  or _84295_ (_34299_, _34298_, _34297_);
  or _84296_ (_34300_, _05053_, _04743_);
  nor _84297_ (_34301_, _12282_, _11355_);
  or _84298_ (_34302_, _34301_, _34292_);
  or _84299_ (_34303_, _34302_, _04444_);
  and _84300_ (_34304_, _05269_, \oc8051_golden_model_1.ACC [2]);
  or _84301_ (_34306_, _34304_, _34292_);
  or _84302_ (_34307_, _34306_, _04427_);
  or _84303_ (_34308_, _04426_, \oc8051_golden_model_1.SP [2]);
  and _84304_ (_34309_, _34308_, _04762_);
  and _84305_ (_34310_, _34309_, _34307_);
  and _84306_ (_34311_, _05110_, _03923_);
  or _84307_ (_34312_, _34311_, _03570_);
  or _84308_ (_34313_, _34312_, _34310_);
  and _84309_ (_34314_, _34313_, _03203_);
  and _84310_ (_34315_, _34314_, _34303_);
  nor _84311_ (_34317_, _12674_, _03203_);
  or _84312_ (_34318_, _34317_, _03568_);
  or _84313_ (_34319_, _34318_, _34315_);
  nand _84314_ (_34320_, _05866_, _03568_);
  and _84315_ (_34321_, _34320_, _34319_);
  or _84316_ (_34322_, _34321_, _03575_);
  or _84317_ (_34323_, _34306_, _03583_);
  and _84318_ (_34324_, _34323_, _04887_);
  and _84319_ (_34325_, _34324_, _34322_);
  or _84320_ (_34326_, _34325_, _34300_);
  nor _84321_ (_34328_, _05110_, _03200_);
  nor _84322_ (_34329_, _34328_, _03223_);
  and _84323_ (_34330_, _34329_, _34326_);
  nand _84324_ (_34331_, _05110_, _03223_);
  nand _84325_ (_34332_, _34331_, _06039_);
  or _84326_ (_34333_, _34332_, _34330_);
  and _84327_ (_34334_, _34333_, _34299_);
  or _84328_ (_34335_, _34334_, _03479_);
  and _84329_ (_34336_, _06718_, _05269_);
  or _84330_ (_34337_, _34292_, _06044_);
  or _84331_ (_34339_, _34337_, _34336_);
  and _84332_ (_34340_, _34339_, _34335_);
  or _84333_ (_34341_, _34340_, _03221_);
  nor _84334_ (_34342_, _12384_, _11355_);
  or _84335_ (_34343_, _34342_, _34292_);
  or _84336_ (_34344_, _34343_, _03474_);
  and _84337_ (_34345_, _34344_, _03438_);
  and _84338_ (_34346_, _34345_, _34341_);
  and _84339_ (_34347_, _05269_, _06261_);
  or _84340_ (_34348_, _34347_, _34292_);
  and _84341_ (_34350_, _34348_, _03437_);
  or _84342_ (_34351_, _34350_, _03189_);
  or _84343_ (_34352_, _34351_, _34346_);
  nand _84344_ (_34353_, _12674_, _03189_);
  and _84345_ (_34354_, _34353_, _34352_);
  or _84346_ (_34355_, _34354_, _03636_);
  and _84347_ (_34356_, _12273_, _05269_);
  or _84348_ (_34357_, _34356_, _34292_);
  or _84349_ (_34358_, _34357_, _04499_);
  and _84350_ (_34359_, _34358_, _04501_);
  and _84351_ (_34361_, _34359_, _34355_);
  or _84352_ (_34362_, _34361_, _34296_);
  and _84353_ (_34363_, _34362_, _05769_);
  or _84354_ (_34364_, _34292_, _05665_);
  and _84355_ (_34365_, _34348_, _04504_);
  and _84356_ (_34366_, _34365_, _34364_);
  or _84357_ (_34367_, _34366_, _34363_);
  and _84358_ (_34368_, _34367_, _09960_);
  and _84359_ (_34369_, _34306_, _03752_);
  and _84360_ (_34370_, _34369_, _34364_);
  and _84361_ (_34372_, _05110_, _03192_);
  or _84362_ (_34373_, _34372_, _03758_);
  or _84363_ (_34374_, _34373_, _34370_);
  or _84364_ (_34375_, _34374_, _34368_);
  nor _84365_ (_34376_, _12272_, _11355_);
  or _84366_ (_34377_, _34376_, _34292_);
  or _84367_ (_34378_, _34377_, _03759_);
  and _84368_ (_34379_, _34378_, _34375_);
  or _84369_ (_34380_, _34379_, _03760_);
  nor _84370_ (_34381_, _12400_, _11355_);
  or _84371_ (_34383_, _34381_, _34292_);
  or _84372_ (_34384_, _34383_, _04517_);
  and _84373_ (_34385_, _34384_, _11403_);
  and _84374_ (_34386_, _34385_, _34380_);
  and _84375_ (_34387_, _12674_, _03775_);
  or _84376_ (_34388_, _34387_, _03179_);
  or _84377_ (_34389_, _34388_, _34386_);
  nand _84378_ (_34390_, _12674_, _03179_);
  and _84379_ (_34391_, _34390_, _03523_);
  and _84380_ (_34392_, _34391_, _34389_);
  and _84381_ (_34394_, _12674_, _03522_);
  or _84382_ (_34395_, _34394_, _03790_);
  or _84383_ (_34396_, _34395_, _34392_);
  or _84384_ (_34397_, _34302_, _04192_);
  and _84385_ (_34398_, _34397_, _04533_);
  and _84386_ (_34399_, _34398_, _34396_);
  nor _84387_ (_34400_, _12674_, _04533_);
  or _84388_ (_34401_, _34400_, _03520_);
  or _84389_ (_34402_, _34401_, _34399_);
  and _84390_ (_34403_, _12456_, _05269_);
  or _84391_ (_34405_, _34292_, _03521_);
  or _84392_ (_34406_, _34405_, _34403_);
  and _84393_ (_34407_, _34406_, _42963_);
  and _84394_ (_34408_, _34407_, _34402_);
  or _84395_ (_43381_, _34408_, _34291_);
  nor _84396_ (_34409_, _42963_, _03567_);
  or _84397_ (_34410_, _05113_, _04533_);
  nor _84398_ (_34411_, _05269_, _03567_);
  nor _84399_ (_34412_, _12486_, _11355_);
  or _84400_ (_34413_, _34412_, _34411_);
  or _84401_ (_34415_, _34413_, _04444_);
  and _84402_ (_34416_, _05269_, \oc8051_golden_model_1.ACC [3]);
  or _84403_ (_34417_, _34416_, _34411_);
  or _84404_ (_34418_, _34417_, _04427_);
  or _84405_ (_34419_, _04426_, \oc8051_golden_model_1.SP [3]);
  and _84406_ (_34420_, _34419_, _04762_);
  and _84407_ (_34421_, _34420_, _34418_);
  and _84408_ (_34422_, _05113_, _03923_);
  or _84409_ (_34423_, _34422_, _03570_);
  or _84410_ (_34424_, _34423_, _34421_);
  and _84411_ (_34426_, _34424_, _03203_);
  and _84412_ (_34427_, _34426_, _34415_);
  nor _84413_ (_34428_, _12678_, _03203_);
  or _84414_ (_34429_, _34428_, _03568_);
  or _84415_ (_34430_, _34429_, _34427_);
  nand _84416_ (_34431_, _05854_, _03568_);
  and _84417_ (_34432_, _34431_, _34430_);
  or _84418_ (_34433_, _34432_, _03575_);
  or _84419_ (_34434_, _34417_, _03583_);
  and _84420_ (_34435_, _34434_, _04887_);
  and _84421_ (_34437_, _34435_, _34433_);
  or _84422_ (_34438_, _34437_, _04891_);
  and _84423_ (_34439_, _34438_, _04745_);
  nand _84424_ (_34440_, _05113_, _04744_);
  nand _84425_ (_34441_, _34440_, _06039_);
  or _84426_ (_34442_, _34441_, _34439_);
  nor _84427_ (_34443_, _11355_, _04843_);
  or _84428_ (_34444_, _34411_, _06039_);
  or _84429_ (_34445_, _34444_, _34443_);
  and _84430_ (_34446_, _34445_, _34442_);
  or _84431_ (_34448_, _34446_, _03479_);
  and _84432_ (_34449_, _06717_, _05269_);
  or _84433_ (_34450_, _34411_, _06044_);
  or _84434_ (_34451_, _34450_, _34449_);
  and _84435_ (_34452_, _34451_, _34448_);
  or _84436_ (_34453_, _34452_, _03221_);
  nor _84437_ (_34454_, _12583_, _11355_);
  or _84438_ (_34455_, _34454_, _34411_);
  or _84439_ (_34456_, _34455_, _03474_);
  and _84440_ (_34457_, _34456_, _34453_);
  or _84441_ (_34459_, _34457_, _03437_);
  and _84442_ (_34460_, _05269_, _06217_);
  or _84443_ (_34461_, _34460_, _34411_);
  or _84444_ (_34462_, _34461_, _03438_);
  and _84445_ (_34463_, _34462_, _11376_);
  and _84446_ (_34464_, _34463_, _34459_);
  and _84447_ (_34465_, _05113_, _03189_);
  or _84448_ (_34466_, _34465_, _03636_);
  or _84449_ (_34467_, _34466_, _34464_);
  and _84450_ (_34468_, _12598_, _05269_);
  or _84451_ (_34470_, _34468_, _34411_);
  or _84452_ (_34471_, _34470_, _04499_);
  and _84453_ (_34472_, _34471_, _34467_);
  or _84454_ (_34473_, _34472_, _03769_);
  and _84455_ (_34474_, _12604_, _05269_);
  or _84456_ (_34475_, _34474_, _34411_);
  or _84457_ (_34476_, _34475_, _04501_);
  and _84458_ (_34477_, _34476_, _05769_);
  and _84459_ (_34478_, _34477_, _34473_);
  or _84460_ (_34479_, _34411_, _05521_);
  and _84461_ (_34481_, _34479_, _03754_);
  and _84462_ (_34482_, _34481_, _34461_);
  or _84463_ (_34483_, _34482_, _34478_);
  and _84464_ (_34484_, _34483_, _09960_);
  and _84465_ (_34485_, _34417_, _03752_);
  and _84466_ (_34486_, _34485_, _34479_);
  and _84467_ (_34487_, _05113_, _03192_);
  or _84468_ (_34488_, _34487_, _03758_);
  or _84469_ (_34489_, _34488_, _34486_);
  or _84470_ (_34490_, _34489_, _34484_);
  nor _84471_ (_34492_, _12597_, _11355_);
  or _84472_ (_34493_, _34492_, _34411_);
  or _84473_ (_34494_, _34493_, _03759_);
  and _84474_ (_34495_, _34494_, _34490_);
  or _84475_ (_34496_, _34495_, _03760_);
  nor _84476_ (_34497_, _12603_, _11355_);
  or _84477_ (_34498_, _34497_, _34411_);
  or _84478_ (_34499_, _34498_, _04517_);
  and _84479_ (_34500_, _34499_, _11403_);
  and _84480_ (_34501_, _34500_, _34496_);
  nor _84481_ (_34503_, _05851_, _03567_);
  or _84482_ (_34504_, _34503_, _05852_);
  and _84483_ (_34505_, _34504_, _03775_);
  or _84484_ (_34506_, _34505_, _03179_);
  or _84485_ (_34507_, _34506_, _34501_);
  nand _84486_ (_34508_, _12678_, _03179_);
  and _84487_ (_34509_, _34508_, _34507_);
  or _84488_ (_34510_, _34509_, _03522_);
  or _84489_ (_34511_, _34504_, _03523_);
  and _84490_ (_34512_, _34511_, _04192_);
  and _84491_ (_34514_, _34512_, _34510_);
  and _84492_ (_34515_, _34413_, _03790_);
  or _84493_ (_34516_, _34515_, _04947_);
  or _84494_ (_34517_, _34516_, _34514_);
  and _84495_ (_34518_, _34517_, _34410_);
  or _84496_ (_34519_, _34518_, _03520_);
  and _84497_ (_34520_, _12658_, _05269_);
  or _84498_ (_34521_, _34411_, _03521_);
  or _84499_ (_34522_, _34521_, _34520_);
  and _84500_ (_34523_, _34522_, _42963_);
  and _84501_ (_34525_, _34523_, _34519_);
  or _84502_ (_34526_, _34525_, _34409_);
  and _84503_ (_43382_, _34526_, _41755_);
  nor _84504_ (_34527_, _05269_, _11330_);
  and _84505_ (_34528_, _12844_, _05269_);
  or _84506_ (_34529_, _34528_, _34527_);
  and _84507_ (_34530_, _34529_, _03769_);
  nor _84508_ (_34531_, _12733_, _11355_);
  or _84509_ (_34532_, _34531_, _34527_);
  or _84510_ (_34533_, _34532_, _04444_);
  and _84511_ (_34535_, _05269_, \oc8051_golden_model_1.ACC [4]);
  or _84512_ (_34536_, _34535_, _34527_);
  or _84513_ (_34537_, _34536_, _04427_);
  or _84514_ (_34538_, _04426_, \oc8051_golden_model_1.SP [4]);
  and _84515_ (_34539_, _34538_, _04762_);
  and _84516_ (_34540_, _34539_, _34537_);
  nor _84517_ (_34541_, _04849_, \oc8051_golden_model_1.SP [4]);
  nor _84518_ (_34542_, _34541_, _11300_);
  and _84519_ (_34543_, _34542_, _03923_);
  or _84520_ (_34544_, _34543_, _03570_);
  or _84521_ (_34546_, _34544_, _34540_);
  and _84522_ (_34547_, _34546_, _03203_);
  and _84523_ (_34548_, _34547_, _34533_);
  and _84524_ (_34549_, _34542_, _04746_);
  or _84525_ (_34550_, _34549_, _03568_);
  or _84526_ (_34551_, _34550_, _34548_);
  and _84527_ (_34552_, _11331_, _03502_);
  nor _84528_ (_34553_, _05853_, _11330_);
  nor _84529_ (_34554_, _34553_, _34552_);
  nand _84530_ (_34555_, _34554_, _03568_);
  and _84531_ (_34557_, _34555_, _34551_);
  or _84532_ (_34558_, _34557_, _03575_);
  or _84533_ (_34559_, _34536_, _03583_);
  and _84534_ (_34560_, _34559_, _04887_);
  and _84535_ (_34561_, _34560_, _34558_);
  and _84536_ (_34562_, _04850_, \oc8051_golden_model_1.SP [4]);
  nor _84537_ (_34563_, _04850_, \oc8051_golden_model_1.SP [4]);
  nor _84538_ (_34564_, _34563_, _34562_);
  and _84539_ (_34565_, _34564_, _03511_);
  or _84540_ (_34566_, _34565_, _04744_);
  or _84541_ (_34568_, _34566_, _34561_);
  or _84542_ (_34569_, _34542_, _04745_);
  and _84543_ (_34570_, _34569_, _06039_);
  and _84544_ (_34571_, _34570_, _34568_);
  nor _84545_ (_34572_, _05712_, _11355_);
  or _84546_ (_34573_, _34572_, _34527_);
  and _84547_ (_34574_, _34573_, _07314_);
  or _84548_ (_34575_, _34574_, _03479_);
  or _84549_ (_34576_, _34575_, _34571_);
  and _84550_ (_34577_, _06722_, _05269_);
  or _84551_ (_34579_, _34527_, _06044_);
  or _84552_ (_34580_, _34579_, _34577_);
  and _84553_ (_34581_, _34580_, _03474_);
  and _84554_ (_34582_, _34581_, _34576_);
  nor _84555_ (_34583_, _12827_, _11355_);
  or _84556_ (_34584_, _34583_, _34527_);
  and _84557_ (_34585_, _34584_, _03221_);
  or _84558_ (_34586_, _34585_, _03437_);
  or _84559_ (_34587_, _34586_, _34582_);
  and _84560_ (_34588_, _06233_, _05269_);
  or _84561_ (_34590_, _34588_, _34527_);
  or _84562_ (_34591_, _34590_, _03438_);
  and _84563_ (_34592_, _34591_, _34587_);
  or _84564_ (_34593_, _34592_, _03189_);
  or _84565_ (_34594_, _34542_, _11376_);
  and _84566_ (_34595_, _34594_, _34593_);
  or _84567_ (_34596_, _34595_, _03636_);
  and _84568_ (_34597_, _12711_, _05269_);
  or _84569_ (_34598_, _34597_, _34527_);
  or _84570_ (_34599_, _34598_, _04499_);
  and _84571_ (_34601_, _34599_, _04501_);
  and _84572_ (_34602_, _34601_, _34596_);
  or _84573_ (_34603_, _34602_, _34530_);
  and _84574_ (_34604_, _34603_, _05769_);
  or _84575_ (_34605_, _34527_, _05761_);
  and _84576_ (_34606_, _34605_, _03754_);
  and _84577_ (_34607_, _34606_, _34590_);
  or _84578_ (_34608_, _34607_, _34604_);
  and _84579_ (_34609_, _34608_, _09960_);
  and _84580_ (_34610_, _34536_, _03752_);
  and _84581_ (_34612_, _34610_, _34605_);
  and _84582_ (_34613_, _34542_, _03192_);
  or _84583_ (_34614_, _34613_, _03758_);
  or _84584_ (_34615_, _34614_, _34612_);
  or _84585_ (_34616_, _34615_, _34609_);
  nor _84586_ (_34617_, _12710_, _11355_);
  or _84587_ (_34618_, _34617_, _34527_);
  or _84588_ (_34619_, _34618_, _03759_);
  and _84589_ (_34620_, _34619_, _34616_);
  or _84590_ (_34621_, _34620_, _03760_);
  nor _84591_ (_34623_, _12843_, _11355_);
  or _84592_ (_34624_, _34623_, _34527_);
  or _84593_ (_34625_, _34624_, _04517_);
  and _84594_ (_34626_, _34625_, _11403_);
  and _84595_ (_34627_, _34626_, _34621_);
  nor _84596_ (_34628_, _05852_, _11330_);
  or _84597_ (_34629_, _34628_, _11331_);
  and _84598_ (_34630_, _34629_, _03775_);
  or _84599_ (_34631_, _34630_, _03179_);
  or _84600_ (_34632_, _34631_, _34627_);
  or _84601_ (_34634_, _34542_, _06328_);
  and _84602_ (_34635_, _34634_, _34632_);
  or _84603_ (_34636_, _34635_, _03522_);
  or _84604_ (_34637_, _34629_, _03523_);
  and _84605_ (_34638_, _34637_, _04192_);
  and _84606_ (_34639_, _34638_, _34636_);
  and _84607_ (_34640_, _34532_, _03790_);
  or _84608_ (_34641_, _34640_, _04947_);
  or _84609_ (_34642_, _34641_, _34639_);
  or _84610_ (_34643_, _34542_, _04533_);
  and _84611_ (_34645_, _34643_, _03521_);
  and _84612_ (_34646_, _34645_, _34642_);
  and _84613_ (_34647_, _12893_, _05269_);
  or _84614_ (_34648_, _34647_, _34527_);
  and _84615_ (_34649_, _34648_, _03520_);
  or _84616_ (_34650_, _34649_, _42967_);
  or _84617_ (_34651_, _34650_, _34646_);
  or _84618_ (_34652_, _42963_, \oc8051_golden_model_1.SP [4]);
  and _84619_ (_34653_, _34652_, _41755_);
  and _84620_ (_43383_, _34653_, _34651_);
  nor _84621_ (_34655_, _05269_, _11329_);
  and _84622_ (_34656_, _13042_, _05269_);
  or _84623_ (_34657_, _34656_, _34655_);
  and _84624_ (_34658_, _34657_, _03769_);
  nor _84625_ (_34659_, _12930_, _11355_);
  or _84626_ (_34660_, _34659_, _34655_);
  or _84627_ (_34661_, _34660_, _04444_);
  and _84628_ (_34662_, _05269_, \oc8051_golden_model_1.ACC [5]);
  or _84629_ (_34663_, _34662_, _34655_);
  or _84630_ (_34664_, _34663_, _04427_);
  or _84631_ (_34666_, _04426_, \oc8051_golden_model_1.SP [5]);
  and _84632_ (_34667_, _34666_, _04762_);
  and _84633_ (_34668_, _34667_, _34664_);
  nor _84634_ (_34669_, _11300_, \oc8051_golden_model_1.SP [5]);
  nor _84635_ (_34670_, _34669_, _11301_);
  and _84636_ (_34671_, _34670_, _03923_);
  or _84637_ (_34672_, _34671_, _03570_);
  or _84638_ (_34673_, _34672_, _34668_);
  and _84639_ (_34674_, _34673_, _03203_);
  and _84640_ (_34675_, _34674_, _34661_);
  and _84641_ (_34677_, _34670_, _04746_);
  or _84642_ (_34678_, _34677_, _03568_);
  or _84643_ (_34679_, _34678_, _34675_);
  and _84644_ (_34680_, _11332_, _03502_);
  nor _84645_ (_34681_, _34552_, _11329_);
  nor _84646_ (_34682_, _34681_, _34680_);
  nand _84647_ (_34683_, _34682_, _03568_);
  and _84648_ (_34684_, _34683_, _34679_);
  or _84649_ (_34685_, _34684_, _03575_);
  or _84650_ (_34686_, _34663_, _03583_);
  and _84651_ (_34688_, _34686_, _04887_);
  and _84652_ (_34689_, _34688_, _34685_);
  nor _84653_ (_34690_, _34562_, \oc8051_golden_model_1.SP [5]);
  nor _84654_ (_34691_, _34690_, _11344_);
  and _84655_ (_34692_, _34691_, _03511_);
  or _84656_ (_34693_, _34692_, _04744_);
  or _84657_ (_34694_, _34693_, _34689_);
  or _84658_ (_34695_, _34670_, _04745_);
  and _84659_ (_34696_, _34695_, _06039_);
  and _84660_ (_34697_, _34696_, _34694_);
  nor _84661_ (_34699_, _05422_, _11355_);
  or _84662_ (_34700_, _34699_, _34655_);
  and _84663_ (_34701_, _34700_, _07314_);
  or _84664_ (_34702_, _34701_, _03479_);
  or _84665_ (_34703_, _34702_, _34697_);
  and _84666_ (_34704_, _06721_, _05269_);
  or _84667_ (_34705_, _34655_, _06044_);
  or _84668_ (_34706_, _34705_, _34704_);
  and _84669_ (_34707_, _34706_, _03474_);
  and _84670_ (_34708_, _34707_, _34703_);
  nor _84671_ (_34710_, _13021_, _11355_);
  or _84672_ (_34711_, _34710_, _34655_);
  and _84673_ (_34712_, _34711_, _03221_);
  or _84674_ (_34713_, _34712_, _03437_);
  or _84675_ (_34714_, _34713_, _34708_);
  and _84676_ (_34715_, _06211_, _05269_);
  or _84677_ (_34716_, _34715_, _34655_);
  or _84678_ (_34717_, _34716_, _03438_);
  and _84679_ (_34718_, _34717_, _34714_);
  or _84680_ (_34719_, _34718_, _03189_);
  or _84681_ (_34721_, _34670_, _11376_);
  and _84682_ (_34722_, _34721_, _34719_);
  or _84683_ (_34723_, _34722_, _03636_);
  and _84684_ (_34724_, _13036_, _05269_);
  or _84685_ (_34725_, _34724_, _34655_);
  or _84686_ (_34726_, _34725_, _04499_);
  and _84687_ (_34727_, _34726_, _04501_);
  and _84688_ (_34728_, _34727_, _34723_);
  or _84689_ (_34729_, _34728_, _34658_);
  and _84690_ (_34730_, _34729_, _05769_);
  or _84691_ (_34732_, _34655_, _05472_);
  and _84692_ (_34733_, _34732_, _03754_);
  and _84693_ (_34734_, _34733_, _34716_);
  or _84694_ (_34735_, _34734_, _34730_);
  and _84695_ (_34736_, _34735_, _09960_);
  and _84696_ (_34737_, _34663_, _03752_);
  and _84697_ (_34738_, _34737_, _34732_);
  and _84698_ (_34739_, _34670_, _03192_);
  or _84699_ (_34740_, _34739_, _03758_);
  or _84700_ (_34741_, _34740_, _34738_);
  or _84701_ (_34743_, _34741_, _34736_);
  nor _84702_ (_34744_, _13035_, _11355_);
  or _84703_ (_34745_, _34744_, _34655_);
  or _84704_ (_34746_, _34745_, _03759_);
  and _84705_ (_34747_, _34746_, _34743_);
  or _84706_ (_34748_, _34747_, _03760_);
  nor _84707_ (_34749_, _13041_, _11355_);
  or _84708_ (_34750_, _34749_, _34655_);
  or _84709_ (_34751_, _34750_, _04517_);
  and _84710_ (_34752_, _34751_, _11403_);
  and _84711_ (_34754_, _34752_, _34748_);
  nor _84712_ (_34755_, _11331_, _11329_);
  or _84713_ (_34756_, _34755_, _11332_);
  and _84714_ (_34757_, _34756_, _03775_);
  or _84715_ (_34758_, _34757_, _03179_);
  or _84716_ (_34759_, _34758_, _34754_);
  or _84717_ (_34760_, _34670_, _06328_);
  and _84718_ (_34761_, _34760_, _34759_);
  or _84719_ (_34762_, _34761_, _03522_);
  or _84720_ (_34763_, _34756_, _03523_);
  and _84721_ (_34765_, _34763_, _04192_);
  and _84722_ (_34766_, _34765_, _34762_);
  and _84723_ (_34767_, _34660_, _03790_);
  or _84724_ (_34768_, _34767_, _04947_);
  or _84725_ (_34769_, _34768_, _34766_);
  or _84726_ (_34770_, _34670_, _04533_);
  and _84727_ (_34771_, _34770_, _03521_);
  and _84728_ (_34772_, _34771_, _34769_);
  and _84729_ (_34773_, _13097_, _05269_);
  or _84730_ (_34774_, _34773_, _34655_);
  and _84731_ (_34776_, _34774_, _03520_);
  or _84732_ (_34777_, _34776_, _42967_);
  or _84733_ (_34778_, _34777_, _34772_);
  or _84734_ (_34779_, _42963_, \oc8051_golden_model_1.SP [5]);
  and _84735_ (_34780_, _34779_, _41755_);
  and _84736_ (_43384_, _34780_, _34778_);
  nor _84737_ (_34781_, _42963_, _11328_);
  nor _84738_ (_34782_, _05269_, _11328_);
  and _84739_ (_34783_, _13259_, _05269_);
  or _84740_ (_34784_, _34783_, _34782_);
  and _84741_ (_34785_, _34784_, _03769_);
  nor _84742_ (_34786_, _05327_, _11355_);
  or _84743_ (_34787_, _34782_, _06039_);
  or _84744_ (_34788_, _34787_, _34786_);
  nor _84745_ (_34789_, _13122_, _11355_);
  or _84746_ (_34790_, _34789_, _34782_);
  or _84747_ (_34791_, _34790_, _04444_);
  and _84748_ (_34792_, _05269_, \oc8051_golden_model_1.ACC [6]);
  or _84749_ (_34793_, _34792_, _34782_);
  or _84750_ (_34794_, _34793_, _04427_);
  or _84751_ (_34797_, _04426_, \oc8051_golden_model_1.SP [6]);
  and _84752_ (_34798_, _34797_, _04762_);
  and _84753_ (_34799_, _34798_, _34794_);
  nor _84754_ (_34800_, _11301_, \oc8051_golden_model_1.SP [6]);
  nor _84755_ (_34801_, _34800_, _11302_);
  and _84756_ (_34802_, _34801_, _03923_);
  or _84757_ (_34803_, _34802_, _03570_);
  or _84758_ (_34804_, _34803_, _34799_);
  and _84759_ (_34805_, _34804_, _03203_);
  and _84760_ (_34806_, _34805_, _34791_);
  and _84761_ (_34808_, _34801_, _04746_);
  or _84762_ (_34809_, _34808_, _03568_);
  or _84763_ (_34810_, _34809_, _34806_);
  nor _84764_ (_34811_, _34680_, _11328_);
  nor _84765_ (_34812_, _34811_, _11334_);
  nand _84766_ (_34813_, _34812_, _03568_);
  and _84767_ (_34814_, _34813_, _34810_);
  or _84768_ (_34815_, _34814_, _03575_);
  or _84769_ (_34816_, _34793_, _03583_);
  and _84770_ (_34817_, _34816_, _04887_);
  and _84771_ (_34819_, _34817_, _34815_);
  nor _84772_ (_34820_, _11344_, \oc8051_golden_model_1.SP [6]);
  nor _84773_ (_34821_, _34820_, _11345_);
  and _84774_ (_34822_, _34821_, _03511_);
  or _84775_ (_34823_, _34822_, _34819_);
  and _84776_ (_34824_, _34823_, _04745_);
  nand _84777_ (_34825_, _34801_, _04744_);
  nand _84778_ (_34826_, _34825_, _06039_);
  or _84779_ (_34827_, _34826_, _34824_);
  and _84780_ (_34828_, _34827_, _34788_);
  or _84781_ (_34830_, _34828_, _03479_);
  and _84782_ (_34831_, _06713_, _05269_);
  or _84783_ (_34832_, _34782_, _06044_);
  or _84784_ (_34833_, _34832_, _34831_);
  and _84785_ (_34834_, _34833_, _03474_);
  and _84786_ (_34835_, _34834_, _34830_);
  nor _84787_ (_34836_, _13237_, _11355_);
  or _84788_ (_34837_, _34836_, _34782_);
  and _84789_ (_34838_, _34837_, _03221_);
  or _84790_ (_34839_, _34838_, _03437_);
  or _84791_ (_34841_, _34839_, _34835_);
  and _84792_ (_34842_, _13244_, _05269_);
  or _84793_ (_34843_, _34842_, _34782_);
  or _84794_ (_34844_, _34843_, _03438_);
  and _84795_ (_34845_, _34844_, _34841_);
  or _84796_ (_34846_, _34845_, _03189_);
  or _84797_ (_34847_, _34801_, _11376_);
  and _84798_ (_34848_, _34847_, _34846_);
  or _84799_ (_34849_, _34848_, _03636_);
  and _84800_ (_34850_, _13253_, _05269_);
  or _84801_ (_34852_, _34850_, _34782_);
  or _84802_ (_34853_, _34852_, _04499_);
  and _84803_ (_34854_, _34853_, _04501_);
  and _84804_ (_34855_, _34854_, _34849_);
  or _84805_ (_34856_, _34855_, _34785_);
  and _84806_ (_34857_, _34856_, _05769_);
  or _84807_ (_34858_, _34782_, _05377_);
  and _84808_ (_34859_, _34858_, _03754_);
  and _84809_ (_34860_, _34859_, _34843_);
  or _84810_ (_34861_, _34860_, _34857_);
  and _84811_ (_34863_, _34861_, _09960_);
  and _84812_ (_34864_, _34793_, _03752_);
  and _84813_ (_34865_, _34864_, _34858_);
  and _84814_ (_34866_, _34801_, _03192_);
  or _84815_ (_34867_, _34866_, _03758_);
  or _84816_ (_34868_, _34867_, _34865_);
  or _84817_ (_34869_, _34868_, _34863_);
  nor _84818_ (_34870_, _13251_, _11355_);
  or _84819_ (_34871_, _34870_, _34782_);
  or _84820_ (_34872_, _34871_, _03759_);
  and _84821_ (_34874_, _34872_, _34869_);
  or _84822_ (_34875_, _34874_, _03760_);
  nor _84823_ (_34876_, _13258_, _11355_);
  or _84824_ (_34877_, _34782_, _04517_);
  or _84825_ (_34878_, _34877_, _34876_);
  and _84826_ (_34879_, _34878_, _11403_);
  and _84827_ (_34880_, _34879_, _34875_);
  nor _84828_ (_34881_, _11332_, _11328_);
  or _84829_ (_34882_, _34881_, _11333_);
  and _84830_ (_34883_, _34882_, _03775_);
  or _84831_ (_34885_, _34883_, _03179_);
  or _84832_ (_34886_, _34885_, _34880_);
  or _84833_ (_34887_, _34801_, _06328_);
  and _84834_ (_34888_, _34887_, _34886_);
  or _84835_ (_34889_, _34888_, _03522_);
  or _84836_ (_34890_, _34882_, _03523_);
  and _84837_ (_34891_, _34890_, _34889_);
  or _84838_ (_34892_, _34891_, _03790_);
  or _84839_ (_34893_, _34790_, _04192_);
  and _84840_ (_34894_, _34893_, _04533_);
  and _84841_ (_34896_, _34894_, _34892_);
  and _84842_ (_34897_, _34801_, _04947_);
  or _84843_ (_34898_, _34897_, _03520_);
  or _84844_ (_34899_, _34898_, _34896_);
  and _84845_ (_34900_, _13312_, _05269_);
  or _84846_ (_34901_, _34782_, _03521_);
  or _84847_ (_34902_, _34901_, _34900_);
  and _84848_ (_34903_, _34902_, _42963_);
  and _84849_ (_34904_, _34903_, _34899_);
  or _84850_ (_34905_, _34904_, _34781_);
  and _84851_ (_43385_, _34905_, _41755_);
  not _84852_ (_34907_, \oc8051_golden_model_1.PSW [0]);
  nor _84853_ (_34908_, _42963_, _34907_);
  nor _84854_ (_34909_, _07444_, _07443_);
  nor _84855_ (_34910_, _34909_, _07346_);
  and _84856_ (_34911_, _34909_, _07346_);
  nor _84857_ (_34912_, _34911_, _34910_);
  nor _84858_ (_34913_, _07364_, _07363_);
  nor _84859_ (_34914_, _34913_, _15368_);
  and _84860_ (_34915_, _34913_, _15368_);
  nor _84861_ (_34917_, _34915_, _34914_);
  and _84862_ (_34918_, _34917_, _34912_);
  nor _84863_ (_34919_, _34917_, _34912_);
  nor _84864_ (_34920_, _34919_, _34918_);
  or _84865_ (_34921_, _34920_, _05834_);
  nand _84866_ (_34922_, _34920_, _05834_);
  and _84867_ (_34923_, _34922_, _34921_);
  or _84868_ (_34924_, _34923_, _04533_);
  not _84869_ (_34925_, _15392_);
  nor _84870_ (_34926_, _15115_, _10375_);
  and _84871_ (_34928_, _15115_, _10375_);
  or _84872_ (_34929_, _34928_, _34926_);
  and _84873_ (_34930_, _34929_, _34925_);
  nor _84874_ (_34931_, _34929_, _34925_);
  nor _84875_ (_34932_, _34931_, _34930_);
  and _84876_ (_34933_, _34932_, _16018_);
  nor _84877_ (_34934_, _34932_, _16018_);
  nor _84878_ (_34935_, _34934_, _34933_);
  nor _84879_ (_34936_, _34935_, _16345_);
  and _84880_ (_34937_, _34935_, _16345_);
  or _84881_ (_34939_, _34937_, _34936_);
  nor _84882_ (_34940_, _34939_, _16696_);
  and _84883_ (_34941_, _34939_, _16696_);
  or _84884_ (_34942_, _34941_, _34940_);
  and _84885_ (_34943_, _34942_, _17033_);
  nor _84886_ (_34944_, _34942_, _17033_);
  nor _84887_ (_34945_, _34944_, _34943_);
  nor _84888_ (_34946_, _34945_, _08642_);
  and _84889_ (_34947_, _34945_, _08642_);
  or _84890_ (_34948_, _34947_, _34946_);
  or _84891_ (_34950_, _34948_, _03526_);
  and _84892_ (_34951_, _34950_, _08598_);
  and _84893_ (_34952_, _15340_, _14860_);
  nor _84894_ (_34953_, _15340_, _14860_);
  nor _84895_ (_34954_, _34953_, _34952_);
  nor _84896_ (_34955_, _34954_, _15664_);
  and _84897_ (_34956_, _34954_, _15664_);
  nor _84898_ (_34957_, _34956_, _34955_);
  and _84899_ (_34958_, _34957_, _15999_);
  nor _84900_ (_34959_, _34957_, _15999_);
  nor _84901_ (_34961_, _34959_, _34958_);
  nor _84902_ (_34962_, _34961_, _16326_);
  and _84903_ (_34963_, _34961_, _16326_);
  or _84904_ (_34964_, _34963_, _34962_);
  nor _84905_ (_34965_, _34964_, _16672_);
  and _84906_ (_34966_, _34964_, _16672_);
  or _84907_ (_34967_, _34966_, _34965_);
  and _84908_ (_34968_, _34967_, _17016_);
  nor _84909_ (_34969_, _34967_, _17016_);
  nor _84910_ (_34970_, _34969_, _34968_);
  and _84911_ (_34972_, _34970_, _08581_);
  nor _84912_ (_34973_, _34970_, _08581_);
  or _84913_ (_34974_, _34973_, _34972_);
  and _84914_ (_34975_, _34974_, _08523_);
  nor _84915_ (_34976_, _14863_, _07887_);
  nor _84916_ (_34977_, _15328_, _15050_);
  nor _84917_ (_34978_, _34977_, _34976_);
  nor _84918_ (_34979_, _34978_, _15651_);
  and _84919_ (_34980_, _34978_, _15651_);
  nor _84920_ (_34981_, _34980_, _34979_);
  and _84921_ (_34983_, _34981_, _15983_);
  nor _84922_ (_34984_, _34981_, _15983_);
  or _84923_ (_34985_, _34984_, _34983_);
  nor _84924_ (_34986_, _34985_, _16314_);
  and _84925_ (_34987_, _34985_, _16314_);
  or _84926_ (_34988_, _34987_, _34986_);
  nor _84927_ (_34989_, _34988_, _16392_);
  and _84928_ (_34990_, _34988_, _16392_);
  or _84929_ (_34991_, _34990_, _34989_);
  nor _84930_ (_34992_, _34991_, _17000_);
  and _84931_ (_34994_, _34991_, _17000_);
  or _84932_ (_34995_, _34994_, _34992_);
  nand _84933_ (_34996_, _34995_, _07907_);
  or _84934_ (_34997_, _34995_, _07907_);
  and _84935_ (_34998_, _34997_, _34996_);
  or _84936_ (_34999_, _34998_, _07828_);
  and _84937_ (_35000_, _34999_, _08490_);
  and _84938_ (_35001_, _03484_, _03182_);
  or _84939_ (_35002_, _07806_, _07803_);
  nand _84940_ (_35003_, _07806_, _07803_);
  and _84941_ (_35005_, _35003_, _35002_);
  nor _84942_ (_35006_, _07799_, _07798_);
  and _84943_ (_35007_, _07799_, _07798_);
  nor _84944_ (_35008_, _35007_, _35006_);
  not _84945_ (_35009_, _35008_);
  and _84946_ (_35010_, _35009_, _35005_);
  nor _84947_ (_35011_, _35009_, _35005_);
  nor _84948_ (_35012_, _35011_, _35010_);
  nor _84949_ (_35013_, _07792_, _07785_);
  and _84950_ (_35014_, _07792_, _07785_);
  nor _84951_ (_35016_, _35014_, _35013_);
  nor _84952_ (_35017_, _35016_, _07791_);
  and _84953_ (_35018_, _35016_, _07791_);
  nor _84954_ (_35019_, _35018_, _35017_);
  not _84955_ (_35020_, _35019_);
  nor _84956_ (_35021_, _35020_, _35012_);
  and _84957_ (_35022_, _35020_, _35012_);
  nor _84958_ (_35023_, _35022_, _35021_);
  nand _84959_ (_35024_, _35023_, _07782_);
  or _84960_ (_35025_, _35023_, _07782_);
  and _84961_ (_35027_, _35025_, _35024_);
  or _84962_ (_35028_, _35027_, _08435_);
  nor _84963_ (_35029_, _10472_, _03744_);
  and _84964_ (_35030_, _35029_, _29345_);
  or _84965_ (_35031_, _35030_, _34923_);
  or _84966_ (_35032_, _34923_, _29147_);
  or _84967_ (_35033_, _06719_, _06570_);
  nand _84968_ (_35034_, _35033_, _12057_);
  or _84969_ (_35035_, _35033_, _12057_);
  nand _84970_ (_35036_, _35035_, _35034_);
  nor _84971_ (_35038_, _06723_, _06662_);
  or _84972_ (_35039_, _06713_, _06004_);
  or _84973_ (_35040_, _06388_, _05935_);
  and _84974_ (_35041_, _35040_, _35039_);
  nand _84975_ (_35042_, _35041_, _35038_);
  or _84976_ (_35043_, _35041_, _35038_);
  nand _84977_ (_35044_, _35043_, _35042_);
  nand _84978_ (_35045_, _35044_, _35036_);
  or _84979_ (_35046_, _35044_, _35036_);
  and _84980_ (_35047_, _35046_, _35045_);
  or _84981_ (_35049_, _35047_, _03043_);
  and _84982_ (_35050_, _35049_, _04458_);
  nor _84983_ (_35051_, _06693_, _05824_);
  and _84984_ (_35052_, _35051_, _12065_);
  nor _84985_ (_35053_, _35051_, _12065_);
  or _84986_ (_35054_, _35053_, _35052_);
  nor _84987_ (_35055_, _06695_, _05822_);
  nor _84988_ (_35056_, _35055_, _06702_);
  and _84989_ (_35057_, _35055_, _06702_);
  nor _84990_ (_35058_, _35057_, _35056_);
  or _84991_ (_35060_, _35058_, _35054_);
  nand _84992_ (_35061_, _35058_, _35054_);
  and _84993_ (_35062_, _35061_, _35060_);
  and _84994_ (_35063_, _35062_, _07928_);
  or _84995_ (_35064_, _35047_, _07936_);
  and _84996_ (_35065_, _05831_, _03208_);
  or _84997_ (_35066_, _35062_, _10288_);
  nor _84998_ (_35067_, _27282_, _03924_);
  nand _84999_ (_35068_, _35067_, _34907_);
  or _85000_ (_35069_, _35067_, _34923_);
  and _85001_ (_35071_, _35069_, _35068_);
  or _85002_ (_35072_, _35071_, _07933_);
  and _85003_ (_35073_, _35072_, _35066_);
  or _85004_ (_35074_, _35073_, _07935_);
  and _85005_ (_35075_, _35074_, _35065_);
  and _85006_ (_35076_, _35075_, _35064_);
  and _85007_ (_35077_, _34923_, _05833_);
  or _85008_ (_35078_, _35077_, _04438_);
  or _85009_ (_35079_, _35078_, _35076_);
  nor _85010_ (_35080_, _34913_, \oc8051_golden_model_1.ACC [6]);
  and _85011_ (_35082_, _34913_, \oc8051_golden_model_1.ACC [6]);
  nor _85012_ (_35083_, _35082_, _35080_);
  nor _85013_ (_35084_, _35083_, \oc8051_golden_model_1.ACC [7]);
  and _85014_ (_35085_, _35083_, \oc8051_golden_model_1.ACC [7]);
  nor _85015_ (_35086_, _35085_, _35084_);
  not _85016_ (_35087_, _35086_);
  nor _85017_ (_35088_, _35087_, _35036_);
  and _85018_ (_35089_, _35087_, _35036_);
  or _85019_ (_35090_, _35089_, _35088_);
  or _85020_ (_35091_, _35090_, _05847_);
  and _85021_ (_35093_, _35091_, _04444_);
  and _85022_ (_35094_, _35093_, _35079_);
  not _85023_ (_35095_, _14903_);
  or _85024_ (_35096_, _15160_, _35095_);
  nand _85025_ (_35097_, _15160_, _35095_);
  and _85026_ (_35098_, _35097_, _35096_);
  nand _85027_ (_35099_, _35098_, _15424_);
  or _85028_ (_35100_, _35098_, _15424_);
  nand _85029_ (_35101_, _35100_, _35099_);
  nand _85030_ (_35102_, _35101_, _16464_);
  or _85031_ (_35104_, _35101_, _16464_);
  and _85032_ (_35105_, _35104_, _35102_);
  nor _85033_ (_35106_, _16112_, _15793_);
  and _85034_ (_35107_, _16112_, _15793_);
  nor _85035_ (_35108_, _35107_, _35106_);
  nand _85036_ (_35109_, _35108_, _35105_);
  or _85037_ (_35110_, _35108_, _35105_);
  nand _85038_ (_35111_, _35110_, _35109_);
  and _85039_ (_35112_, _35111_, _16798_);
  nor _85040_ (_35113_, _35111_, _16798_);
  or _85041_ (_35115_, _35113_, _35112_);
  and _85042_ (_35116_, _35115_, _07950_);
  nor _85043_ (_35117_, _35115_, _07950_);
  or _85044_ (_35118_, _35117_, _35116_);
  and _85045_ (_35119_, _35118_, _03570_);
  or _85046_ (_35120_, _35119_, _07948_);
  or _85047_ (_35121_, _35120_, _35094_);
  and _85048_ (_35122_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor _85049_ (_35123_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or _85050_ (_35124_, _35123_, _35122_);
  and _85051_ (_35126_, _35124_, _15166_);
  nor _85052_ (_35127_, _35124_, _15166_);
  nor _85053_ (_35128_, _35127_, _35126_);
  and _85054_ (_35129_, _16118_, _15800_);
  nor _85055_ (_35130_, _16118_, _15800_);
  nor _85056_ (_35131_, _35130_, _35129_);
  nor _85057_ (_35132_, _35131_, _35128_);
  and _85058_ (_35133_, _35131_, _35128_);
  or _85059_ (_35134_, _35133_, _35132_);
  nor _85060_ (_35135_, _35134_, _07972_);
  and _85061_ (_35137_, _35134_, _07972_);
  or _85062_ (_35138_, _35137_, _35135_);
  and _85063_ (_35139_, _35138_, _16470_);
  nor _85064_ (_35140_, _35138_, _16470_);
  or _85065_ (_35141_, _35140_, _35139_);
  nor _85066_ (_35142_, _35141_, _16806_);
  and _85067_ (_35143_, _35141_, _16806_);
  or _85068_ (_35144_, _35143_, _35142_);
  or _85069_ (_35145_, _35144_, _11538_);
  and _85070_ (_35146_, _35145_, _35121_);
  or _85071_ (_35148_, _35146_, _10254_);
  or _85072_ (_35149_, _34923_, _11551_);
  and _85073_ (_35150_, _35149_, _03517_);
  and _85074_ (_35151_, _35150_, _35148_);
  not _85075_ (_35152_, _07979_);
  and _85076_ (_35153_, _15173_, _14909_);
  nor _85077_ (_35154_, _15173_, _14909_);
  or _85078_ (_35155_, _35154_, _35153_);
  nor _85079_ (_35156_, _16813_, _16125_);
  and _85080_ (_35157_, _16813_, _16125_);
  nor _85081_ (_35159_, _35157_, _35156_);
  nor _85082_ (_35160_, _35159_, _35155_);
  and _85083_ (_35161_, _35159_, _35155_);
  or _85084_ (_35162_, _35161_, _35160_);
  not _85085_ (_35163_, _16475_);
  nor _85086_ (_35164_, _15805_, _15438_);
  and _85087_ (_35165_, _15805_, _15438_);
  nor _85088_ (_35166_, _35165_, _35164_);
  nor _85089_ (_35167_, _35166_, _35163_);
  and _85090_ (_35168_, _35166_, _35163_);
  nor _85091_ (_35170_, _35168_, _35167_);
  and _85092_ (_35171_, _35170_, _35162_);
  nor _85093_ (_35172_, _35170_, _35162_);
  nor _85094_ (_35173_, _35172_, _35171_);
  nand _85095_ (_35174_, _35173_, _35152_);
  or _85096_ (_35175_, _35173_, _35152_);
  and _85097_ (_35176_, _35175_, _03516_);
  and _85098_ (_35177_, _35176_, _35174_);
  or _85099_ (_35178_, _35177_, _28712_);
  or _85100_ (_35179_, _35178_, _35151_);
  not _85101_ (_35181_, _16756_);
  and _85102_ (_35182_, _35181_, _07920_);
  nor _85103_ (_35183_, _35181_, _07920_);
  nor _85104_ (_35184_, _35183_, _35182_);
  and _85105_ (_35185_, _15132_, _14885_);
  nor _85106_ (_35186_, _15132_, _14885_);
  nor _85107_ (_35187_, _35186_, _35185_);
  and _85108_ (_35188_, _35187_, _15407_);
  nor _85109_ (_35189_, _35187_, _15407_);
  or _85110_ (_35190_, _35189_, _35188_);
  and _85111_ (_35192_, _35190_, _15754_);
  nor _85112_ (_35193_, _35190_, _15754_);
  or _85113_ (_35194_, _35193_, _35192_);
  not _85114_ (_35195_, _16410_);
  and _85115_ (_35196_, _35195_, _16084_);
  nor _85116_ (_35197_, _35195_, _16084_);
  nor _85117_ (_35198_, _35197_, _35196_);
  and _85118_ (_35199_, _35198_, _35194_);
  nor _85119_ (_35200_, _35198_, _35194_);
  nor _85120_ (_35201_, _35200_, _35199_);
  or _85121_ (_35203_, _35201_, _35184_);
  nand _85122_ (_35204_, _35201_, _35184_);
  and _85123_ (_35205_, _35204_, _35203_);
  or _85124_ (_35206_, _35205_, _03983_);
  or _85125_ (_35207_, _34923_, _03203_);
  and _85126_ (_35208_, _35207_, _07927_);
  and _85127_ (_35209_, _35208_, _35206_);
  and _85128_ (_35210_, _35209_, _35179_);
  or _85129_ (_35211_, _35210_, _35063_);
  and _85130_ (_35212_, _35211_, _07987_);
  or _85131_ (_35214_, _35212_, _35050_);
  not _85132_ (_35215_, _04004_);
  or _85133_ (_35216_, _35047_, _35215_);
  and _85134_ (_35217_, _35216_, _04718_);
  or _85135_ (_35218_, _35217_, _03205_);
  and _85136_ (_35219_, _35218_, _35214_);
  and _85137_ (_35220_, _08222_, _08205_);
  nor _85138_ (_35221_, _35220_, _08223_);
  and _85139_ (_35222_, _35221_, _08143_);
  nor _85140_ (_35223_, _35221_, _08143_);
  nor _85141_ (_35225_, _35223_, _35222_);
  and _85142_ (_35226_, _08178_, _08163_);
  and _85143_ (_35227_, _08177_, _08164_);
  nor _85144_ (_35228_, _35227_, _35226_);
  and _85145_ (_35229_, _08191_, _08125_);
  nor _85146_ (_35230_, _08191_, _08125_);
  or _85147_ (_35231_, _35230_, _35229_);
  and _85148_ (_35232_, _35231_, _35228_);
  nor _85149_ (_35233_, _35231_, _35228_);
  or _85150_ (_35234_, _35233_, _35232_);
  nor _85151_ (_35236_, _35234_, _35225_);
  and _85152_ (_35237_, _35234_, _35225_);
  nor _85153_ (_35238_, _35237_, _35236_);
  nand _85154_ (_35239_, _35238_, _11721_);
  or _85155_ (_35240_, _35238_, _11721_);
  and _85156_ (_35241_, _35240_, _03575_);
  and _85157_ (_35242_, _35241_, _35239_);
  or _85158_ (_35243_, _35242_, _26220_);
  or _85159_ (_35244_, _35243_, _35219_);
  or _85160_ (_35245_, _34923_, _10316_);
  and _85161_ (_35247_, _35245_, _03513_);
  and _85162_ (_35248_, _35247_, _35244_);
  not _85163_ (_35249_, _15456_);
  nor _85164_ (_35250_, _15191_, _14873_);
  and _85165_ (_35251_, _15191_, _14873_);
  nor _85166_ (_35252_, _35251_, _35250_);
  nor _85167_ (_35253_, _35252_, _35249_);
  and _85168_ (_35254_, _35252_, _35249_);
  or _85169_ (_35255_, _35254_, _35253_);
  and _85170_ (_35256_, _35255_, _15826_);
  nor _85171_ (_35258_, _35255_, _15826_);
  or _85172_ (_35259_, _35258_, _35256_);
  and _85173_ (_35260_, _35259_, _16145_);
  nor _85174_ (_35261_, _35259_, _16145_);
  or _85175_ (_35262_, _35261_, _35260_);
  and _85176_ (_35263_, _35262_, _16495_);
  nor _85177_ (_35264_, _35262_, _16495_);
  or _85178_ (_35265_, _35264_, _35263_);
  and _85179_ (_35266_, _35265_, _16832_);
  nor _85180_ (_35267_, _35265_, _16832_);
  or _85181_ (_35269_, _35267_, _35266_);
  and _85182_ (_35270_, _35269_, _07999_);
  nor _85183_ (_35271_, _35269_, _07999_);
  or _85184_ (_35272_, _35271_, _35270_);
  nand _85185_ (_35273_, _35272_, _03512_);
  nor _85186_ (_35274_, _03962_, _03929_);
  and _85187_ (_35275_, _35274_, _10250_);
  nand _85188_ (_35276_, _35275_, _35273_);
  or _85189_ (_35277_, _35276_, _35248_);
  and _85190_ (_35278_, _03661_, _03504_);
  nor _85191_ (_35280_, _35275_, _34923_);
  nor _85192_ (_35281_, _35280_, _35278_);
  and _85193_ (_35282_, _35281_, _35277_);
  nand _85194_ (_35283_, _34923_, _35278_);
  nor _85195_ (_35284_, _09947_, _03199_);
  nor _85196_ (_35285_, _35284_, _29019_);
  nand _85197_ (_35286_, _35285_, _35283_);
  or _85198_ (_35287_, _35286_, _35282_);
  or _85199_ (_35288_, _35285_, _34923_);
  and _85200_ (_35289_, _35288_, _03506_);
  and _85201_ (_35291_, _35289_, _35287_);
  nor _85202_ (_35292_, _15773_, _35095_);
  and _85203_ (_35293_, _15773_, _35095_);
  nor _85204_ (_35294_, _35293_, _35292_);
  nor _85205_ (_35295_, _35294_, _16150_);
  and _85206_ (_35296_, _35294_, _16150_);
  or _85207_ (_35297_, _35296_, _35295_);
  not _85208_ (_35298_, _15461_);
  and _85209_ (_35299_, _35298_, _15196_);
  nor _85210_ (_35300_, _35298_, _15196_);
  nor _85211_ (_35302_, _35300_, _35299_);
  nor _85212_ (_35303_, _35302_, _16447_);
  and _85213_ (_35304_, _35302_, _16447_);
  nor _85214_ (_35305_, _35304_, _35303_);
  and _85215_ (_35306_, _35305_, _35297_);
  nor _85216_ (_35307_, _35305_, _35297_);
  nor _85217_ (_35308_, _35307_, _35306_);
  not _85218_ (_35309_, _16838_);
  and _85219_ (_35310_, _35309_, _08004_);
  nor _85220_ (_35311_, _35309_, _08004_);
  nor _85221_ (_35313_, _35311_, _35310_);
  nand _85222_ (_35314_, _35313_, _35308_);
  or _85223_ (_35315_, _35313_, _35308_);
  and _85224_ (_35316_, _35315_, _03505_);
  nand _85225_ (_35317_, _35316_, _35314_);
  nor _85226_ (_35318_, _26278_, _04743_);
  and _85227_ (_35319_, _35318_, _26277_);
  nand _85228_ (_35320_, _35319_, _35317_);
  or _85229_ (_35321_, _35320_, _35291_);
  or _85230_ (_35322_, _35319_, _34923_);
  and _85231_ (_35324_, _35322_, _26275_);
  and _85232_ (_35325_, _35324_, _35321_);
  nor _85233_ (_35326_, _10412_, _04478_);
  not _85234_ (_35327_, _26275_);
  nand _85235_ (_35328_, _34923_, _35327_);
  nand _85236_ (_35329_, _35328_, _35326_);
  or _85237_ (_35330_, _35329_, _35325_);
  or _85238_ (_35331_, _35326_, _34923_);
  and _85239_ (_35332_, _35331_, _06800_);
  and _85240_ (_35333_, _35332_, _35330_);
  nor _85241_ (_35335_, _03607_, _10420_);
  nand _85242_ (_35336_, _35335_, _09771_);
  nor _85243_ (_35337_, _15202_, _14934_);
  and _85244_ (_35338_, _15202_, _14934_);
  or _85245_ (_35339_, _35338_, _35337_);
  nor _85246_ (_35340_, _35339_, _15466_);
  and _85247_ (_35341_, _35339_, _15466_);
  nor _85248_ (_35342_, _35341_, _35340_);
  nor _85249_ (_35343_, _35342_, _15833_);
  and _85250_ (_35344_, _35342_, _15833_);
  nor _85251_ (_35346_, _35344_, _35343_);
  not _85252_ (_35347_, _35346_);
  nor _85253_ (_35348_, _35347_, _16156_);
  and _85254_ (_35349_, _35347_, _16156_);
  nor _85255_ (_35350_, _35349_, _35348_);
  nor _85256_ (_35351_, _35350_, _16502_);
  and _85257_ (_35352_, _35350_, _16502_);
  or _85258_ (_35353_, _35352_, _35351_);
  and _85259_ (_35354_, _35353_, _16843_);
  nor _85260_ (_35355_, _35353_, _16843_);
  nor _85261_ (_35357_, _35355_, _35354_);
  or _85262_ (_35358_, _35357_, _08009_);
  nand _85263_ (_35359_, _35357_, _08009_);
  and _85264_ (_35360_, _35359_, _06794_);
  and _85265_ (_35361_, _35360_, _35358_);
  or _85266_ (_35362_, _35361_, _35336_);
  or _85267_ (_35363_, _35362_, _35333_);
  not _85268_ (_35364_, _35336_);
  or _85269_ (_35365_, _35364_, _34923_);
  and _85270_ (_35366_, _35365_, _11467_);
  and _85271_ (_35368_, _35366_, _35363_);
  and _85272_ (_35369_, _34923_, _03606_);
  or _85273_ (_35370_, _35369_, _07923_);
  or _85274_ (_35371_, _35370_, _35368_);
  nor _85275_ (_35372_, _15210_, _14863_);
  and _85276_ (_35373_, _15210_, _14863_);
  or _85277_ (_35374_, _35373_, _35372_);
  and _85278_ (_35375_, _35374_, _15484_);
  nor _85279_ (_35376_, _35374_, _15484_);
  or _85280_ (_35377_, _35376_, _35375_);
  and _85281_ (_35379_, _35377_, _15849_);
  nor _85282_ (_35380_, _35377_, _15849_);
  or _85283_ (_35381_, _35380_, _35379_);
  or _85284_ (_35382_, _35381_, _16174_);
  nand _85285_ (_35383_, _35381_, _16174_);
  and _85286_ (_35384_, _35383_, _35382_);
  nor _85287_ (_35385_, _35384_, _16442_);
  and _85288_ (_35386_, _35384_, _16442_);
  or _85289_ (_35387_, _35386_, _35385_);
  nor _85290_ (_35388_, _35387_, _16860_);
  and _85291_ (_35390_, _35387_, _16860_);
  nor _85292_ (_35391_, _35390_, _35388_);
  or _85293_ (_35392_, _35391_, _08033_);
  and _85294_ (_35393_, _08032_, _07923_);
  nand _85295_ (_35394_, _35393_, _35391_);
  and _85296_ (_35395_, _35394_, _08037_);
  and _85297_ (_35396_, _35395_, _35392_);
  and _85298_ (_35397_, _35396_, _35371_);
  not _85299_ (_35398_, _16193_);
  or _85300_ (_35399_, _15141_, _14943_);
  nand _85301_ (_35401_, _15141_, _14943_);
  and _85302_ (_35402_, _35401_, _35399_);
  nor _85303_ (_35403_, _35402_, _15503_);
  and _85304_ (_35404_, _35402_, _15503_);
  nor _85305_ (_35405_, _35404_, _35403_);
  and _85306_ (_35406_, _35405_, _15867_);
  nor _85307_ (_35407_, _35405_, _15867_);
  or _85308_ (_35408_, _35407_, _35406_);
  nand _85309_ (_35409_, _35408_, _35398_);
  or _85310_ (_35410_, _35408_, _35398_);
  and _85311_ (_35412_, _35410_, _35409_);
  or _85312_ (_35413_, _35412_, _16522_);
  nand _85313_ (_35414_, _35412_, _16522_);
  and _85314_ (_35415_, _35414_, _35413_);
  nor _85315_ (_35416_, _35415_, _16783_);
  and _85316_ (_35417_, _35415_, _16783_);
  nor _85317_ (_35418_, _35417_, _35416_);
  not _85318_ (_35419_, _35418_);
  nand _85319_ (_35420_, _35419_, _08104_);
  or _85320_ (_35421_, _35419_, _08104_);
  and _85321_ (_35423_, _35421_, _08035_);
  and _85322_ (_35424_, _35423_, _35420_);
  or _85323_ (_35425_, _35424_, _03614_);
  or _85324_ (_35426_, _35425_, _35397_);
  nand _85325_ (_35427_, _15220_, _14948_);
  or _85326_ (_35428_, _15220_, _14948_);
  and _85327_ (_35429_, _35428_, _35427_);
  and _85328_ (_35430_, _35429_, _15517_);
  nor _85329_ (_35431_, _35429_, _15517_);
  or _85330_ (_35432_, _35431_, _35430_);
  nor _85331_ (_35434_, _35432_, _15880_);
  and _85332_ (_35435_, _35432_, _15880_);
  or _85333_ (_35436_, _35435_, _35434_);
  and _85334_ (_35437_, _35436_, _16095_);
  nor _85335_ (_35438_, _35436_, _16095_);
  or _85336_ (_35439_, _35438_, _35437_);
  nor _85337_ (_35440_, _35439_, _16534_);
  and _85338_ (_35441_, _35439_, _16534_);
  or _85339_ (_35442_, _35441_, _35440_);
  nor _85340_ (_35443_, _35442_, _16767_);
  and _85341_ (_35445_, _35442_, _16767_);
  or _85342_ (_35446_, _35445_, _35443_);
  nor _85343_ (_35447_, _35446_, _08284_);
  and _85344_ (_35448_, _35446_, _08284_);
  or _85345_ (_35449_, _35448_, _35447_);
  or _85346_ (_35450_, _35449_, _03619_);
  and _85347_ (_35451_, _35450_, _08109_);
  and _85348_ (_35452_, _35451_, _35426_);
  nand _85349_ (_35453_, _15228_, _14860_);
  or _85350_ (_35454_, _15228_, _14860_);
  and _85351_ (_35456_, _35454_, _35453_);
  nand _85352_ (_35457_, _35456_, _15535_);
  or _85353_ (_35458_, _35456_, _15535_);
  and _85354_ (_35459_, _35458_, _35457_);
  nor _85355_ (_35460_, _35459_, _15767_);
  and _85356_ (_35461_, _35459_, _15767_);
  or _85357_ (_35462_, _35461_, _35460_);
  and _85358_ (_35463_, _16425_, _16211_);
  nor _85359_ (_35464_, _16425_, _16211_);
  or _85360_ (_35465_, _35464_, _35463_);
  and _85361_ (_35467_, _35465_, _35462_);
  nor _85362_ (_35468_, _35465_, _35462_);
  nor _85363_ (_35469_, _35468_, _35467_);
  nor _85364_ (_35470_, _35469_, _16877_);
  and _85365_ (_35471_, _35469_, _16877_);
  nor _85366_ (_35472_, _35471_, _35470_);
  nor _85367_ (_35473_, _35472_, _08351_);
  and _85368_ (_35474_, _35472_, _08351_);
  or _85369_ (_35475_, _35474_, _35473_);
  and _85370_ (_35476_, _35475_, _08108_);
  or _85371_ (_35478_, _35476_, _03311_);
  or _85372_ (_35479_, _35478_, _35452_);
  nor _85373_ (_35480_, _05181_, _03562_);
  nor _85374_ (_35481_, _05191_, _05183_);
  nor _85375_ (_35482_, _05232_, _05196_);
  nor _85376_ (_35483_, _05187_, _05206_);
  nor _85377_ (_35484_, _35483_, _35482_);
  and _85378_ (_35485_, _35483_, _35482_);
  nor _85379_ (_35486_, _35485_, _35484_);
  nor _85380_ (_35487_, _35486_, _35481_);
  and _85381_ (_35489_, _35486_, _35481_);
  nor _85382_ (_35490_, _35489_, _35487_);
  not _85383_ (_35491_, _35490_);
  nor _85384_ (_35492_, _35491_, _35480_);
  and _85385_ (_35493_, _35491_, _35480_);
  or _85386_ (_35494_, _35493_, _35492_);
  or _85387_ (_35495_, _35494_, _03254_);
  and _85388_ (_35496_, _35495_, _03500_);
  and _85389_ (_35497_, _35496_, _35479_);
  not _85390_ (_35498_, _15891_);
  and _85391_ (_35500_, _35498_, _15544_);
  nor _85392_ (_35501_, _35498_, _15544_);
  nor _85393_ (_35502_, _35501_, _35500_);
  nor _85394_ (_35503_, _16545_, _16220_);
  and _85395_ (_35504_, _16545_, _16220_);
  nor _85396_ (_35505_, _35504_, _35503_);
  nor _85397_ (_35506_, _35505_, _35502_);
  and _85398_ (_35507_, _35505_, _35502_);
  nor _85399_ (_35508_, _35507_, _35506_);
  and _85400_ (_35509_, _15236_, _14958_);
  nor _85401_ (_35512_, _15236_, _14958_);
  nor _85402_ (_35513_, _35512_, _35509_);
  and _85403_ (_35514_, _16886_, _08360_);
  nor _85404_ (_35515_, _16886_, _08360_);
  nor _85405_ (_35516_, _35515_, _35514_);
  not _85406_ (_35517_, _35516_);
  and _85407_ (_35518_, _35517_, _35513_);
  nor _85408_ (_35519_, _35517_, _35513_);
  nor _85409_ (_35520_, _35519_, _35518_);
  nand _85410_ (_35521_, _35520_, _35508_);
  or _85411_ (_35523_, _35520_, _35508_);
  and _85412_ (_35524_, _35523_, _03499_);
  and _85413_ (_35525_, _35524_, _35521_);
  or _85414_ (_35526_, _35525_, _29148_);
  or _85415_ (_35527_, _35526_, _35497_);
  nand _85416_ (_35528_, _35527_, _35032_);
  and _85417_ (_35529_, _03664_, _03186_);
  not _85418_ (_35530_, _35529_);
  and _85419_ (_35531_, _35530_, _03492_);
  nand _85420_ (_35532_, _35531_, _35528_);
  nor _85421_ (_35535_, _35531_, _35205_);
  nor _85422_ (_35536_, _35535_, _04070_);
  and _85423_ (_35537_, _35536_, _35532_);
  and _85424_ (_35538_, _35205_, _04070_);
  or _85425_ (_35539_, _35538_, _03479_);
  or _85426_ (_35540_, _35539_, _35537_);
  not _85427_ (_35541_, _16894_);
  and _85428_ (_35542_, _35541_, _08367_);
  nor _85429_ (_35543_, _35541_, _08367_);
  nor _85430_ (_35544_, _35543_, _35542_);
  not _85431_ (_35546_, _16553_);
  and _85432_ (_35547_, _35546_, _16227_);
  nor _85433_ (_35548_, _35546_, _16227_);
  nor _85434_ (_35549_, _35548_, _35547_);
  and _85435_ (_35550_, _15243_, _14965_);
  nor _85436_ (_35551_, _15243_, _14965_);
  nor _85437_ (_35552_, _35551_, _35550_);
  not _85438_ (_35553_, _35552_);
  not _85439_ (_35554_, _15898_);
  and _85440_ (_35555_, _35554_, _15552_);
  nor _85441_ (_35558_, _35554_, _15552_);
  nor _85442_ (_35559_, _35558_, _35555_);
  and _85443_ (_35560_, _35559_, _35553_);
  nor _85444_ (_35561_, _35559_, _35553_);
  nor _85445_ (_35562_, _35561_, _35560_);
  nor _85446_ (_35563_, _35562_, _35549_);
  and _85447_ (_35564_, _35562_, _35549_);
  nor _85448_ (_35565_, _35564_, _35563_);
  or _85449_ (_35566_, _35565_, _35544_);
  nand _85450_ (_35567_, _35565_, _35544_);
  and _85451_ (_35569_, _35567_, _35566_);
  or _85452_ (_35570_, _35569_, _06044_);
  and _85453_ (_35571_, _35570_, _03474_);
  and _85454_ (_35572_, _35571_, _35540_);
  not _85455_ (_35573_, _16899_);
  and _85456_ (_35574_, _35573_, _08372_);
  nor _85457_ (_35575_, _35573_, _08372_);
  nor _85458_ (_35576_, _35575_, _35574_);
  not _85459_ (_35577_, _16558_);
  and _85460_ (_35578_, _35577_, _16233_);
  nor _85461_ (_35581_, _35577_, _16233_);
  nor _85462_ (_35582_, _35581_, _35578_);
  not _85463_ (_35583_, _35582_);
  and _85464_ (_35584_, _15248_, _14882_);
  nor _85465_ (_35585_, _15248_, _14882_);
  nor _85466_ (_35586_, _35585_, _35584_);
  not _85467_ (_35587_, _15904_);
  and _85468_ (_35588_, _35587_, _15557_);
  nor _85469_ (_35589_, _35587_, _15557_);
  nor _85470_ (_35590_, _35589_, _35588_);
  nor _85471_ (_35592_, _35590_, _35586_);
  and _85472_ (_35593_, _35590_, _35586_);
  nor _85473_ (_35594_, _35593_, _35592_);
  nor _85474_ (_35595_, _35594_, _35583_);
  and _85475_ (_35596_, _35594_, _35583_);
  nor _85476_ (_35597_, _35596_, _35595_);
  nand _85477_ (_35598_, _35597_, _35576_);
  or _85478_ (_35599_, _35597_, _35576_);
  and _85479_ (_35600_, _35599_, _03221_);
  and _85480_ (_35601_, _35600_, _35598_);
  or _85481_ (_35603_, _35601_, _35572_);
  and _85482_ (_35604_, _35603_, _07677_);
  nor _85483_ (_35605_, _07520_, _07466_);
  and _85484_ (_35606_, _07520_, _07466_);
  nor _85485_ (_35607_, _35606_, _35605_);
  nor _85486_ (_35608_, _35607_, _07412_);
  and _85487_ (_35609_, _35607_, _07412_);
  nor _85488_ (_35610_, _35609_, _35608_);
  and _85489_ (_35611_, _35610_, _16905_);
  nor _85490_ (_35612_, _35610_, _16905_);
  nor _85491_ (_35614_, _35612_, _35611_);
  and _85492_ (_35615_, _07382_, _08379_);
  nor _85493_ (_35616_, _07382_, _08379_);
  nor _85494_ (_35617_, _35616_, _35615_);
  and _85495_ (_35618_, _35617_, _35614_);
  nor _85496_ (_35619_, _35617_, _35614_);
  or _85497_ (_35620_, _35619_, _35618_);
  and _85498_ (_35621_, _35620_, _07596_);
  nor _85499_ (_35622_, _35620_, _07596_);
  nor _85500_ (_35623_, _35622_, _35621_);
  and _85501_ (_35625_, _35623_, _07675_);
  nor _85502_ (_35626_, _35623_, _07675_);
  or _85503_ (_35627_, _35626_, _35625_);
  and _85504_ (_35628_, _35627_, _07328_);
  or _85505_ (_35629_, _35628_, _03231_);
  or _85506_ (_35630_, _35629_, _35604_);
  or _85507_ (_35631_, _35494_, _03232_);
  and _85508_ (_35632_, _35631_, _27421_);
  and _85509_ (_35633_, _35632_, _35630_);
  nand _85510_ (_35634_, _34923_, _03745_);
  nor _85511_ (_35636_, _28687_, _04739_);
  nor _85512_ (_35637_, _03483_, _03633_);
  or _85513_ (_35638_, _35637_, _04657_);
  and _85514_ (_35639_, _35638_, _35636_);
  nand _85515_ (_35640_, _35639_, _35634_);
  or _85516_ (_35641_, _35640_, _35633_);
  and _85517_ (_35642_, _03487_, _03188_);
  nor _85518_ (_35643_, _35639_, _34923_);
  nor _85519_ (_35644_, _35643_, _35642_);
  and _85520_ (_35645_, _35644_, _35641_);
  nand _85521_ (_35647_, _34923_, _35642_);
  nand _85522_ (_35648_, _35647_, _04731_);
  or _85523_ (_35649_, _35648_, _35645_);
  nor _85524_ (_35650_, _34923_, _04731_);
  nor _85525_ (_35651_, _35650_, _04758_);
  and _85526_ (_35652_, _35651_, _35649_);
  or _85527_ (_35653_, _04489_, _04758_);
  or _85528_ (_35654_, _34923_, _04489_);
  and _85529_ (_35655_, _35654_, _35653_);
  or _85530_ (_35656_, _35655_, _35652_);
  or _85531_ (_35658_, _34923_, _04910_);
  and _85532_ (_35659_, _35658_, _03438_);
  and _85533_ (_35660_, _35659_, _35656_);
  nor _85534_ (_35661_, _15258_, _14976_);
  and _85535_ (_35662_, _15258_, _14976_);
  or _85536_ (_35663_, _35662_, _35661_);
  nor _85537_ (_35664_, _15915_, _15568_);
  and _85538_ (_35665_, _15915_, _15568_);
  nor _85539_ (_35666_, _35665_, _35664_);
  nor _85540_ (_35667_, _35666_, _35663_);
  and _85541_ (_35669_, _35666_, _35663_);
  or _85542_ (_35670_, _35669_, _35667_);
  nor _85543_ (_35671_, _16569_, _16244_);
  and _85544_ (_35672_, _16569_, _16244_);
  nor _85545_ (_35673_, _35672_, _35671_);
  and _85546_ (_35674_, _35673_, _16913_);
  nor _85547_ (_35675_, _35673_, _16913_);
  nor _85548_ (_35676_, _35675_, _35674_);
  and _85549_ (_35677_, _35676_, _35670_);
  nor _85550_ (_35678_, _35676_, _35670_);
  or _85551_ (_35680_, _35678_, _35677_);
  or _85552_ (_35681_, _35680_, _08388_);
  nand _85553_ (_35682_, _35680_, _08388_);
  and _85554_ (_35683_, _35682_, _03437_);
  and _85555_ (_35684_, _35683_, _35681_);
  or _85556_ (_35685_, _35684_, _35660_);
  and _85557_ (_35686_, _35685_, _08386_);
  nand _85558_ (_35687_, _35494_, _08385_);
  nand _85559_ (_35688_, _35687_, _35030_);
  or _85560_ (_35689_, _35688_, _35686_);
  nand _85561_ (_35691_, _35689_, _35031_);
  nand _85562_ (_35692_, _35691_, _16251_);
  not _85563_ (_35693_, _04347_);
  nor _85564_ (_35694_, _16923_, _07784_);
  and _85565_ (_35695_, _16923_, _07784_);
  nor _85566_ (_35696_, _35695_, _35694_);
  and _85567_ (_35697_, _14983_, _07805_);
  nor _85568_ (_35698_, _35697_, _15477_);
  and _85569_ (_35699_, _15724_, _07801_);
  nor _85570_ (_35700_, _15724_, _07801_);
  nor _85571_ (_35702_, _35700_, _35699_);
  nor _85572_ (_35703_, _35702_, _35698_);
  and _85573_ (_35704_, _35702_, _35698_);
  nor _85574_ (_35705_, _35704_, _35703_);
  and _85575_ (_35706_, _16406_, _07794_);
  nor _85576_ (_35707_, _16406_, _07794_);
  nor _85577_ (_35708_, _35707_, _35706_);
  nor _85578_ (_35709_, _35708_, _35705_);
  and _85579_ (_35710_, _35708_, _35705_);
  nor _85580_ (_35711_, _35710_, _35709_);
  nor _85581_ (_35713_, _35711_, _35696_);
  and _85582_ (_35714_, _35711_, _35696_);
  or _85583_ (_35715_, _35714_, _35713_);
  or _85584_ (_35716_, _35715_, _16251_);
  and _85585_ (_35717_, _35716_, _35693_);
  and _85586_ (_35718_, _35717_, _35692_);
  and _85587_ (_35719_, _35715_, _04347_);
  or _85588_ (_35720_, _35719_, _15268_);
  or _85589_ (_35721_, _35720_, _35718_);
  or _85590_ (_35722_, _35715_, _14992_);
  and _85591_ (_35724_, _35722_, _15582_);
  and _85592_ (_35725_, _35724_, _35721_);
  and _85593_ (_35726_, _35715_, _04129_);
  or _85594_ (_35727_, _35726_, _08405_);
  or _85595_ (_35728_, _35727_, _35725_);
  and _85596_ (_35729_, _15748_, _07752_);
  nor _85597_ (_35730_, _15748_, _07752_);
  nor _85598_ (_35731_, _35730_, _35729_);
  and _85599_ (_35732_, _14878_, _07756_);
  nor _85600_ (_35733_, _35732_, _15495_);
  nor _85601_ (_35735_, _35733_, _35731_);
  and _85602_ (_35736_, _35733_, _35731_);
  nor _85603_ (_35737_, _35736_, _35735_);
  and _85604_ (_35738_, _07745_, _07741_);
  nor _85605_ (_35739_, _07745_, _07741_);
  nor _85606_ (_35740_, _35739_, _35738_);
  nor _85607_ (_35741_, _35740_, _35737_);
  and _85608_ (_35742_, _35740_, _35737_);
  nor _85609_ (_35743_, _35742_, _35741_);
  nand _85610_ (_35744_, _07738_, _07735_);
  or _85611_ (_35746_, _07738_, _07735_);
  and _85612_ (_35747_, _35746_, _35744_);
  nand _85613_ (_35748_, _35747_, _35743_);
  or _85614_ (_35749_, _35747_, _35743_);
  and _85615_ (_35750_, _35749_, _35748_);
  or _85616_ (_35751_, _35750_, _08406_);
  and _85617_ (_35752_, _35751_, _03768_);
  and _85618_ (_35753_, _35752_, _35728_);
  not _85619_ (_35754_, _13259_);
  and _85620_ (_35755_, _35754_, _06311_);
  nor _85621_ (_35757_, _35754_, _06311_);
  nor _85622_ (_35758_, _35757_, _35755_);
  not _85623_ (_35759_, _13042_);
  and _85624_ (_35760_, _35759_, _12844_);
  nor _85625_ (_35761_, _35759_, _12844_);
  nor _85626_ (_35762_, _35761_, _35760_);
  nor _85627_ (_35763_, _12197_, _11995_);
  and _85628_ (_35764_, _12197_, _11995_);
  nor _85629_ (_35765_, _35764_, _35763_);
  not _85630_ (_35766_, _12604_);
  and _85631_ (_35768_, _35766_, _12401_);
  nor _85632_ (_35769_, _35766_, _12401_);
  nor _85633_ (_35770_, _35769_, _35768_);
  nor _85634_ (_35771_, _35770_, _35765_);
  and _85635_ (_35772_, _35770_, _35765_);
  nor _85636_ (_35773_, _35772_, _35771_);
  nor _85637_ (_35774_, _35773_, _35762_);
  and _85638_ (_35775_, _35773_, _35762_);
  nor _85639_ (_35776_, _35775_, _35774_);
  and _85640_ (_35777_, _35776_, _35758_);
  nor _85641_ (_35779_, _35776_, _35758_);
  or _85642_ (_35780_, _35779_, _35777_);
  or _85643_ (_35781_, _35780_, _08415_);
  and _85644_ (_35782_, _35781_, _10524_);
  or _85645_ (_35783_, _35782_, _35753_);
  and _85646_ (_35784_, _08652_, _08656_);
  nor _85647_ (_35785_, _35784_, _10389_);
  not _85648_ (_35786_, _35785_);
  and _85649_ (_35787_, _10392_, _08661_);
  nor _85650_ (_35788_, _35787_, _10393_);
  and _85651_ (_35790_, _10395_, _08665_);
  nor _85652_ (_35791_, _35790_, _10396_);
  and _85653_ (_35792_, _35791_, _35788_);
  nor _85654_ (_35793_, _35791_, _35788_);
  nor _85655_ (_35794_, _35793_, _35792_);
  nor _85656_ (_35795_, _35794_, _35786_);
  and _85657_ (_35796_, _35794_, _35786_);
  nor _85658_ (_35797_, _35796_, _35795_);
  and _85659_ (_35798_, _08649_, _08422_);
  nor _85660_ (_35799_, _35798_, _10390_);
  nor _85661_ (_35801_, _35799_, _35797_);
  and _85662_ (_35802_, _35799_, _35797_);
  or _85663_ (_35803_, _35802_, _35801_);
  or _85664_ (_35804_, _35803_, _08416_);
  and _85665_ (_35805_, _35804_, _04499_);
  and _85666_ (_35806_, _35805_, _35783_);
  nor _85667_ (_35807_, _15128_, _14875_);
  and _85668_ (_35808_, _15128_, _14875_);
  nor _85669_ (_35809_, _35808_, _35807_);
  not _85670_ (_35810_, _35809_);
  not _85671_ (_35812_, _15745_);
  and _85672_ (_35813_, _35812_, _15402_);
  nor _85673_ (_35814_, _35812_, _15402_);
  nor _85674_ (_35815_, _35814_, _35813_);
  and _85675_ (_35816_, _35815_, _35810_);
  nor _85676_ (_35817_, _35815_, _35810_);
  or _85677_ (_35818_, _35817_, _35816_);
  nor _85678_ (_35819_, _16750_, _16399_);
  and _85679_ (_35820_, _16750_, _16399_);
  nor _85680_ (_35821_, _35820_, _35819_);
  not _85681_ (_35823_, _16079_);
  and _85682_ (_35824_, _35823_, _08427_);
  nor _85683_ (_35825_, _35823_, _08427_);
  nor _85684_ (_35826_, _35825_, _35824_);
  nor _85685_ (_35827_, _35826_, _35821_);
  and _85686_ (_35828_, _35826_, _35821_);
  nor _85687_ (_35829_, _35828_, _35827_);
  or _85688_ (_35830_, _35829_, _35818_);
  nand _85689_ (_35831_, _35829_, _35818_);
  and _85690_ (_35832_, _35831_, _03636_);
  and _85691_ (_35834_, _35832_, _35830_);
  or _85692_ (_35835_, _35834_, _35806_);
  and _85693_ (_35836_, _35835_, _10531_);
  nor _85694_ (_35837_, _05227_, _04501_);
  or _85695_ (_35838_, _35837_, _03194_);
  and _85696_ (_35839_, _35838_, _34923_);
  or _85697_ (_35840_, _35839_, _35836_);
  and _85698_ (_35841_, _35840_, _10535_);
  nand _85699_ (_35842_, _34923_, _10534_);
  nand _85700_ (_35843_, _35842_, _08435_);
  or _85701_ (_35845_, _35843_, _35841_);
  and _85702_ (_35846_, _35845_, _35028_);
  or _85703_ (_35847_, _35846_, _04135_);
  or _85704_ (_35848_, _35027_, _08440_);
  and _85705_ (_35849_, _35848_, _08446_);
  and _85706_ (_35850_, _35849_, _35847_);
  not _85707_ (_35851_, _07734_);
  or _85708_ (_35852_, _07757_, _07754_);
  nand _85709_ (_35853_, _07757_, _07754_);
  and _85710_ (_35854_, _35853_, _35852_);
  nor _85711_ (_35856_, _07750_, _07749_);
  and _85712_ (_35857_, _07750_, _07749_);
  nor _85713_ (_35858_, _35857_, _35856_);
  not _85714_ (_35859_, _35858_);
  and _85715_ (_35860_, _35859_, _35854_);
  nor _85716_ (_35861_, _35859_, _35854_);
  nor _85717_ (_35862_, _35861_, _35860_);
  not _85718_ (_35863_, _07739_);
  nor _85719_ (_35864_, _07743_, _07736_);
  and _85720_ (_35865_, _07743_, _07736_);
  nor _85721_ (_35867_, _35865_, _35864_);
  nor _85722_ (_35868_, _35867_, _35863_);
  and _85723_ (_35869_, _35867_, _35863_);
  nor _85724_ (_35870_, _35869_, _35868_);
  not _85725_ (_35871_, _35870_);
  nor _85726_ (_35872_, _35871_, _35862_);
  and _85727_ (_35873_, _35871_, _35862_);
  or _85728_ (_35874_, _35873_, _35872_);
  nand _85729_ (_35875_, _35874_, _35851_);
  or _85730_ (_35876_, _35874_, _35851_);
  and _85731_ (_35878_, _35876_, _08445_);
  and _85732_ (_35879_, _35878_, _35875_);
  or _85733_ (_35880_, _35879_, _03755_);
  or _85734_ (_35881_, _35880_, _35850_);
  nor _85735_ (_35882_, _12195_, _11994_);
  and _85736_ (_35883_, _12195_, _11994_);
  nor _85737_ (_35884_, _35883_, _35882_);
  not _85738_ (_35885_, _35884_);
  not _85739_ (_35886_, _12602_);
  and _85740_ (_35887_, _35886_, _12399_);
  nor _85741_ (_35889_, _35886_, _12399_);
  nor _85742_ (_35890_, _35889_, _35887_);
  nor _85743_ (_35891_, _35890_, _35885_);
  and _85744_ (_35892_, _35890_, _35885_);
  nor _85745_ (_35893_, _35892_, _35891_);
  not _85746_ (_35894_, _13257_);
  nor _85747_ (_35895_, _13040_, _12842_);
  and _85748_ (_35896_, _13040_, _12842_);
  nor _85749_ (_35897_, _35896_, _35895_);
  nor _85750_ (_35898_, _35897_, _35894_);
  and _85751_ (_35900_, _35897_, _35894_);
  nor _85752_ (_35901_, _35900_, _35898_);
  not _85753_ (_35902_, _35901_);
  nor _85754_ (_35903_, _35902_, _35893_);
  and _85755_ (_35904_, _35902_, _35893_);
  or _85756_ (_35905_, _35904_, _35903_);
  and _85757_ (_35906_, _35905_, _06309_);
  nor _85758_ (_35907_, _35905_, _06309_);
  or _85759_ (_35908_, _35907_, _35906_);
  or _85760_ (_35909_, _35908_, _07911_);
  and _85761_ (_35911_, _35909_, _07910_);
  and _85762_ (_35912_, _35911_, _35881_);
  not _85763_ (_35913_, _08654_);
  or _85764_ (_35914_, _08666_, _08663_);
  nand _85765_ (_35915_, _08666_, _08663_);
  and _85766_ (_35916_, _35915_, _35914_);
  not _85767_ (_35917_, _08657_);
  and _85768_ (_35918_, _35917_, _08659_);
  nor _85769_ (_35919_, _35917_, _08659_);
  nor _85770_ (_35920_, _35919_, _35918_);
  not _85771_ (_35922_, _35920_);
  and _85772_ (_35923_, _35922_, _35916_);
  nor _85773_ (_35924_, _35922_, _35916_);
  nor _85774_ (_35925_, _35924_, _35923_);
  nand _85775_ (_35926_, _35925_, _35913_);
  or _85776_ (_35927_, _35925_, _35913_);
  and _85777_ (_35928_, _35927_, _35926_);
  or _85778_ (_35929_, _35928_, _08650_);
  nand _85779_ (_35930_, _35928_, _08650_);
  and _85780_ (_35931_, _35930_, _35929_);
  nor _85781_ (_35933_, _35931_, _08646_);
  and _85782_ (_35934_, _35931_, _08646_);
  or _85783_ (_35935_, _35934_, _35933_);
  or _85784_ (_35936_, _35935_, _08421_);
  nand _85785_ (_35937_, _35935_, _08421_);
  and _85786_ (_35938_, _35937_, _07909_);
  and _85787_ (_35939_, _35938_, _35936_);
  or _85788_ (_35940_, _35939_, _35912_);
  and _85789_ (_35941_, _35940_, _05769_);
  and _85790_ (_35942_, _09960_, _09959_);
  nor _85791_ (_35944_, _15623_, _15021_);
  and _85792_ (_35945_, _15623_, _15021_);
  nor _85793_ (_35946_, _35945_, _35944_);
  nor _85794_ (_35947_, _16971_, _16286_);
  and _85795_ (_35948_, _16971_, _16286_);
  nor _85796_ (_35949_, _35948_, _35947_);
  and _85797_ (_35950_, _35949_, _35946_);
  nor _85798_ (_35951_, _35949_, _35946_);
  nor _85799_ (_35952_, _35951_, _35950_);
  not _85800_ (_35953_, _15959_);
  and _85801_ (_35955_, _35953_, _15302_);
  nor _85802_ (_35956_, _35953_, _15302_);
  nor _85803_ (_35957_, _35956_, _35955_);
  nor _85804_ (_35958_, _16630_, _08459_);
  and _85805_ (_35959_, _16630_, _08459_);
  nor _85806_ (_35960_, _35959_, _35958_);
  and _85807_ (_35961_, _35960_, _35957_);
  nor _85808_ (_35962_, _35960_, _35957_);
  nor _85809_ (_35963_, _35962_, _35961_);
  or _85810_ (_35964_, _35963_, _35952_);
  nand _85811_ (_35966_, _35963_, _35952_);
  and _85812_ (_35967_, _35966_, _04504_);
  nand _85813_ (_35968_, _35967_, _35964_);
  nand _85814_ (_35969_, _35968_, _35942_);
  or _85815_ (_35970_, _35969_, _35941_);
  or _85816_ (_35971_, _34923_, _35942_);
  and _85817_ (_35972_, _35971_, _35970_);
  or _85818_ (_35973_, _35972_, _35001_);
  not _85819_ (_35974_, _03487_);
  nor _85820_ (_35975_, _14866_, _07804_);
  and _85821_ (_35977_, _14866_, _07804_);
  nor _85822_ (_35978_, _35977_, _35975_);
  not _85823_ (_35979_, _35978_);
  nor _85824_ (_35980_, _07800_, _07796_);
  and _85825_ (_35981_, _07800_, _07796_);
  nor _85826_ (_35982_, _35981_, _35980_);
  nor _85827_ (_35983_, _35982_, _35979_);
  and _85828_ (_35984_, _35982_, _35979_);
  nor _85829_ (_35985_, _35984_, _35983_);
  nor _85830_ (_35986_, _07793_, _07786_);
  and _85831_ (_35988_, _07793_, _07786_);
  nor _85832_ (_35989_, _35988_, _35986_);
  nor _85833_ (_35990_, _35989_, _07789_);
  and _85834_ (_35991_, _35989_, _07789_);
  nor _85835_ (_35992_, _35991_, _35990_);
  not _85836_ (_35993_, _35992_);
  nor _85837_ (_35994_, _35993_, _35985_);
  and _85838_ (_35995_, _35993_, _35985_);
  nor _85839_ (_35996_, _35995_, _35994_);
  nand _85840_ (_35997_, _35996_, _07783_);
  or _85841_ (_35999_, _35996_, _07783_);
  and _85842_ (_36000_, _35999_, _35997_);
  nand _85843_ (_36001_, _36000_, _35974_);
  nand _85844_ (_36002_, _36001_, _08456_);
  and _85845_ (_36003_, _36002_, _15026_);
  and _85846_ (_36004_, _36003_, _35973_);
  and _85847_ (_36005_, _03487_, _03182_);
  or _85848_ (_36006_, _15027_, _36005_);
  and _85849_ (_36007_, _36006_, _36000_);
  or _85850_ (_36008_, _36007_, _04161_);
  or _85851_ (_36010_, _36008_, _36004_);
  nor _85852_ (_36011_, _36000_, _15029_);
  nor _85853_ (_36012_, _36011_, _26429_);
  and _85854_ (_36013_, _36012_, _36010_);
  nor _85855_ (_36014_, _14877_, _07755_);
  and _85856_ (_36015_, _14877_, _07755_);
  nor _85857_ (_36016_, _36015_, _36014_);
  not _85858_ (_36017_, _36016_);
  nor _85859_ (_36018_, _07751_, _07747_);
  and _85860_ (_36019_, _07751_, _07747_);
  nor _85861_ (_36021_, _36019_, _36018_);
  nor _85862_ (_36022_, _36021_, _36017_);
  and _85863_ (_36023_, _36021_, _36017_);
  nor _85864_ (_36024_, _36023_, _36022_);
  not _85865_ (_36025_, _07740_);
  nor _85866_ (_36026_, _07744_, _07737_);
  and _85867_ (_36027_, _07744_, _07737_);
  nor _85868_ (_36028_, _36027_, _36026_);
  nor _85869_ (_36029_, _36028_, _36025_);
  and _85870_ (_36030_, _36028_, _36025_);
  nor _85871_ (_36032_, _36030_, _36029_);
  nor _85872_ (_36033_, _36032_, _36024_);
  and _85873_ (_36034_, _36032_, _36024_);
  or _85874_ (_36035_, _36034_, _36033_);
  nand _85875_ (_36036_, _36035_, _07733_);
  or _85876_ (_36037_, _36035_, _07733_);
  and _85877_ (_36038_, _36037_, _36036_);
  and _85878_ (_36039_, _36038_, _26429_);
  or _85879_ (_36040_, _36039_, _04165_);
  or _85880_ (_36041_, _36040_, _36013_);
  not _85881_ (_36043_, _04165_);
  or _85882_ (_36044_, _36038_, _36043_);
  and _85883_ (_36045_, _36044_, _08473_);
  and _85884_ (_36046_, _36045_, _36041_);
  nor _85885_ (_36047_, _12196_, _11870_);
  and _85886_ (_36048_, _12196_, _11870_);
  nor _85887_ (_36049_, _36048_, _36047_);
  and _85888_ (_36050_, _36049_, _12400_);
  nor _85889_ (_36051_, _36049_, _12400_);
  or _85890_ (_36052_, _36051_, _36050_);
  nand _85891_ (_36054_, _36052_, _12603_);
  or _85892_ (_36055_, _36052_, _12603_);
  and _85893_ (_36056_, _36055_, _36054_);
  nor _85894_ (_36057_, _13041_, _12843_);
  and _85895_ (_36058_, _13041_, _12843_);
  nor _85896_ (_36059_, _36058_, _36057_);
  nor _85897_ (_36060_, _36059_, _13258_);
  and _85898_ (_36061_, _36059_, _13258_);
  nor _85899_ (_36062_, _36061_, _36060_);
  and _85900_ (_36063_, _36062_, _36056_);
  nor _85901_ (_36065_, _36062_, _36056_);
  nor _85902_ (_36066_, _36065_, _36063_);
  and _85903_ (_36067_, _36066_, _06310_);
  nor _85904_ (_36068_, _36066_, _06310_);
  or _85905_ (_36069_, _36068_, _36067_);
  and _85906_ (_36070_, _36069_, _03761_);
  or _85907_ (_36071_, _36070_, _08477_);
  or _85908_ (_36072_, _36071_, _36046_);
  nor _85909_ (_36073_, _10394_, _08664_);
  and _85910_ (_36074_, _10394_, _08664_);
  nor _85911_ (_36076_, _36074_, _36073_);
  not _85912_ (_36077_, _36076_);
  not _85913_ (_36078_, _08658_);
  and _85914_ (_36079_, _36078_, _08660_);
  nor _85915_ (_36080_, _36078_, _08660_);
  nor _85916_ (_36081_, _36080_, _36079_);
  nor _85917_ (_36082_, _36081_, _36077_);
  and _85918_ (_36083_, _36081_, _36077_);
  nor _85919_ (_36084_, _36083_, _36082_);
  and _85920_ (_36085_, _36084_, _08655_);
  nor _85921_ (_36087_, _36084_, _08655_);
  or _85922_ (_36088_, _36087_, _36085_);
  and _85923_ (_36089_, _36088_, _08651_);
  nor _85924_ (_36090_, _36088_, _08651_);
  or _85925_ (_36091_, _36090_, _36089_);
  and _85926_ (_36092_, _36091_, _08647_);
  nor _85927_ (_36093_, _36091_, _08647_);
  or _85928_ (_36094_, _36093_, _36092_);
  nor _85929_ (_36095_, _36094_, _08420_);
  and _85930_ (_36096_, _36094_, _08420_);
  or _85931_ (_36098_, _36096_, _36095_);
  or _85932_ (_36099_, _36098_, _08480_);
  and _85933_ (_36100_, _36099_, _03759_);
  and _85934_ (_36101_, _36100_, _36072_);
  and _85935_ (_36102_, _10577_, _10573_);
  nor _85936_ (_36103_, _15323_, _15046_);
  and _85937_ (_36104_, _15323_, _15046_);
  or _85938_ (_36105_, _36104_, _36103_);
  nor _85939_ (_36106_, _15732_, _15645_);
  and _85940_ (_36107_, _15732_, _15645_);
  nor _85941_ (_36109_, _36107_, _36106_);
  nor _85942_ (_36110_, _36109_, _36105_);
  and _85943_ (_36111_, _36109_, _36105_);
  nor _85944_ (_36112_, _36111_, _36110_);
  nor _85945_ (_36113_, _16994_, _16653_);
  and _85946_ (_36114_, _16994_, _16653_);
  nor _85947_ (_36115_, _36114_, _36113_);
  not _85948_ (_36116_, _16309_);
  and _85949_ (_36117_, _36116_, _08488_);
  nor _85950_ (_36118_, _36116_, _08488_);
  nor _85951_ (_36120_, _36118_, _36117_);
  nor _85952_ (_36121_, _36120_, _36115_);
  and _85953_ (_36122_, _36120_, _36115_);
  nor _85954_ (_36123_, _36122_, _36121_);
  not _85955_ (_36124_, _36123_);
  nand _85956_ (_36125_, _36124_, _36112_);
  or _85957_ (_36126_, _36124_, _36112_);
  and _85958_ (_36127_, _36126_, _03758_);
  nand _85959_ (_36128_, _36127_, _36125_);
  nand _85960_ (_36129_, _36128_, _36102_);
  or _85961_ (_36131_, _36129_, _36101_);
  or _85962_ (_36132_, _34923_, _36102_);
  and _85963_ (_36133_, _36132_, _07826_);
  and _85964_ (_36134_, _36133_, _36131_);
  or _85965_ (_36135_, _36134_, _35000_);
  or _85966_ (_36136_, _34998_, _07829_);
  and _85967_ (_36137_, _36136_, _08495_);
  and _85968_ (_36138_, _36137_, _36135_);
  not _85969_ (_36139_, _15988_);
  nor _85970_ (_36140_, _15333_, _14943_);
  and _85971_ (_36142_, _15333_, _14943_);
  or _85972_ (_36143_, _36142_, _36140_);
  nor _85973_ (_36144_, _36143_, _15396_);
  and _85974_ (_36145_, _36143_, _15396_);
  nor _85975_ (_36146_, _36145_, _36144_);
  and _85976_ (_36147_, _36146_, _36139_);
  nor _85977_ (_36148_, _36146_, _36139_);
  nor _85978_ (_36149_, _36148_, _36147_);
  and _85979_ (_36150_, _36149_, _16320_);
  nor _85980_ (_36151_, _36149_, _16320_);
  nor _85981_ (_36153_, _36151_, _36150_);
  nor _85982_ (_36154_, _36153_, _16661_);
  and _85983_ (_36155_, _36153_, _16661_);
  or _85984_ (_36156_, _36155_, _36154_);
  nor _85985_ (_36157_, _36156_, _17005_);
  and _85986_ (_36158_, _36156_, _17005_);
  or _85987_ (_36159_, _36158_, _36157_);
  and _85988_ (_36160_, _36159_, _08519_);
  nor _85989_ (_36161_, _36159_, _08519_);
  or _85990_ (_36162_, _36161_, _36160_);
  and _85991_ (_36164_, _36162_, _07825_);
  or _85992_ (_36165_, _36164_, _03765_);
  or _85993_ (_36166_, _36165_, _36138_);
  not _85994_ (_36167_, _15994_);
  nor _85995_ (_36168_, _15119_, _14948_);
  and _85996_ (_36169_, _15119_, _14948_);
  or _85997_ (_36170_, _36169_, _36168_);
  nor _85998_ (_36171_, _36170_, _15658_);
  and _85999_ (_36172_, _36170_, _15658_);
  nor _86000_ (_36173_, _36172_, _36171_);
  and _86001_ (_36175_, _36173_, _36167_);
  nor _86002_ (_36176_, _36173_, _36167_);
  nor _86003_ (_36177_, _36176_, _36175_);
  nor _86004_ (_36178_, _36177_, _16068_);
  and _86005_ (_36179_, _36177_, _16068_);
  or _86006_ (_36180_, _36179_, _36178_);
  and _86007_ (_36181_, _36180_, _16666_);
  nor _86008_ (_36182_, _36180_, _16666_);
  nor _86009_ (_36183_, _36182_, _36181_);
  nor _86010_ (_36184_, _36183_, _17011_);
  and _86011_ (_36186_, _36183_, _17011_);
  or _86012_ (_36187_, _36186_, _36184_);
  nor _86013_ (_36188_, _36187_, _08551_);
  and _86014_ (_36189_, _36187_, _08551_);
  or _86015_ (_36190_, _36189_, _36188_);
  or _86016_ (_36191_, _36190_, _03766_);
  and _86017_ (_36192_, _36191_, _08557_);
  and _86018_ (_36193_, _36192_, _36166_);
  or _86019_ (_36194_, _36193_, _34975_);
  and _86020_ (_36195_, _36194_, _08556_);
  nor _86021_ (_36197_, _15135_, _15134_);
  nor _86022_ (_36198_, _15430_, \oc8051_golden_model_1.ACC [3]);
  and _86023_ (_36199_, _15430_, \oc8051_golden_model_1.ACC [3]);
  nor _86024_ (_36200_, _36199_, _36198_);
  and _86025_ (_36201_, _36200_, _35083_);
  nor _86026_ (_36202_, _36200_, _35083_);
  nor _86027_ (_36203_, _36202_, _36201_);
  not _86028_ (_36204_, _36203_);
  nand _86029_ (_36205_, _36204_, _36197_);
  or _86030_ (_36206_, _36204_, _36197_);
  and _86031_ (_36208_, _36206_, _36205_);
  nand _86032_ (_36209_, _36208_, _08555_);
  and _86033_ (_36210_, _29266_, _11403_);
  nand _86034_ (_36211_, _36210_, _36209_);
  or _86035_ (_36212_, _36211_, _36195_);
  or _86036_ (_36213_, _36210_, _34923_);
  and _86037_ (_36214_, _36213_, _07779_);
  and _86038_ (_36215_, _36214_, _36212_);
  not _86039_ (_36216_, _07779_);
  and _86040_ (_36217_, _14866_, _07805_);
  nor _86041_ (_36219_, _14866_, _07805_);
  or _86042_ (_36220_, _36219_, _36217_);
  and _86043_ (_36221_, _36220_, _15672_);
  nor _86044_ (_36222_, _36220_, _15672_);
  nor _86045_ (_36223_, _36222_, _36221_);
  and _86046_ (_36224_, _36223_, _15728_);
  nor _86047_ (_36225_, _36223_, _15728_);
  nor _86048_ (_36226_, _36225_, _36224_);
  and _86049_ (_36227_, _36226_, _16334_);
  nor _86050_ (_36228_, _36226_, _16334_);
  nor _86051_ (_36230_, _36228_, _36227_);
  nor _86052_ (_36231_, _36230_, _16682_);
  and _86053_ (_36232_, _36230_, _16682_);
  nor _86054_ (_36233_, _36232_, _36231_);
  nor _86055_ (_36234_, _36233_, _17025_);
  and _86056_ (_36235_, _36233_, _17025_);
  or _86057_ (_36236_, _36235_, _36234_);
  nand _86058_ (_36237_, _36236_, _07821_);
  or _86059_ (_36238_, _36236_, _07821_);
  and _86060_ (_36239_, _36238_, _36237_);
  and _86061_ (_36241_, _36239_, _36216_);
  or _86062_ (_36242_, _36241_, _07774_);
  or _86063_ (_36243_, _36242_, _36215_);
  or _86064_ (_36244_, _36239_, _07775_);
  and _86065_ (_36245_, _36244_, _07732_);
  and _86066_ (_36246_, _36245_, _36243_);
  not _86067_ (_36247_, _14877_);
  and _86068_ (_36248_, _36247_, _07756_);
  nor _86069_ (_36249_, _36247_, _07756_);
  nor _86070_ (_36250_, _36249_, _36248_);
  and _86071_ (_36252_, _36250_, _15677_);
  nor _86072_ (_36253_, _36250_, _15677_);
  nor _86073_ (_36254_, _36253_, _36252_);
  and _86074_ (_36255_, _36254_, _16012_);
  nor _86075_ (_36256_, _36254_, _16012_);
  nor _86076_ (_36257_, _36256_, _36255_);
  and _86077_ (_36258_, _36257_, _16339_);
  nor _86078_ (_36259_, _36257_, _16339_);
  nor _86079_ (_36260_, _36259_, _36258_);
  nor _86080_ (_36261_, _36260_, _16690_);
  and _86081_ (_36263_, _36260_, _16690_);
  or _86082_ (_36264_, _36263_, _36261_);
  and _86083_ (_36265_, _36264_, _16743_);
  nor _86084_ (_36266_, _36264_, _16743_);
  or _86085_ (_36267_, _36266_, _36265_);
  nor _86086_ (_36268_, _36267_, _07772_);
  and _86087_ (_36269_, _36267_, _07772_);
  or _86088_ (_36270_, _36269_, _36268_);
  and _86089_ (_36271_, _36270_, _07731_);
  or _86090_ (_36272_, _36271_, _03524_);
  or _86091_ (_36274_, _36272_, _36246_);
  and _86092_ (_36275_, _36274_, _34951_);
  nor _86093_ (_36276_, _15359_, _10395_);
  nor _86094_ (_36277_, _36276_, _35790_);
  nor _86095_ (_36278_, _36277_, _15684_);
  and _86096_ (_36279_, _36277_, _15684_);
  or _86097_ (_36280_, _36279_, _36278_);
  nor _86098_ (_36281_, _36280_, _16025_);
  and _86099_ (_36282_, _36280_, _16025_);
  or _86100_ (_36283_, _36282_, _36281_);
  and _86101_ (_36285_, _36283_, _16350_);
  nor _86102_ (_36286_, _36283_, _16350_);
  nor _86103_ (_36287_, _36286_, _36285_);
  nor _86104_ (_36288_, _36287_, _16701_);
  and _86105_ (_36289_, _36287_, _16701_);
  or _86106_ (_36290_, _36289_, _36288_);
  nor _86107_ (_36291_, _36290_, _17038_);
  and _86108_ (_36292_, _36290_, _17038_);
  or _86109_ (_36293_, _36292_, _36291_);
  not _86110_ (_36294_, _36293_);
  nor _86111_ (_36296_, _36294_, _08681_);
  and _86112_ (_36297_, _36294_, _08681_);
  or _86113_ (_36298_, _36297_, _36296_);
  nand _86114_ (_36299_, _36298_, _08597_);
  and _86115_ (_36300_, _03655_, _03010_);
  nor _86116_ (_36301_, _07729_, _36300_);
  and _86117_ (_36302_, _36301_, _03523_);
  and _86118_ (_36303_, _36302_, _29288_);
  nand _86119_ (_36304_, _36303_, _36299_);
  or _86120_ (_36305_, _36304_, _36275_);
  or _86121_ (_36307_, _36303_, _34923_);
  nor _86122_ (_36308_, _09947_, _12061_);
  not _86123_ (_36309_, _36308_);
  not _86124_ (_36310_, _04193_);
  nor _86125_ (_36311_, _04707_, _03970_);
  and _86126_ (_36312_, _36311_, _36310_);
  and _86127_ (_36313_, _36312_, _36309_);
  and _86128_ (_36314_, _36313_, _36307_);
  and _86129_ (_36315_, _36314_, _36305_);
  not _86130_ (_36316_, _36313_);
  and _86131_ (_36318_, _36316_, _34923_);
  or _86132_ (_36319_, _36318_, _03790_);
  or _86133_ (_36320_, _36319_, _36315_);
  or _86134_ (_36321_, _35118_, _04192_);
  and _86135_ (_36322_, _36321_, _08688_);
  and _86136_ (_36323_, _36322_, _36320_);
  not _86137_ (_36324_, _08693_);
  and _86138_ (_36325_, _15430_, _36324_);
  and _86139_ (_36326_, _36325_, \oc8051_golden_model_1.ACC [3]);
  nor _86140_ (_36327_, _36325_, \oc8051_golden_model_1.ACC [3]);
  nor _86141_ (_36329_, _36327_, _36326_);
  and _86142_ (_36330_, _36329_, _16364_);
  nor _86143_ (_36331_, _36329_, _16364_);
  nor _86144_ (_36332_, _36331_, _36330_);
  and _86145_ (_36333_, _16712_, _07346_);
  nor _86146_ (_36334_, _16712_, _07346_);
  nor _86147_ (_36335_, _36334_, _36333_);
  nor _86148_ (_36336_, _36335_, _36332_);
  and _86149_ (_36337_, _36335_, _36332_);
  or _86150_ (_36338_, _36337_, _36336_);
  nor _86151_ (_36340_, _36338_, _08699_);
  and _86152_ (_36341_, _36338_, _08699_);
  or _86153_ (_36342_, _36341_, _36340_);
  and _86154_ (_36343_, _36342_, _08687_);
  or _86155_ (_36344_, _36343_, _36323_);
  and _86156_ (_36345_, _36344_, _11839_);
  and _86157_ (_36346_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor _86158_ (_36347_, _36346_, _07969_);
  nand _86159_ (_36348_, _36347_, _36203_);
  or _86160_ (_36349_, _36347_, _36203_);
  and _86161_ (_36351_, _36349_, _36348_);
  nand _86162_ (_36352_, _36351_, _08692_);
  nand _86163_ (_36353_, _36352_, _04533_);
  or _86164_ (_36354_, _36353_, _36345_);
  and _86165_ (_36355_, _36354_, _34924_);
  or _86166_ (_36356_, _36355_, _03151_);
  nor _86167_ (_36357_, _35272_, _03152_);
  nor _86168_ (_36358_, _36357_, _03949_);
  and _86169_ (_36359_, _36358_, _36356_);
  nand _86170_ (_36360_, _34923_, _03949_);
  and _86171_ (_36362_, _03483_, _03165_);
  nor _86172_ (_36363_, _26159_, _36362_);
  and _86173_ (_36364_, _36363_, _06712_);
  and _86174_ (_36365_, _06691_, _04208_);
  and _86175_ (_36366_, _36365_, _36364_);
  nand _86176_ (_36367_, _36366_, _36360_);
  or _86177_ (_36368_, _36367_, _36359_);
  or _86178_ (_36369_, _36366_, _34923_);
  and _86179_ (_36370_, _36369_, _03521_);
  and _86180_ (_36371_, _36370_, _36368_);
  not _86181_ (_36373_, _16049_);
  nor _86182_ (_36374_, _15378_, _14903_);
  and _86183_ (_36375_, _15378_, _14903_);
  nor _86184_ (_36376_, _36375_, _36374_);
  and _86185_ (_36377_, _36376_, _15708_);
  nor _86186_ (_36378_, _36376_, _15708_);
  nor _86187_ (_36379_, _36378_, _36377_);
  nor _86188_ (_36380_, _36379_, _36373_);
  and _86189_ (_36381_, _36379_, _36373_);
  or _86190_ (_36382_, _36381_, _36380_);
  and _86191_ (_36384_, _36382_, _16376_);
  nor _86192_ (_36385_, _36382_, _16376_);
  or _86193_ (_36386_, _36385_, _36384_);
  and _86194_ (_36387_, _36386_, _16726_);
  nor _86195_ (_36388_, _36386_, _16726_);
  or _86196_ (_36389_, _36388_, _36387_);
  and _86197_ (_36390_, _36389_, _17061_);
  nor _86198_ (_36391_, _36389_, _17061_);
  or _86199_ (_36392_, _36391_, _36390_);
  and _86200_ (_36393_, _36392_, _08712_);
  nor _86201_ (_36395_, _36392_, _08712_);
  or _86202_ (_36396_, _36395_, _36393_);
  and _86203_ (_36397_, _36396_, _03520_);
  or _86204_ (_36398_, _36397_, _08709_);
  or _86205_ (_36399_, _36398_, _36371_);
  not _86206_ (_36400_, _08717_);
  and _86207_ (_36401_, _15430_, _36400_);
  and _86208_ (_36402_, _36401_, _07500_);
  nor _86209_ (_36403_, _36401_, _07500_);
  nor _86210_ (_36404_, _36403_, _36402_);
  nor _86211_ (_36406_, _36404_, _16381_);
  and _86212_ (_36407_, _36404_, _16381_);
  or _86213_ (_36408_, _36407_, _36406_);
  nor _86214_ (_36409_, _36408_, _17067_);
  and _86215_ (_36410_, _36408_, _17067_);
  or _86216_ (_36411_, _36410_, _36409_);
  not _86217_ (_36412_, _36411_);
  nor _86218_ (_36413_, _16731_, _08724_);
  and _86219_ (_36414_, _16731_, _08724_);
  nor _86220_ (_36415_, _36414_, _36413_);
  nor _86221_ (_36417_, _36415_, _36412_);
  nand _86222_ (_36418_, _36415_, _36412_);
  nand _86223_ (_36419_, _36418_, _08709_);
  nor _86224_ (_36420_, _36419_, _36417_);
  nor _86225_ (_36421_, _03148_, _03079_);
  and _86226_ (_36422_, _36421_, _03165_);
  nor _86227_ (_36423_, _36422_, _36420_);
  and _86228_ (_36424_, _36423_, _36399_);
  and _86229_ (_36425_, _36422_, _34923_);
  or _86230_ (_36426_, _36425_, _10862_);
  or _86231_ (_36428_, _36426_, _36424_);
  or _86232_ (_36429_, _34923_, _10863_);
  and _86233_ (_36430_, _36429_, _42963_);
  and _86234_ (_36431_, _36430_, _36428_);
  or _86235_ (_36432_, _36431_, _34908_);
  and _86236_ (_43388_, _36432_, _41755_);
  and _86237_ (_36433_, _42967_, \oc8051_golden_model_1.PSW [1]);
  or _86238_ (_36434_, _05218_, \oc8051_golden_model_1.PSW [1]);
  and _86239_ (_36435_, _12252_, _05218_);
  not _86240_ (_36436_, _36435_);
  and _86241_ (_36438_, _36436_, _36434_);
  or _86242_ (_36439_, _36438_, _04444_);
  nand _86243_ (_36440_, _05218_, _03233_);
  and _86244_ (_36441_, _36440_, _36434_);
  and _86245_ (_36442_, _36441_, _04426_);
  and _86246_ (_36443_, _04427_, \oc8051_golden_model_1.PSW [1]);
  or _86247_ (_36444_, _36443_, _03570_);
  or _86248_ (_36445_, _36444_, _36442_);
  and _86249_ (_36446_, _36445_, _03517_);
  and _86250_ (_36447_, _36446_, _36439_);
  and _86251_ (_36449_, _12083_, _05783_);
  not _86252_ (_36450_, _05783_);
  and _86253_ (_36451_, _36450_, \oc8051_golden_model_1.PSW [1]);
  or _86254_ (_36452_, _36451_, _03568_);
  or _86255_ (_36453_, _36452_, _36449_);
  and _86256_ (_36454_, _36453_, _14165_);
  or _86257_ (_36455_, _36454_, _36447_);
  nand _86258_ (_36456_, _05218_, _04603_);
  and _86259_ (_36457_, _36456_, _36434_);
  or _86260_ (_36458_, _36457_, _03983_);
  and _86261_ (_36460_, _36458_, _36455_);
  or _86262_ (_36461_, _36460_, _03575_);
  or _86263_ (_36462_, _36441_, _03583_);
  and _86264_ (_36463_, _36462_, _03513_);
  and _86265_ (_36464_, _36463_, _36461_);
  and _86266_ (_36465_, _12069_, _05783_);
  or _86267_ (_36466_, _36465_, _36451_);
  and _86268_ (_36467_, _36466_, _03512_);
  or _86269_ (_36468_, _36467_, _03505_);
  or _86270_ (_36469_, _36468_, _36464_);
  and _86271_ (_36471_, _36449_, _12098_);
  or _86272_ (_36472_, _36451_, _03506_);
  or _86273_ (_36473_, _36472_, _36471_);
  and _86274_ (_36474_, _36473_, _36469_);
  and _86275_ (_36475_, _36474_, _03500_);
  nor _86276_ (_36476_, _12116_, _36450_);
  or _86277_ (_36477_, _36451_, _36476_);
  and _86278_ (_36478_, _36477_, _03499_);
  or _86279_ (_36479_, _36478_, _07314_);
  or _86280_ (_36480_, _36479_, _36475_);
  or _86281_ (_36482_, _36457_, _06039_);
  and _86282_ (_36483_, _36482_, _36480_);
  or _86283_ (_36484_, _36483_, _03479_);
  or _86284_ (_36485_, _06714_, _11451_);
  and _86285_ (_36486_, _36485_, _36434_);
  or _86286_ (_36487_, _36486_, _06044_);
  and _86287_ (_36488_, _36487_, _03474_);
  and _86288_ (_36489_, _36488_, _36484_);
  nand _86289_ (_36490_, _12176_, _05218_);
  and _86290_ (_36491_, _36434_, _03221_);
  and _86291_ (_36493_, _36491_, _36490_);
  or _86292_ (_36494_, _36493_, _36489_);
  and _86293_ (_36495_, _36494_, _03438_);
  nand _86294_ (_36496_, _05218_, _04317_);
  and _86295_ (_36497_, _36434_, _03437_);
  and _86296_ (_36498_, _36497_, _36496_);
  or _86297_ (_36499_, _36498_, _36495_);
  and _86298_ (_36500_, _36499_, _04499_);
  or _86299_ (_36501_, _12191_, _11451_);
  and _86300_ (_36502_, _36434_, _03636_);
  and _86301_ (_36504_, _36502_, _36501_);
  or _86302_ (_36505_, _36504_, _36500_);
  and _86303_ (_36506_, _36505_, _04501_);
  or _86304_ (_36507_, _12197_, _11451_);
  and _86305_ (_36508_, _36434_, _03769_);
  and _86306_ (_36509_, _36508_, _36507_);
  or _86307_ (_36510_, _36509_, _36506_);
  and _86308_ (_36511_, _36510_, _05769_);
  or _86309_ (_36512_, _12190_, _11451_);
  and _86310_ (_36513_, _36512_, _03754_);
  and _86311_ (_36515_, _36513_, _36434_);
  or _86312_ (_36516_, _36515_, _36511_);
  and _86313_ (_36517_, _36516_, _03753_);
  and _86314_ (_36518_, _11451_, \oc8051_golden_model_1.PSW [1]);
  or _86315_ (_36519_, _36518_, _05569_);
  and _86316_ (_36520_, _36441_, _03752_);
  and _86317_ (_36521_, _36520_, _36519_);
  or _86318_ (_36522_, _36521_, _36517_);
  and _86319_ (_36523_, _36522_, _03759_);
  or _86320_ (_36524_, _36496_, _05569_);
  and _86321_ (_36526_, _36434_, _03758_);
  and _86322_ (_36527_, _36526_, _36524_);
  or _86323_ (_36528_, _36527_, _36523_);
  and _86324_ (_36529_, _36528_, _04517_);
  or _86325_ (_36530_, _36440_, _05569_);
  and _86326_ (_36531_, _36434_, _03760_);
  and _86327_ (_36532_, _36531_, _36530_);
  or _86328_ (_36533_, _36532_, _03790_);
  or _86329_ (_36534_, _36533_, _36529_);
  or _86330_ (_36535_, _36438_, _04192_);
  and _86331_ (_36537_, _36535_, _03152_);
  and _86332_ (_36538_, _36537_, _36534_);
  and _86333_ (_36539_, _36466_, _03151_);
  or _86334_ (_36540_, _36539_, _03520_);
  or _86335_ (_36541_, _36540_, _36538_);
  or _86336_ (_36542_, _36518_, _03521_);
  or _86337_ (_36543_, _36542_, _36435_);
  and _86338_ (_36544_, _36543_, _42963_);
  and _86339_ (_36545_, _36544_, _36541_);
  or _86340_ (_36546_, _36545_, _36433_);
  and _86341_ (_43389_, _36546_, _41755_);
  and _86342_ (_36548_, _42967_, \oc8051_golden_model_1.PSW [2]);
  and _86343_ (_36549_, _08292_, \oc8051_golden_model_1.ACC [7]);
  and _86344_ (_36550_, _36549_, _08578_);
  nor _86345_ (_36551_, _08292_, \oc8051_golden_model_1.ACC [7]);
  nor _86346_ (_36552_, _36551_, _36549_);
  not _86347_ (_36553_, _36552_);
  nor _86348_ (_36554_, _36553_, _11808_);
  nor _86349_ (_36555_, _36554_, _36549_);
  and _86350_ (_36556_, _36555_, _08581_);
  or _86351_ (_36558_, _36556_, _36550_);
  and _86352_ (_36559_, _36558_, _08523_);
  and _86353_ (_36560_, _11572_, _03177_);
  and _86354_ (_36561_, _08039_, \oc8051_golden_model_1.ACC [7]);
  and _86355_ (_36562_, _36561_, _08516_);
  nor _86356_ (_36563_, _08039_, \oc8051_golden_model_1.ACC [7]);
  or _86357_ (_36564_, _36563_, _36561_);
  nor _86358_ (_36565_, _36564_, _11797_);
  nor _86359_ (_36566_, _36565_, _36561_);
  and _86360_ (_36567_, _36566_, _08519_);
  or _86361_ (_36569_, _36567_, _36562_);
  and _86362_ (_36570_, _36569_, _36560_);
  and _86363_ (_36571_, _11451_, \oc8051_golden_model_1.PSW [2]);
  nor _86364_ (_36572_, _11451_, _05026_);
  or _86365_ (_36573_, _36572_, _36571_);
  or _86366_ (_36574_, _36573_, _06039_);
  and _86367_ (_36575_, _07834_, \oc8051_golden_model_1.ACC [7]);
  nor _86368_ (_36576_, _07834_, \oc8051_golden_model_1.ACC [7]);
  or _86369_ (_36577_, _36576_, _36575_);
  and _86370_ (_36578_, _36577_, _11711_);
  nor _86371_ (_36580_, _36577_, _11711_);
  nor _86372_ (_36581_, _36580_, _36578_);
  nor _86373_ (_36582_, _36581_, _08032_);
  and _86374_ (_36583_, _36581_, _08032_);
  or _86375_ (_36584_, _36583_, _07922_);
  or _86376_ (_36585_, _36584_, _36582_);
  and _86377_ (_36586_, _36450_, \oc8051_golden_model_1.PSW [2]);
  and _86378_ (_36587_, _12278_, _05783_);
  and _86379_ (_36588_, _36587_, _12309_);
  or _86380_ (_36589_, _36588_, _36586_);
  and _86381_ (_36591_, _36589_, _03505_);
  and _86382_ (_36592_, _12276_, _05783_);
  or _86383_ (_36593_, _36592_, _36586_);
  and _86384_ (_36594_, _36593_, _03512_);
  or _86385_ (_36595_, _36573_, _03983_);
  nor _86386_ (_36596_, _12282_, _11451_);
  or _86387_ (_36597_, _36596_, _36571_);
  or _86388_ (_36598_, _36597_, _04444_);
  and _86389_ (_36599_, _05218_, \oc8051_golden_model_1.ACC [2]);
  or _86390_ (_36600_, _36599_, _36571_);
  and _86391_ (_36602_, _36600_, _04426_);
  and _86392_ (_36603_, _04427_, \oc8051_golden_model_1.PSW [2]);
  or _86393_ (_36604_, _36603_, _03570_);
  or _86394_ (_36605_, _36604_, _36602_);
  and _86395_ (_36606_, _36605_, _03517_);
  and _86396_ (_36607_, _36606_, _36598_);
  or _86397_ (_36608_, _36587_, _36586_);
  and _86398_ (_36609_, _36608_, _03516_);
  or _86399_ (_36610_, _36609_, _03568_);
  or _86400_ (_36611_, _36610_, _36607_);
  and _86401_ (_36613_, _36611_, _36595_);
  or _86402_ (_36614_, _36613_, _03575_);
  or _86403_ (_36615_, _36600_, _03583_);
  and _86404_ (_36616_, _36615_, _03513_);
  and _86405_ (_36617_, _36616_, _36614_);
  or _86406_ (_36618_, _36617_, _36594_);
  and _86407_ (_36619_, _36618_, _03506_);
  or _86408_ (_36620_, _36619_, _36591_);
  and _86409_ (_36621_, _36620_, _06800_);
  or _86410_ (_36622_, _14192_, _14084_);
  or _86411_ (_36624_, _36622_, _14313_);
  or _86412_ (_36625_, _36624_, _14431_);
  or _86413_ (_36626_, _36625_, _14549_);
  or _86414_ (_36627_, _36626_, _14667_);
  or _86415_ (_36628_, _36627_, _14788_);
  or _86416_ (_36629_, _36628_, _07310_);
  and _86417_ (_36630_, _36629_, _06794_);
  or _86418_ (_36631_, _36630_, _07923_);
  or _86419_ (_36632_, _36631_, _36621_);
  and _86420_ (_36633_, _36632_, _08037_);
  and _86421_ (_36635_, _36633_, _36585_);
  or _86422_ (_36636_, _36564_, _11464_);
  nand _86423_ (_36637_, _36564_, _11464_);
  and _86424_ (_36638_, _36637_, _36636_);
  and _86425_ (_36639_, _36638_, _08104_);
  nor _86426_ (_36640_, _36638_, _08104_);
  or _86427_ (_36641_, _36640_, _36639_);
  and _86428_ (_36642_, _36641_, _08035_);
  or _86429_ (_36643_, _36642_, _36635_);
  and _86430_ (_36644_, _36643_, _03619_);
  not _86431_ (_36646_, _08227_);
  and _86432_ (_36647_, _11729_, _36646_);
  nor _86433_ (_36648_, _11729_, _36646_);
  or _86434_ (_36649_, _36648_, _36647_);
  nand _86435_ (_36650_, _36649_, _08281_);
  or _86436_ (_36651_, _36649_, _08281_);
  and _86437_ (_36652_, _36651_, _36650_);
  or _86438_ (_36653_, _36652_, _08108_);
  and _86439_ (_36654_, _36653_, _10431_);
  or _86440_ (_36655_, _36654_, _36644_);
  or _86441_ (_36657_, _36553_, _11739_);
  nand _86442_ (_36658_, _36553_, _11739_);
  and _86443_ (_36659_, _36658_, _36657_);
  and _86444_ (_36660_, _36659_, _08351_);
  nor _86445_ (_36661_, _36659_, _08351_);
  or _86446_ (_36662_, _36661_, _36660_);
  or _86447_ (_36663_, _36662_, _08109_);
  and _86448_ (_36664_, _36663_, _03500_);
  and _86449_ (_36665_, _36664_, _36655_);
  nor _86450_ (_36666_, _12326_, _36450_);
  or _86451_ (_36668_, _36666_, _36586_);
  and _86452_ (_36669_, _36668_, _03499_);
  or _86453_ (_36670_, _36669_, _07314_);
  or _86454_ (_36671_, _36670_, _36665_);
  and _86455_ (_36672_, _36671_, _36574_);
  or _86456_ (_36673_, _36672_, _03479_);
  and _86457_ (_36674_, _06718_, _05218_);
  or _86458_ (_36675_, _36571_, _06044_);
  or _86459_ (_36676_, _36675_, _36674_);
  and _86460_ (_36677_, _36676_, _03474_);
  and _86461_ (_36679_, _36677_, _36673_);
  nor _86462_ (_36680_, _12384_, _11451_);
  or _86463_ (_36681_, _36680_, _36571_);
  and _86464_ (_36682_, _36681_, _03221_);
  or _86465_ (_36683_, _36682_, _07328_);
  or _86466_ (_36684_, _36683_, _36679_);
  nand _86467_ (_36685_, _07344_, _07340_);
  nand _86468_ (_36686_, _36685_, _07328_);
  and _86469_ (_36687_, _36686_, _36684_);
  or _86470_ (_36688_, _36687_, _03437_);
  and _86471_ (_36690_, _05218_, _06261_);
  or _86472_ (_36691_, _36690_, _36571_);
  or _86473_ (_36692_, _36691_, _03438_);
  and _86474_ (_36693_, _36692_, _04499_);
  and _86475_ (_36694_, _36693_, _36688_);
  and _86476_ (_36695_, _12273_, _05218_);
  or _86477_ (_36696_, _36695_, _36571_);
  and _86478_ (_36697_, _36696_, _03636_);
  or _86479_ (_36698_, _36697_, _03769_);
  or _86480_ (_36699_, _36698_, _36694_);
  and _86481_ (_36701_, _12401_, _05218_);
  or _86482_ (_36702_, _36701_, _36571_);
  or _86483_ (_36703_, _36702_, _04501_);
  and _86484_ (_36704_, _36703_, _05769_);
  and _86485_ (_36705_, _36704_, _36699_);
  or _86486_ (_36706_, _36571_, _05665_);
  and _86487_ (_36707_, _36706_, _03754_);
  and _86488_ (_36708_, _36707_, _36691_);
  or _86489_ (_36709_, _36708_, _36705_);
  and _86490_ (_36710_, _36709_, _03753_);
  and _86491_ (_36712_, _36600_, _03752_);
  and _86492_ (_36713_, _36712_, _36706_);
  or _86493_ (_36714_, _36713_, _03758_);
  or _86494_ (_36715_, _36714_, _36710_);
  nor _86495_ (_36716_, _12272_, _11451_);
  or _86496_ (_36717_, _36571_, _03759_);
  or _86497_ (_36718_, _36717_, _36716_);
  and _86498_ (_36719_, _36718_, _04517_);
  and _86499_ (_36720_, _36719_, _36715_);
  nor _86500_ (_36721_, _12400_, _11451_);
  or _86501_ (_36723_, _36721_, _36571_);
  and _86502_ (_36724_, _36723_, _03760_);
  or _86503_ (_36725_, _36724_, _08490_);
  or _86504_ (_36726_, _36725_, _36720_);
  not _86505_ (_36727_, _36560_);
  nor _86506_ (_36728_, _36577_, _11444_);
  nor _86507_ (_36729_, _36728_, _36575_);
  and _86508_ (_36730_, _36729_, _07907_);
  and _86509_ (_36731_, _36575_, _07904_);
  or _86510_ (_36732_, _36731_, _07830_);
  or _86511_ (_36734_, _36732_, _36730_);
  and _86512_ (_36735_, _36734_, _36727_);
  and _86513_ (_36736_, _36735_, _36726_);
  or _86514_ (_36737_, _36736_, _36570_);
  and _86515_ (_36738_, _36737_, _04154_);
  and _86516_ (_36739_, _36569_, _04153_);
  or _86517_ (_36740_, _36739_, _03765_);
  or _86518_ (_36741_, _36740_, _36738_);
  and _86519_ (_36742_, _08226_, \oc8051_golden_model_1.ACC [7]);
  and _86520_ (_36743_, _36742_, _08548_);
  nor _86521_ (_36745_, _08226_, \oc8051_golden_model_1.ACC [7]);
  nor _86522_ (_36746_, _36745_, _11802_);
  nor _86523_ (_36747_, _36746_, _36742_);
  and _86524_ (_36748_, _36747_, _08551_);
  or _86525_ (_36749_, _36748_, _36743_);
  or _86526_ (_36750_, _36749_, _03766_);
  and _86527_ (_36751_, _36750_, _08557_);
  and _86528_ (_36752_, _36751_, _36741_);
  or _86529_ (_36753_, _36752_, _36559_);
  and _86530_ (_36754_, _36753_, _07780_);
  nand _86531_ (_36756_, _07818_, _11437_);
  and _86532_ (_36757_, _36756_, _11439_);
  or _86533_ (_36758_, _36757_, _15068_);
  or _86534_ (_36759_, _36758_, _36754_);
  nand _86535_ (_36760_, _07769_, _35851_);
  or _86536_ (_36761_, _07769_, _07733_);
  and _86537_ (_36762_, _36761_, _36760_);
  or _86538_ (_36763_, _36762_, _15075_);
  and _86539_ (_36764_, _36763_, _36759_);
  or _86540_ (_36765_, _36764_, _15073_);
  or _86541_ (_36767_, _36762_, _15074_);
  and _86542_ (_36768_, _36767_, _09936_);
  and _86543_ (_36769_, _36768_, _36765_);
  or _86544_ (_36770_, _08639_, _08599_);
  and _86545_ (_36771_, _36770_, _11829_);
  nand _86546_ (_36772_, _08678_, _11833_);
  and _86547_ (_36773_, _36772_, _11835_);
  or _86548_ (_36774_, _36773_, _03790_);
  or _86549_ (_36775_, _36774_, _36771_);
  or _86550_ (_36776_, _36775_, _36769_);
  or _86551_ (_36778_, _36597_, _04192_);
  and _86552_ (_36779_, _36778_, _03152_);
  and _86553_ (_36780_, _36779_, _36776_);
  and _86554_ (_36781_, _36593_, _03151_);
  or _86555_ (_36782_, _36781_, _03520_);
  or _86556_ (_36783_, _36782_, _36780_);
  and _86557_ (_36784_, _12456_, _05218_);
  or _86558_ (_36785_, _36571_, _03521_);
  or _86559_ (_36786_, _36785_, _36784_);
  and _86560_ (_36787_, _36786_, _42963_);
  and _86561_ (_36789_, _36787_, _36783_);
  or _86562_ (_36790_, _36789_, _36548_);
  and _86563_ (_43390_, _36790_, _41755_);
  nor _86564_ (_36791_, _42963_, _04856_);
  nor _86565_ (_36792_, _05218_, _04856_);
  nor _86566_ (_36793_, _12486_, _11451_);
  or _86567_ (_36794_, _36793_, _36792_);
  or _86568_ (_36795_, _36794_, _04444_);
  and _86569_ (_36796_, _05218_, \oc8051_golden_model_1.ACC [3]);
  or _86570_ (_36797_, _36796_, _36792_);
  and _86571_ (_36799_, _36797_, _04426_);
  nor _86572_ (_36800_, _04426_, _04856_);
  or _86573_ (_36801_, _36800_, _03570_);
  or _86574_ (_36802_, _36801_, _36799_);
  and _86575_ (_36803_, _36802_, _03517_);
  and _86576_ (_36804_, _36803_, _36795_);
  nor _86577_ (_36805_, _05783_, _04856_);
  and _86578_ (_36806_, _12490_, _05783_);
  or _86579_ (_36807_, _36806_, _36805_);
  and _86580_ (_36808_, _36807_, _03516_);
  or _86581_ (_36810_, _36808_, _03568_);
  or _86582_ (_36811_, _36810_, _36804_);
  nor _86583_ (_36812_, _11451_, _04843_);
  or _86584_ (_36813_, _36812_, _36792_);
  or _86585_ (_36814_, _36813_, _03983_);
  and _86586_ (_36815_, _36814_, _36811_);
  or _86587_ (_36816_, _36815_, _03575_);
  or _86588_ (_36817_, _36797_, _03583_);
  and _86589_ (_36818_, _36817_, _03513_);
  and _86590_ (_36819_, _36818_, _36816_);
  and _86591_ (_36821_, _12500_, _05783_);
  or _86592_ (_36822_, _36821_, _36805_);
  and _86593_ (_36823_, _36822_, _03512_);
  or _86594_ (_36824_, _36823_, _03505_);
  or _86595_ (_36825_, _36824_, _36819_);
  or _86596_ (_36826_, _36805_, _12507_);
  and _86597_ (_36827_, _36826_, _36807_);
  or _86598_ (_36828_, _36827_, _03506_);
  and _86599_ (_36829_, _36828_, _03500_);
  and _86600_ (_36830_, _36829_, _36825_);
  nor _86601_ (_36832_, _12525_, _36450_);
  or _86602_ (_36833_, _36832_, _36805_);
  and _86603_ (_36834_, _36833_, _03499_);
  or _86604_ (_36835_, _36834_, _07314_);
  or _86605_ (_36836_, _36835_, _36830_);
  or _86606_ (_36837_, _36813_, _06039_);
  and _86607_ (_36838_, _36837_, _06044_);
  and _86608_ (_36839_, _36838_, _36836_);
  and _86609_ (_36840_, _06717_, _05218_);
  or _86610_ (_36841_, _36840_, _36792_);
  and _86611_ (_36843_, _36841_, _03479_);
  or _86612_ (_36844_, _36843_, _03221_);
  or _86613_ (_36845_, _36844_, _36839_);
  nor _86614_ (_36846_, _12583_, _11451_);
  or _86615_ (_36847_, _36846_, _36792_);
  or _86616_ (_36848_, _36847_, _03474_);
  and _86617_ (_36849_, _36848_, _03438_);
  and _86618_ (_36850_, _36849_, _36845_);
  and _86619_ (_36851_, _05218_, _06217_);
  or _86620_ (_36852_, _36851_, _36792_);
  and _86621_ (_36854_, _36852_, _03437_);
  or _86622_ (_36855_, _36854_, _03636_);
  or _86623_ (_36856_, _36855_, _36850_);
  and _86624_ (_36857_, _12598_, _05218_);
  or _86625_ (_36858_, _36857_, _36792_);
  or _86626_ (_36859_, _36858_, _04499_);
  and _86627_ (_36860_, _36859_, _36856_);
  or _86628_ (_36861_, _36860_, _03769_);
  and _86629_ (_36862_, _12604_, _05218_);
  or _86630_ (_36863_, _36862_, _36792_);
  or _86631_ (_36865_, _36863_, _04501_);
  and _86632_ (_36866_, _36865_, _05769_);
  and _86633_ (_36867_, _36866_, _36861_);
  or _86634_ (_36868_, _36792_, _05521_);
  and _86635_ (_36869_, _36852_, _04504_);
  and _86636_ (_36870_, _36869_, _36868_);
  or _86637_ (_36871_, _36870_, _36867_);
  and _86638_ (_36872_, _36871_, _03753_);
  and _86639_ (_36873_, _36797_, _03752_);
  and _86640_ (_36874_, _36873_, _36868_);
  or _86641_ (_36876_, _36874_, _03758_);
  or _86642_ (_36877_, _36876_, _36872_);
  nor _86643_ (_36878_, _12597_, _11451_);
  or _86644_ (_36879_, _36792_, _03759_);
  or _86645_ (_36880_, _36879_, _36878_);
  and _86646_ (_36881_, _36880_, _04517_);
  and _86647_ (_36882_, _36881_, _36877_);
  nor _86648_ (_36883_, _12603_, _11451_);
  or _86649_ (_36884_, _36883_, _36792_);
  and _86650_ (_36885_, _36884_, _03760_);
  or _86651_ (_36887_, _36885_, _03790_);
  or _86652_ (_36888_, _36887_, _36882_);
  or _86653_ (_36889_, _36794_, _04192_);
  and _86654_ (_36890_, _36889_, _03152_);
  and _86655_ (_36891_, _36890_, _36888_);
  and _86656_ (_36892_, _36822_, _03151_);
  or _86657_ (_36893_, _36892_, _03520_);
  or _86658_ (_36894_, _36893_, _36891_);
  and _86659_ (_36895_, _12658_, _05218_);
  or _86660_ (_36896_, _36792_, _03521_);
  or _86661_ (_36898_, _36896_, _36895_);
  and _86662_ (_36899_, _36898_, _42963_);
  and _86663_ (_36900_, _36899_, _36894_);
  or _86664_ (_36901_, _36900_, _36791_);
  and _86665_ (_43393_, _36901_, _41755_);
  and _86666_ (_36902_, _42967_, \oc8051_golden_model_1.PSW [4]);
  and _86667_ (_36903_, _11451_, \oc8051_golden_model_1.PSW [4]);
  and _86668_ (_36904_, _06722_, _05218_);
  or _86669_ (_36905_, _36904_, _36903_);
  or _86670_ (_36906_, _36905_, _06044_);
  nor _86671_ (_36908_, _05712_, _11451_);
  or _86672_ (_36909_, _36908_, _36903_);
  or _86673_ (_36910_, _36909_, _06039_);
  nor _86674_ (_36911_, _12733_, _11451_);
  or _86675_ (_36912_, _36911_, _36903_);
  or _86676_ (_36913_, _36912_, _04444_);
  and _86677_ (_36914_, _05218_, \oc8051_golden_model_1.ACC [4]);
  or _86678_ (_36915_, _36914_, _36903_);
  and _86679_ (_36916_, _36915_, _04426_);
  and _86680_ (_36917_, _04427_, \oc8051_golden_model_1.PSW [4]);
  or _86681_ (_36919_, _36917_, _03570_);
  or _86682_ (_36920_, _36919_, _36916_);
  and _86683_ (_36921_, _36920_, _03517_);
  and _86684_ (_36922_, _36921_, _36913_);
  and _86685_ (_36923_, _36450_, \oc8051_golden_model_1.PSW [4]);
  and _86686_ (_36924_, _12737_, _05783_);
  or _86687_ (_36925_, _36924_, _36923_);
  and _86688_ (_36926_, _36925_, _03516_);
  or _86689_ (_36927_, _36926_, _03568_);
  or _86690_ (_36928_, _36927_, _36922_);
  or _86691_ (_36930_, _36909_, _03983_);
  and _86692_ (_36931_, _36930_, _36928_);
  or _86693_ (_36932_, _36931_, _03575_);
  or _86694_ (_36933_, _36915_, _03583_);
  and _86695_ (_36934_, _36933_, _03513_);
  and _86696_ (_36935_, _36934_, _36932_);
  and _86697_ (_36936_, _12718_, _05783_);
  or _86698_ (_36937_, _36936_, _36923_);
  and _86699_ (_36938_, _36937_, _03512_);
  or _86700_ (_36939_, _36938_, _03505_);
  or _86701_ (_36941_, _36939_, _36935_);
  or _86702_ (_36942_, _36923_, _12752_);
  and _86703_ (_36943_, _36942_, _36925_);
  or _86704_ (_36944_, _36943_, _03506_);
  and _86705_ (_36945_, _36944_, _03500_);
  and _86706_ (_36946_, _36945_, _36941_);
  nor _86707_ (_36947_, _12716_, _36450_);
  or _86708_ (_36948_, _36947_, _36923_);
  and _86709_ (_36949_, _36948_, _03499_);
  or _86710_ (_36950_, _36949_, _07314_);
  or _86711_ (_36952_, _36950_, _36946_);
  and _86712_ (_36953_, _36952_, _36910_);
  and _86713_ (_36954_, _11572_, _03186_);
  and _86714_ (_36955_, _36905_, _04069_);
  or _86715_ (_36956_, _36955_, _36954_);
  or _86716_ (_36957_, _36956_, _36953_);
  and _86717_ (_36958_, _36957_, _36906_);
  or _86718_ (_36959_, _36958_, _03221_);
  nor _86719_ (_36960_, _12827_, _11451_);
  or _86720_ (_36961_, _36960_, _36903_);
  or _86721_ (_36963_, _36961_, _03474_);
  and _86722_ (_36964_, _36963_, _36959_);
  or _86723_ (_36965_, _36964_, _03437_);
  and _86724_ (_36966_, _06233_, _05218_);
  or _86725_ (_36967_, _36966_, _36903_);
  or _86726_ (_36968_, _36967_, _03438_);
  and _86727_ (_36969_, _36968_, _04499_);
  and _86728_ (_36970_, _36969_, _36965_);
  and _86729_ (_36971_, _12711_, _05218_);
  or _86730_ (_36972_, _36971_, _36903_);
  and _86731_ (_36974_, _36972_, _03636_);
  or _86732_ (_36975_, _36974_, _03769_);
  or _86733_ (_36976_, _36975_, _36970_);
  and _86734_ (_36977_, _12844_, _05218_);
  or _86735_ (_36978_, _36977_, _36903_);
  or _86736_ (_36979_, _36978_, _04501_);
  and _86737_ (_36980_, _36979_, _05769_);
  and _86738_ (_36981_, _36980_, _36976_);
  or _86739_ (_36982_, _36903_, _05761_);
  and _86740_ (_36983_, _36982_, _03754_);
  and _86741_ (_36985_, _36983_, _36967_);
  or _86742_ (_36986_, _36985_, _36981_);
  and _86743_ (_36987_, _36986_, _03753_);
  and _86744_ (_36988_, _36915_, _03752_);
  and _86745_ (_36989_, _36988_, _36982_);
  or _86746_ (_36990_, _36989_, _03758_);
  or _86747_ (_36991_, _36990_, _36987_);
  nor _86748_ (_36992_, _12710_, _11451_);
  or _86749_ (_36993_, _36903_, _03759_);
  or _86750_ (_36994_, _36993_, _36992_);
  and _86751_ (_36996_, _36994_, _04517_);
  and _86752_ (_36997_, _36996_, _36991_);
  nor _86753_ (_36998_, _12843_, _11451_);
  or _86754_ (_36999_, _36998_, _36903_);
  and _86755_ (_37000_, _36999_, _03760_);
  or _86756_ (_37001_, _37000_, _03790_);
  or _86757_ (_37002_, _37001_, _36997_);
  or _86758_ (_37003_, _36912_, _04192_);
  and _86759_ (_37004_, _37003_, _03152_);
  and _86760_ (_37005_, _37004_, _37002_);
  and _86761_ (_37007_, _36937_, _03151_);
  or _86762_ (_37008_, _37007_, _03520_);
  or _86763_ (_37009_, _37008_, _37005_);
  and _86764_ (_37010_, _12893_, _05218_);
  or _86765_ (_37011_, _36903_, _03521_);
  or _86766_ (_37012_, _37011_, _37010_);
  and _86767_ (_37013_, _37012_, _42963_);
  and _86768_ (_37014_, _37013_, _37009_);
  or _86769_ (_37015_, _37014_, _36902_);
  and _86770_ (_43394_, _37015_, _41755_);
  and _86771_ (_37017_, _42967_, \oc8051_golden_model_1.PSW [5]);
  and _86772_ (_37018_, _11451_, \oc8051_golden_model_1.PSW [5]);
  nor _86773_ (_37019_, _12930_, _11451_);
  or _86774_ (_37020_, _37019_, _37018_);
  or _86775_ (_37021_, _37020_, _04444_);
  and _86776_ (_37022_, _05218_, \oc8051_golden_model_1.ACC [5]);
  or _86777_ (_37023_, _37022_, _37018_);
  and _86778_ (_37024_, _37023_, _04426_);
  and _86779_ (_37025_, _04427_, \oc8051_golden_model_1.PSW [5]);
  or _86780_ (_37026_, _37025_, _03570_);
  or _86781_ (_37028_, _37026_, _37024_);
  and _86782_ (_37029_, _37028_, _03517_);
  and _86783_ (_37030_, _37029_, _37021_);
  and _86784_ (_37031_, _36450_, \oc8051_golden_model_1.PSW [5]);
  and _86785_ (_37032_, _12934_, _05783_);
  or _86786_ (_37033_, _37032_, _37031_);
  and _86787_ (_37034_, _37033_, _03516_);
  or _86788_ (_37035_, _37034_, _03568_);
  or _86789_ (_37036_, _37035_, _37030_);
  nor _86790_ (_37037_, _05422_, _11451_);
  or _86791_ (_37039_, _37037_, _37018_);
  or _86792_ (_37040_, _37039_, _03983_);
  and _86793_ (_37041_, _37040_, _37036_);
  or _86794_ (_37042_, _37041_, _03575_);
  or _86795_ (_37043_, _37023_, _03583_);
  and _86796_ (_37044_, _37043_, _03513_);
  and _86797_ (_37045_, _37044_, _37042_);
  and _86798_ (_37046_, _12914_, _05783_);
  or _86799_ (_37047_, _37046_, _37031_);
  and _86800_ (_37048_, _37047_, _03512_);
  or _86801_ (_37050_, _37048_, _03505_);
  or _86802_ (_37051_, _37050_, _37045_);
  or _86803_ (_37052_, _37031_, _12949_);
  and _86804_ (_37053_, _37052_, _37033_);
  or _86805_ (_37054_, _37053_, _03506_);
  and _86806_ (_37055_, _37054_, _03500_);
  and _86807_ (_37056_, _37055_, _37051_);
  nor _86808_ (_37057_, _12912_, _36450_);
  or _86809_ (_37058_, _37057_, _37031_);
  and _86810_ (_37059_, _37058_, _03499_);
  or _86811_ (_37061_, _37059_, _07314_);
  or _86812_ (_37062_, _37061_, _37056_);
  or _86813_ (_37063_, _37039_, _06039_);
  and _86814_ (_37064_, _37063_, _06044_);
  and _86815_ (_37065_, _37064_, _37062_);
  and _86816_ (_37066_, _06721_, _05218_);
  or _86817_ (_37067_, _37066_, _37018_);
  and _86818_ (_37068_, _37067_, _03479_);
  or _86819_ (_37069_, _37068_, _03221_);
  or _86820_ (_37070_, _37069_, _37065_);
  nor _86821_ (_37072_, _13021_, _11451_);
  or _86822_ (_37073_, _37072_, _37018_);
  or _86823_ (_37074_, _37073_, _03474_);
  and _86824_ (_37075_, _37074_, _03438_);
  and _86825_ (_37076_, _37075_, _37070_);
  and _86826_ (_37077_, _06211_, _05218_);
  or _86827_ (_37078_, _37077_, _37018_);
  and _86828_ (_37079_, _37078_, _03437_);
  or _86829_ (_37080_, _37079_, _03636_);
  or _86830_ (_37081_, _37080_, _37076_);
  and _86831_ (_37083_, _13036_, _05218_);
  or _86832_ (_37084_, _37083_, _37018_);
  or _86833_ (_37085_, _37084_, _04499_);
  and _86834_ (_37086_, _37085_, _37081_);
  or _86835_ (_37087_, _37086_, _03769_);
  and _86836_ (_37088_, _13042_, _05218_);
  or _86837_ (_37089_, _37088_, _37018_);
  or _86838_ (_37090_, _37089_, _04501_);
  and _86839_ (_37091_, _37090_, _05769_);
  and _86840_ (_37092_, _37091_, _37087_);
  or _86841_ (_37094_, _37018_, _05472_);
  and _86842_ (_37095_, _37078_, _04504_);
  and _86843_ (_37096_, _37095_, _37094_);
  or _86844_ (_37097_, _37096_, _37092_);
  and _86845_ (_37098_, _37097_, _03753_);
  and _86846_ (_37099_, _37023_, _03752_);
  and _86847_ (_37100_, _37099_, _37094_);
  or _86848_ (_37101_, _37100_, _03758_);
  or _86849_ (_37102_, _37101_, _37098_);
  nor _86850_ (_37103_, _13035_, _11451_);
  or _86851_ (_37105_, _37018_, _03759_);
  or _86852_ (_37106_, _37105_, _37103_);
  and _86853_ (_37107_, _37106_, _04517_);
  and _86854_ (_37108_, _37107_, _37102_);
  nor _86855_ (_37109_, _13041_, _11451_);
  or _86856_ (_37110_, _37109_, _37018_);
  and _86857_ (_37111_, _37110_, _03760_);
  or _86858_ (_37112_, _37111_, _03790_);
  or _86859_ (_37113_, _37112_, _37108_);
  or _86860_ (_37114_, _37020_, _04192_);
  and _86861_ (_37116_, _37114_, _03152_);
  and _86862_ (_37117_, _37116_, _37113_);
  and _86863_ (_37118_, _37047_, _03151_);
  or _86864_ (_37119_, _37118_, _03520_);
  or _86865_ (_37120_, _37119_, _37117_);
  and _86866_ (_37121_, _13097_, _05218_);
  or _86867_ (_37122_, _37018_, _03521_);
  or _86868_ (_37123_, _37122_, _37121_);
  and _86869_ (_37124_, _37123_, _42963_);
  and _86870_ (_37125_, _37124_, _37120_);
  or _86871_ (_37127_, _37125_, _37017_);
  and _86872_ (_43395_, _37127_, _41755_);
  nor _86873_ (_37128_, _42963_, _15797_);
  or _86874_ (_37129_, _07898_, _07850_);
  and _86875_ (_37130_, _03489_, _03177_);
  and _86876_ (_37131_, _03664_, _03177_);
  nor _86877_ (_37132_, _37131_, _37130_);
  not _86878_ (_37133_, _37132_);
  and _86879_ (_37134_, _37133_, _37129_);
  and _86880_ (_37135_, _37129_, _03953_);
  nor _86881_ (_37137_, _13251_, _11451_);
  nor _86882_ (_37138_, _05218_, _15797_);
  or _86883_ (_37139_, _37138_, _03759_);
  or _86884_ (_37140_, _37139_, _37137_);
  nor _86885_ (_37141_, _05783_, _15797_);
  and _86886_ (_37142_, _13145_, _05783_);
  or _86887_ (_37143_, _37142_, _37141_);
  or _86888_ (_37144_, _37141_, _13160_);
  and _86889_ (_37145_, _37144_, _37143_);
  or _86890_ (_37146_, _37145_, _03506_);
  nor _86891_ (_37148_, _13122_, _11451_);
  or _86892_ (_37149_, _37148_, _37138_);
  or _86893_ (_37150_, _37149_, _04444_);
  and _86894_ (_37151_, _05218_, \oc8051_golden_model_1.ACC [6]);
  or _86895_ (_37152_, _37151_, _37138_);
  and _86896_ (_37153_, _37152_, _04426_);
  nor _86897_ (_37154_, _04426_, _15797_);
  or _86898_ (_37155_, _37154_, _03570_);
  or _86899_ (_37156_, _37155_, _37153_);
  and _86900_ (_37157_, _37156_, _03517_);
  and _86901_ (_37159_, _37157_, _37150_);
  and _86902_ (_37160_, _37143_, _03516_);
  or _86903_ (_37161_, _37160_, _03568_);
  or _86904_ (_37162_, _37161_, _37159_);
  nor _86905_ (_37163_, _05327_, _11451_);
  or _86906_ (_37164_, _37163_, _37138_);
  or _86907_ (_37165_, _37164_, _03983_);
  and _86908_ (_37166_, _37165_, _37162_);
  or _86909_ (_37167_, _37166_, _03575_);
  or _86910_ (_37168_, _37152_, _03583_);
  and _86911_ (_37170_, _37168_, _03513_);
  and _86912_ (_37171_, _37170_, _37167_);
  and _86913_ (_37172_, _13130_, _05783_);
  or _86914_ (_37173_, _37172_, _37141_);
  and _86915_ (_37174_, _37173_, _03512_);
  or _86916_ (_37175_, _37174_, _03505_);
  or _86917_ (_37176_, _37175_, _37171_);
  and _86918_ (_37177_, _37176_, _37146_);
  and _86919_ (_37178_, _37177_, _07922_);
  or _86920_ (_37179_, _08022_, _07850_);
  and _86921_ (_37181_, _37179_, _07923_);
  or _86922_ (_37182_, _37181_, _08035_);
  or _86923_ (_37183_, _37182_, _37178_);
  or _86924_ (_37184_, _08057_, _08037_);
  or _86925_ (_37185_, _37184_, _08094_);
  and _86926_ (_37186_, _37185_, _37183_);
  or _86927_ (_37187_, _37186_, _10431_);
  or _86928_ (_37188_, _08195_, _03619_);
  or _86929_ (_37189_, _37188_, _08275_);
  or _86930_ (_37190_, _08289_, _08109_);
  or _86931_ (_37192_, _37190_, _08341_);
  and _86932_ (_37193_, _37192_, _03500_);
  and _86933_ (_37194_, _37193_, _37189_);
  and _86934_ (_37195_, _37194_, _37187_);
  nor _86935_ (_37196_, _13178_, _36450_);
  or _86936_ (_37197_, _37196_, _37141_);
  and _86937_ (_37198_, _37197_, _03499_);
  or _86938_ (_37199_, _37198_, _07314_);
  or _86939_ (_37200_, _37199_, _37195_);
  or _86940_ (_37201_, _37164_, _06039_);
  and _86941_ (_37203_, _37201_, _06044_);
  and _86942_ (_37204_, _37203_, _37200_);
  and _86943_ (_37205_, _06713_, _05218_);
  or _86944_ (_37206_, _37205_, _37138_);
  and _86945_ (_37207_, _37206_, _03479_);
  or _86946_ (_37208_, _37207_, _03221_);
  or _86947_ (_37209_, _37208_, _37204_);
  nor _86948_ (_37210_, _13237_, _11451_);
  or _86949_ (_37211_, _37210_, _37138_);
  or _86950_ (_37212_, _37211_, _03474_);
  and _86951_ (_37214_, _37212_, _03438_);
  and _86952_ (_37215_, _37214_, _37209_);
  and _86953_ (_37216_, _13244_, _05218_);
  or _86954_ (_37217_, _37216_, _37138_);
  and _86955_ (_37218_, _37217_, _03437_);
  or _86956_ (_37219_, _37218_, _03636_);
  or _86957_ (_37220_, _37219_, _37215_);
  and _86958_ (_37221_, _13253_, _05218_);
  or _86959_ (_37222_, _37221_, _37138_);
  or _86960_ (_37223_, _37222_, _04499_);
  and _86961_ (_37225_, _37223_, _37220_);
  or _86962_ (_37226_, _37225_, _03769_);
  and _86963_ (_37227_, _13259_, _05218_);
  or _86964_ (_37228_, _37227_, _37138_);
  or _86965_ (_37229_, _37228_, _04501_);
  and _86966_ (_37230_, _37229_, _05769_);
  and _86967_ (_37231_, _37230_, _37226_);
  or _86968_ (_37232_, _37138_, _05377_);
  and _86969_ (_37233_, _37217_, _04504_);
  and _86970_ (_37234_, _37233_, _37232_);
  or _86971_ (_37236_, _37234_, _37231_);
  and _86972_ (_37237_, _37236_, _03753_);
  and _86973_ (_37238_, _37152_, _03752_);
  and _86974_ (_37239_, _37238_, _37232_);
  or _86975_ (_37240_, _37239_, _03758_);
  or _86976_ (_37241_, _37240_, _37237_);
  and _86977_ (_37242_, _37241_, _37140_);
  or _86978_ (_37243_, _37242_, _03760_);
  nor _86979_ (_37244_, _13258_, _11451_);
  or _86980_ (_37245_, _37138_, _04517_);
  nor _86981_ (_37247_, _37245_, _37244_);
  nor _86982_ (_37248_, _37247_, _03953_);
  and _86983_ (_37249_, _37248_, _37243_);
  nor _86984_ (_37250_, _37249_, _37135_);
  nor _86985_ (_37251_, _37250_, _03958_);
  and _86986_ (_37252_, _37129_, _03958_);
  or _86987_ (_37253_, _37252_, _03973_);
  or _86988_ (_37254_, _37253_, _37251_);
  not _86989_ (_37255_, _03973_);
  or _86990_ (_37256_, _37129_, _37255_);
  and _86991_ (_37258_, _37256_, _37132_);
  and _86992_ (_37259_, _37258_, _37254_);
  nor _86993_ (_37260_, _37259_, _37134_);
  nor _86994_ (_37261_, _37260_, _04155_);
  and _86995_ (_37262_, _37129_, _04155_);
  or _86996_ (_37263_, _37262_, _36560_);
  or _86997_ (_37264_, _37263_, _37261_);
  or _86998_ (_37265_, _08510_, _08057_);
  or _86999_ (_37266_, _37265_, _36727_);
  and _87000_ (_37267_, _37266_, _04154_);
  and _87001_ (_37269_, _37267_, _37264_);
  and _87002_ (_37270_, _37265_, _04153_);
  or _87003_ (_37271_, _37270_, _03765_);
  or _87004_ (_37272_, _37271_, _37269_);
  or _87005_ (_37273_, _08195_, _03766_);
  or _87006_ (_37274_, _37273_, _08542_);
  and _87007_ (_37275_, _37274_, _08557_);
  and _87008_ (_37276_, _37275_, _37272_);
  or _87009_ (_37277_, _08572_, _08289_);
  and _87010_ (_37278_, _37277_, _08523_);
  or _87011_ (_37280_, _37278_, _15069_);
  or _87012_ (_37281_, _37280_, _37276_);
  or _87013_ (_37282_, _07812_, _07780_);
  and _87014_ (_37283_, _37282_, _07732_);
  and _87015_ (_37284_, _37283_, _37281_);
  and _87016_ (_37285_, _07763_, _07731_);
  or _87017_ (_37286_, _37285_, _03524_);
  or _87018_ (_37287_, _37286_, _37284_);
  or _87019_ (_37288_, _08633_, _03526_);
  and _87020_ (_37289_, _37288_, _08598_);
  and _87021_ (_37291_, _37289_, _37287_);
  and _87022_ (_37292_, _08672_, _08597_);
  or _87023_ (_37293_, _37292_, _03790_);
  or _87024_ (_37294_, _37293_, _37291_);
  or _87025_ (_37295_, _37149_, _04192_);
  and _87026_ (_37296_, _37295_, _03152_);
  and _87027_ (_37297_, _37296_, _37294_);
  and _87028_ (_37298_, _37173_, _03151_);
  or _87029_ (_37299_, _37298_, _03520_);
  or _87030_ (_37300_, _37299_, _37297_);
  and _87031_ (_37302_, _13312_, _05218_);
  or _87032_ (_37303_, _37138_, _03521_);
  or _87033_ (_37304_, _37303_, _37302_);
  and _87034_ (_37305_, _37304_, _42963_);
  and _87035_ (_37306_, _37305_, _37300_);
  or _87036_ (_37307_, _37306_, _37128_);
  and _87037_ (_43396_, _37307_, _41755_);
  and _87038_ (_37308_, _42967_, \oc8051_golden_model_1.P0INREG [0]);
  or _87039_ (_37309_, _37308_, _00816_);
  and _87040_ (_43397_, _37309_, _41755_);
  and _87041_ (_37311_, _42967_, \oc8051_golden_model_1.P0INREG [1]);
  or _87042_ (_37312_, _37311_, _00839_);
  and _87043_ (_43398_, _37312_, _41755_);
  and _87044_ (_37313_, _42967_, \oc8051_golden_model_1.P0INREG [2]);
  or _87045_ (_37314_, _37313_, _00831_);
  and _87046_ (_43399_, _37314_, _41755_);
  and _87047_ (_37315_, _42967_, \oc8051_golden_model_1.P0INREG [3]);
  or _87048_ (_37316_, _37315_, _00824_);
  and _87049_ (_43400_, _37316_, _41755_);
  and _87050_ (_37317_, _42967_, \oc8051_golden_model_1.P0INREG [4]);
  or _87051_ (_37319_, _37317_, _00854_);
  and _87052_ (_43401_, _37319_, _41755_);
  and _87053_ (_37320_, _42967_, \oc8051_golden_model_1.P0INREG [5]);
  or _87054_ (_37321_, _37320_, _00877_);
  and _87055_ (_43402_, _37321_, _41755_);
  and _87056_ (_37322_, _42967_, \oc8051_golden_model_1.P0INREG [6]);
  or _87057_ (_37323_, _37322_, _00870_);
  and _87058_ (_43403_, _37323_, _41755_);
  and _87059_ (_37324_, _42967_, \oc8051_golden_model_1.P1INREG [0]);
  or _87060_ (_37325_, _37324_, _00997_);
  and _87061_ (_43406_, _37325_, _41755_);
  and _87062_ (_37327_, _42967_, \oc8051_golden_model_1.P1INREG [1]);
  or _87063_ (_37328_, _37327_, _01019_);
  and _87064_ (_43407_, _37328_, _41755_);
  and _87065_ (_37329_, _42967_, \oc8051_golden_model_1.P1INREG [2]);
  or _87066_ (_37330_, _37329_, _01012_);
  and _87067_ (_43408_, _37330_, _41755_);
  and _87068_ (_37331_, _42967_, \oc8051_golden_model_1.P1INREG [3]);
  or _87069_ (_37332_, _37331_, _01005_);
  and _87070_ (_43409_, _37332_, _41755_);
  and _87071_ (_37334_, _42967_, \oc8051_golden_model_1.P1INREG [4]);
  or _87072_ (_37335_, _37334_, _00961_);
  and _87073_ (_43410_, _37335_, _41755_);
  and _87074_ (_37336_, _42967_, \oc8051_golden_model_1.P1INREG [5]);
  or _87075_ (_37337_, _37336_, _00983_);
  and _87076_ (_43413_, _37337_, _41755_);
  and _87077_ (_37338_, _42967_, \oc8051_golden_model_1.P1INREG [6]);
  or _87078_ (_37339_, _37338_, _00976_);
  and _87079_ (_43414_, _37339_, _41755_);
  and _87080_ (_37340_, _42967_, \oc8051_golden_model_1.P2INREG [0]);
  or _87081_ (_37342_, _37340_, _00889_);
  and _87082_ (_43415_, _37342_, _41755_);
  and _87083_ (_37343_, _42967_, \oc8051_golden_model_1.P2INREG [1]);
  or _87084_ (_37344_, _37343_, _00905_);
  and _87085_ (_43416_, _37344_, _41755_);
  and _87086_ (_37345_, _42967_, \oc8051_golden_model_1.P2INREG [2]);
  or _87087_ (_37346_, _37345_, _00912_);
  and _87088_ (_43417_, _37346_, _41755_);
  and _87089_ (_37347_, _42967_, \oc8051_golden_model_1.P2INREG [3]);
  or _87090_ (_37348_, _37347_, _00898_);
  and _87091_ (_43418_, _37348_, _41755_);
  and _87092_ (_37350_, _42967_, \oc8051_golden_model_1.P2INREG [4]);
  or _87093_ (_37351_, _37350_, _00926_);
  and _87094_ (_43419_, _37351_, _41755_);
  and _87095_ (_37352_, _42967_, \oc8051_golden_model_1.P2INREG [5]);
  or _87096_ (_37353_, _37352_, _00941_);
  and _87097_ (_43420_, _37353_, _41755_);
  and _87098_ (_37354_, _42967_, \oc8051_golden_model_1.P2INREG [6]);
  or _87099_ (_37355_, _37354_, _00948_);
  and _87100_ (_43421_, _37355_, _41755_);
  and _87101_ (_37357_, _42967_, \oc8051_golden_model_1.P3INREG [0]);
  or _87102_ (_37358_, _37357_, _01072_);
  and _87103_ (_43424_, _37358_, _41755_);
  and _87104_ (_37359_, _42967_, \oc8051_golden_model_1.P3INREG [1]);
  or _87105_ (_37360_, _37359_, _01087_);
  and _87106_ (_43425_, _37360_, _41755_);
  and _87107_ (_37361_, _42967_, \oc8051_golden_model_1.P3INREG [2]);
  or _87108_ (_37362_, _37361_, _01094_);
  and _87109_ (_43426_, _37362_, _41755_);
  and _87110_ (_37363_, _42967_, \oc8051_golden_model_1.P3INREG [3]);
  or _87111_ (_37365_, _37363_, _01080_);
  and _87112_ (_43427_, _37365_, _41755_);
  and _87113_ (_37366_, _42967_, \oc8051_golden_model_1.P3INREG [4]);
  or _87114_ (_37367_, _37366_, _01107_);
  and _87115_ (_43428_, _37367_, _41755_);
  and _87116_ (_37368_, _42967_, \oc8051_golden_model_1.P3INREG [5]);
  or _87117_ (_37369_, _37368_, _01122_);
  and _87118_ (_43429_, _37369_, _41755_);
  and _87119_ (_37370_, _42967_, \oc8051_golden_model_1.P3INREG [6]);
  or _87120_ (_37371_, _37370_, _01129_);
  and _87121_ (_43430_, _37371_, _41755_);
  and _87122_ (_00005_[6], _01130_, _41755_);
  and _87123_ (_00005_[5], _01123_, _41755_);
  and _87124_ (_00005_[4], _01108_, _41755_);
  and _87125_ (_00005_[3], _01081_, _41755_);
  and _87126_ (_00005_[2], _01095_, _41755_);
  and _87127_ (_00005_[1], _01088_, _41755_);
  and _87128_ (_00005_[0], _01073_, _41755_);
  and _87129_ (_00004_[6], _00949_, _41755_);
  and _87130_ (_00004_[5], _00942_, _41755_);
  and _87131_ (_00004_[4], _00927_, _41755_);
  and _87132_ (_00004_[3], _00899_, _41755_);
  and _87133_ (_00004_[2], _00913_, _41755_);
  and _87134_ (_00004_[1], _00906_, _41755_);
  and _87135_ (_00004_[0], _00890_, _41755_);
  and _87136_ (_00003_[6], _00977_, _41755_);
  and _87137_ (_00003_[5], _00984_, _41755_);
  and _87138_ (_00003_[4], _00962_, _41755_);
  and _87139_ (_00003_[3], _01006_, _41755_);
  and _87140_ (_00003_[2], _01013_, _41755_);
  and _87141_ (_00003_[1], _01020_, _41755_);
  and _87142_ (_00003_[0], _00998_, _41755_);
  and _87143_ (_00002_[6], _00871_, _41755_);
  and _87144_ (_00002_[5], _00878_, _41755_);
  and _87145_ (_00002_[4], _00855_, _41755_);
  and _87146_ (_00002_[3], _00825_, _41755_);
  and _87147_ (_00002_[2], _00832_, _41755_);
  and _87148_ (_00002_[1], _00840_, _41755_);
  and _87149_ (_00002_[0], _00817_, _41755_);
  nor _87150_ (_37375_, _09114_, _08918_);
  nor _87151_ (_37377_, _09740_, _09632_);
  and _87152_ (_37378_, _37377_, _37375_);
  not _87153_ (_37379_, _23980_);
  and _87154_ (_37380_, _37379_, _19334_);
  or _87155_ (_37381_, _24452_, _23759_);
  or _87156_ (_37382_, _37381_, _24567_);
  nor _87157_ (_37383_, _37382_, _17915_);
  and _87158_ (_37384_, _37383_, _37380_);
  nor _87159_ (_37385_, _19681_, _18264_);
  nor _87160_ (_37386_, _24336_, _23529_);
  and _87161_ (_37388_, _37386_, _37385_);
  nor _87162_ (_37389_, _17246_, _09522_);
  not _87163_ (_37390_, _18670_);
  and _87164_ (_37391_, _37390_, _17799_);
  and _87165_ (_37392_, _37391_, _37389_);
  nor _87166_ (_37393_, _09441_, _09360_);
  nor _87167_ (_37394_, _09278_, _09196_);
  and _87168_ (_37395_, _37394_, _37393_);
  and _87169_ (_37396_, _37395_, _37392_);
  or _87170_ (_37397_, _23301_, _22528_);
  nor _87171_ (_37399_, _37397_, _24097_);
  nor _87172_ (_37400_, _20684_, _20086_);
  nor _87173_ (_37401_, _21911_, _21289_);
  and _87174_ (_37402_, _37401_, _37400_);
  and _87175_ (_37403_, _37402_, _37399_);
  and _87176_ (_37404_, _37403_, _37396_);
  nand _87177_ (_37405_, _37404_, _37388_);
  nor _87178_ (_37406_, _37405_, _23191_);
  nor _87179_ (_37407_, _19797_, _18497_);
  nor _87180_ (_37408_, _23644_, _19914_);
  and _87181_ (_37410_, _37408_, _37407_);
  nor _87182_ (_37411_, _18147_, _18030_);
  nor _87183_ (_37412_, _22352_, _22263_);
  nor _87184_ (_37413_, _22970_, _22882_);
  and _87185_ (_37414_, _37413_, _37412_);
  nor _87186_ (_37415_, _21117_, _21029_);
  nor _87187_ (_37416_, _21737_, _21648_);
  and _87188_ (_37417_, _37416_, _37415_);
  and _87189_ (_37418_, _37417_, _37414_);
  and _87190_ (_37419_, _37418_, _37411_);
  nor _87191_ (_37421_, _09006_, _08809_);
  nor _87192_ (_37422_, _20854_, _20768_);
  nor _87193_ (_37423_, _20174_, _18759_);
  and _87194_ (_37424_, _37423_, _37422_);
  nor _87195_ (_37425_, _17423_, _17335_);
  nor _87196_ (_37426_, _21198_, _20598_);
  nor _87197_ (_37427_, _22435_, _21819_);
  and _87198_ (_37428_, _37427_, _37426_);
  or _87199_ (_37429_, _03643_, _02945_);
  or _87200_ (_37430_, _37429_, _10534_);
  nor _87201_ (_37432_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor _87202_ (_37433_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and _87203_ (_37434_, _37433_, _37432_);
  nor _87204_ (_37435_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor _87205_ (_37436_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and _87206_ (_37437_, _37436_, _37435_);
  and _87207_ (_37438_, _37437_, _37434_);
  nor _87208_ (_37439_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor _87209_ (_37440_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and _87210_ (_37441_, _37440_, _37439_);
  nor _87211_ (_37443_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor _87212_ (_37444_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and _87213_ (_37445_, _37444_, _37443_);
  and _87214_ (_37446_, _37445_, _37441_);
  and _87215_ (_37447_, _37446_, _37438_);
  nor _87216_ (_37448_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor _87217_ (_37449_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor _87218_ (_37450_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and _87219_ (_37451_, _37450_, _37449_);
  and _87220_ (_37452_, _37451_, _37448_);
  nor _87221_ (_37454_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor _87222_ (_37455_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and _87223_ (_37456_, _37455_, _37454_);
  nor _87224_ (_37457_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor _87225_ (_37458_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and _87226_ (_37459_, _37458_, _37457_);
  and _87227_ (_37460_, _37459_, _37456_);
  and _87228_ (_37461_, _37460_, _37452_);
  and _87229_ (_37462_, _37461_, _37447_);
  nor _87230_ (_37463_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor _87231_ (_37465_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and _87232_ (_37466_, _37465_, _37463_);
  nor _87233_ (_37467_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  nor _87234_ (_37468_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  and _87235_ (_37469_, _37468_, _37467_);
  and _87236_ (_37470_, _37469_, _37466_);
  nor _87237_ (_37471_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor _87238_ (_37472_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and _87239_ (_37473_, _37472_, _37471_);
  nor _87240_ (_37474_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor _87241_ (_37476_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and _87242_ (_37477_, _37476_, _37474_);
  and _87243_ (_37478_, _37477_, _37473_);
  and _87244_ (_37479_, _37478_, _37470_);
  nor _87245_ (_37480_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor _87246_ (_37481_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and _87247_ (_37482_, _37481_, _37480_);
  nor _87248_ (_37483_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor _87249_ (_37484_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and _87250_ (_37485_, _37484_, _37483_);
  and _87251_ (_37487_, _37485_, _37482_);
  nor _87252_ (_37488_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  nor _87253_ (_37489_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  and _87254_ (_37490_, _37489_, _37488_);
  nor _87255_ (_37491_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor _87256_ (_37492_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and _87257_ (_37493_, _37492_, _37491_);
  and _87258_ (_37494_, _37493_, _37490_);
  and _87259_ (_37495_, _37494_, _37487_);
  and _87260_ (_37496_, _37495_, _37479_);
  nor _87261_ (_37498_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and _87262_ (_37499_, _37498_, op0_cnst);
  nor _87263_ (_37500_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor _87264_ (_37501_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and _87265_ (_37502_, _37501_, _37500_);
  nor _87266_ (_37503_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor _87267_ (_37504_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and _87268_ (_37505_, _37504_, _37503_);
  and _87269_ (_37506_, _37505_, _37502_);
  and _87270_ (_37507_, _37506_, _37499_);
  nor _87271_ (_37509_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor _87272_ (_37510_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and _87273_ (_37511_, _37510_, _37509_);
  nor _87274_ (_37512_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor _87275_ (_37513_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and _87276_ (_37514_, _37513_, _37512_);
  and _87277_ (_37515_, _37514_, _37511_);
  and _87278_ (_37516_, \oc8051_golden_model_1.TCON [1], _19117_);
  nor _87279_ (_37517_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and _87280_ (_37518_, _37517_, _37516_);
  nor _87281_ (_37520_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor _87282_ (_37521_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and _87283_ (_37522_, _37521_, _37520_);
  and _87284_ (_37523_, _37522_, _37518_);
  and _87285_ (_37524_, _37523_, _37515_);
  and _87286_ (_37525_, _37524_, _37507_);
  and _87287_ (_37526_, _37525_, _37496_);
  and _87288_ (_37527_, _37526_, _37462_);
  nand _87289_ (_37528_, _37527_, _37430_);
  nor _87290_ (_37529_, _37528_, _17155_);
  nor _87291_ (_37531_, _19994_, _18578_);
  and _87292_ (_37532_, _37531_, _37529_);
  and _87293_ (_37533_, _37532_, _37428_);
  and _87294_ (_37534_, _37533_, _37425_);
  and _87295_ (_37535_, _37534_, _37424_);
  nor _87296_ (_37536_, _22704_, _22617_);
  nor _87297_ (_37537_, _21998_, _21376_);
  and _87298_ (_37538_, _37537_, _37536_);
  and _87299_ (_37539_, _37538_, _23864_);
  and _87300_ (_37540_, _37539_, _37535_);
  nor _87301_ (_37542_, _20942_, _20348_);
  nor _87302_ (_37543_, _21560_, _21465_);
  and _87303_ (_37544_, _37543_, _37542_);
  nor _87304_ (_37545_, _20262_, _18934_);
  nor _87305_ (_37546_, _18847_, _17513_);
  and _87306_ (_37547_, _37546_, _37545_);
  and _87307_ (_37548_, _37547_, _37544_);
  and _87308_ (_37549_, _37548_, _37540_);
  and _87309_ (_37550_, _37549_, _37421_);
  nor _87310_ (_37551_, _19219_, _19113_);
  nor _87311_ (_37553_, _20521_, _20435_);
  and _87312_ (_37554_, _37553_, _37551_);
  nor _87313_ (_37555_, _22174_, _22086_);
  nor _87314_ (_37556_, _23076_, _22793_);
  nand _87315_ (_37557_, _37556_, _37555_);
  nor _87316_ (_37558_, _37557_, _17603_);
  nor _87317_ (_37559_, _19023_, _17692_);
  and _87318_ (_37560_, _37559_, _37558_);
  and _87319_ (_37561_, _37560_, _37554_);
  and _87320_ (_37562_, _37561_, _37550_);
  and _87321_ (_37564_, _37562_, _37419_);
  nor _87322_ (_37565_, _19565_, _19449_);
  nor _87323_ (_37566_, _24216_, _23416_);
  nand _87324_ (_37567_, _37566_, _37565_);
  nor _87325_ (_37568_, _37567_, _18380_);
  and _87326_ (_37569_, _37568_, _37564_);
  and _87327_ (_37570_, _37569_, _37410_);
  and _87328_ (_37571_, _37570_, _37406_);
  and _87329_ (_37572_, _37571_, _37384_);
  and _87330_ (_37573_, _37572_, _37378_);
  or _87331_ (_00001_, _37573_, rst);
  and _87332_ (_00005_[7], _01116_, _41755_);
  and _87333_ (_00004_[7], _00935_, _41755_);
  and _87334_ (_00003_[7], _00970_, _41755_);
  and _87335_ (_00002_[7], _00864_, _41755_);
  and _87336_ (_37575_, _37573_, inst_finished_r);
  nor _87337_ (_37576_, word_in[3], word_in[2]);
  not _87338_ (_37577_, _37576_);
  not _87339_ (_37578_, word_in[1]);
  and _87340_ (_37579_, _37578_, word_in[0]);
  and _87341_ (_37581_, _37579_, \oc8051_golden_model_1.IRAM[1] [0]);
  nor _87342_ (_37582_, _37578_, word_in[0]);
  and _87343_ (_37583_, _37582_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor _87344_ (_37584_, _37583_, _37581_);
  nor _87345_ (_37585_, word_in[1], word_in[0]);
  and _87346_ (_37586_, _37585_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _87347_ (_37587_, word_in[1], word_in[0]);
  and _87348_ (_37588_, _37587_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor _87349_ (_37589_, _37588_, _37586_);
  and _87350_ (_37590_, _37589_, _37584_);
  nor _87351_ (_37592_, _37590_, _37577_);
  not _87352_ (_37593_, word_in[3]);
  nor _87353_ (_37594_, _37593_, word_in[2]);
  not _87354_ (_37595_, _37594_);
  and _87355_ (_37596_, _37579_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _87356_ (_37597_, _37582_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor _87357_ (_37598_, _37597_, _37596_);
  and _87358_ (_37599_, _37585_, \oc8051_golden_model_1.IRAM[8] [0]);
  and _87359_ (_37600_, _37587_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor _87360_ (_37601_, _37600_, _37599_);
  and _87361_ (_37603_, _37601_, _37598_);
  nor _87362_ (_37604_, _37603_, _37595_);
  nor _87363_ (_37605_, _37604_, _37592_);
  and _87364_ (_37606_, _37593_, word_in[2]);
  not _87365_ (_37607_, _37606_);
  and _87366_ (_37608_, _37579_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _87367_ (_37609_, _37582_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor _87368_ (_37610_, _37609_, _37608_);
  and _87369_ (_37611_, _37585_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _87370_ (_37612_, _37587_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor _87371_ (_37614_, _37612_, _37611_);
  and _87372_ (_37615_, _37614_, _37610_);
  nor _87373_ (_37616_, _37615_, _37607_);
  and _87374_ (_37617_, word_in[3], word_in[2]);
  not _87375_ (_37618_, _37617_);
  and _87376_ (_37619_, _37579_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _87377_ (_37620_, _37582_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor _87378_ (_37621_, _37620_, _37619_);
  and _87379_ (_37622_, _37585_, \oc8051_golden_model_1.IRAM[12] [0]);
  and _87380_ (_37623_, _37587_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor _87381_ (_37625_, _37623_, _37622_);
  and _87382_ (_37626_, _37625_, _37621_);
  nor _87383_ (_37627_, _37626_, _37618_);
  nor _87384_ (_37628_, _37627_, _37616_);
  and _87385_ (_37629_, _37628_, _37605_);
  and _87386_ (_37630_, _37617_, _37579_);
  and _87387_ (_37631_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _87388_ (_37632_, _37594_, _37587_);
  and _87389_ (_37633_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _87390_ (_37634_, _37633_, _37631_);
  and _87391_ (_37636_, _37585_, _37606_);
  and _87392_ (_37637_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _87393_ (_37638_, _37576_, _37585_);
  and _87394_ (_37639_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _87395_ (_37640_, _37639_, _37637_);
  and _87396_ (_37641_, _37640_, _37634_);
  and _87397_ (_37642_, _37594_, _37582_);
  and _87398_ (_37643_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _87399_ (_37644_, _37594_, _37579_);
  and _87400_ (_37645_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _87401_ (_37647_, _37645_, _37643_);
  and _87402_ (_37648_, _37617_, _37582_);
  and _87403_ (_37649_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and _87404_ (_37650_, _37617_, _37585_);
  and _87405_ (_37651_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _87406_ (_37652_, _37651_, _37649_);
  and _87407_ (_37653_, _37652_, _37647_);
  and _87408_ (_37654_, _37653_, _37641_);
  and _87409_ (_37655_, _37587_, _37606_);
  and _87410_ (_37656_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and _87411_ (_37658_, _37582_, _37606_);
  and _87412_ (_37659_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor _87413_ (_37660_, _37659_, _37656_);
  and _87414_ (_37661_, _37579_, _37606_);
  and _87415_ (_37662_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and _87416_ (_37663_, _37576_, _37587_);
  and _87417_ (_37664_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _87418_ (_37665_, _37664_, _37662_);
  and _87419_ (_37666_, _37665_, _37660_);
  and _87420_ (_37667_, _37576_, _37582_);
  and _87421_ (_37669_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and _87422_ (_37670_, _37576_, _37579_);
  and _87423_ (_37671_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _87424_ (_37672_, _37671_, _37669_);
  and _87425_ (_37673_, _37617_, _37587_);
  and _87426_ (_37674_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _87427_ (_37675_, _37594_, _37585_);
  and _87428_ (_37676_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _87429_ (_37677_, _37676_, _37674_);
  and _87430_ (_37678_, _37677_, _37672_);
  and _87431_ (_37680_, _37678_, _37666_);
  and _87432_ (_37681_, _37680_, _37654_);
  nand _87433_ (_37682_, _37681_, _37629_);
  or _87434_ (_37683_, _37681_, _37629_);
  and _87435_ (_37684_, _37683_, _37682_);
  and _87436_ (_37685_, _37579_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _87437_ (_37686_, _37582_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor _87438_ (_37687_, _37686_, _37685_);
  and _87439_ (_37688_, _37585_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _87440_ (_37689_, _37587_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor _87441_ (_37691_, _37689_, _37688_);
  and _87442_ (_37692_, _37691_, _37687_);
  nor _87443_ (_37693_, _37692_, _37577_);
  and _87444_ (_37694_, _37579_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _87445_ (_37695_, _37582_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor _87446_ (_37696_, _37695_, _37694_);
  and _87447_ (_37697_, _37585_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _87448_ (_37698_, _37587_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor _87449_ (_37699_, _37698_, _37697_);
  and _87450_ (_37700_, _37699_, _37696_);
  nor _87451_ (_37702_, _37700_, _37618_);
  nor _87452_ (_37703_, _37702_, _37693_);
  and _87453_ (_37704_, _37579_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _87454_ (_37705_, _37582_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor _87455_ (_37706_, _37705_, _37704_);
  and _87456_ (_37707_, _37585_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _87457_ (_37708_, _37587_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor _87458_ (_37709_, _37708_, _37707_);
  and _87459_ (_37710_, _37709_, _37706_);
  nor _87460_ (_37711_, _37710_, _37607_);
  and _87461_ (_37713_, _37579_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _87462_ (_37714_, _37582_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor _87463_ (_37715_, _37714_, _37713_);
  and _87464_ (_37716_, _37585_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _87465_ (_37717_, _37587_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor _87466_ (_37718_, _37717_, _37716_);
  and _87467_ (_37719_, _37718_, _37715_);
  nor _87468_ (_37720_, _37719_, _37595_);
  nor _87469_ (_37721_, _37720_, _37711_);
  and _87470_ (_37722_, _37721_, _37703_);
  and _87471_ (_37724_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _87472_ (_37725_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _87473_ (_37726_, _37725_, _37724_);
  and _87474_ (_37727_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _87475_ (_37728_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _87476_ (_37729_, _37728_, _37727_);
  and _87477_ (_37730_, _37729_, _37726_);
  and _87478_ (_37731_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and _87479_ (_37732_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _87480_ (_37733_, _37732_, _37731_);
  and _87481_ (_37735_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and _87482_ (_37736_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _87483_ (_37737_, _37736_, _37735_);
  and _87484_ (_37738_, _37737_, _37733_);
  and _87485_ (_37739_, _37738_, _37730_);
  and _87486_ (_37740_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _87487_ (_37741_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _87488_ (_37742_, _37741_, _37740_);
  and _87489_ (_37743_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _87490_ (_37744_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _87491_ (_37746_, _37744_, _37743_);
  and _87492_ (_37747_, _37746_, _37742_);
  and _87493_ (_37748_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and _87494_ (_37749_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _87495_ (_37750_, _37749_, _37748_);
  and _87496_ (_37751_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _87497_ (_37752_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor _87498_ (_37753_, _37752_, _37751_);
  and _87499_ (_37754_, _37753_, _37750_);
  and _87500_ (_37755_, _37754_, _37747_);
  and _87501_ (_37757_, _37755_, _37739_);
  nand _87502_ (_37758_, _37757_, _37722_);
  or _87503_ (_37759_, _37757_, _37722_);
  and _87504_ (_37760_, _37759_, _37758_);
  or _87505_ (_37761_, _37760_, _37684_);
  and _87506_ (_37762_, _37579_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _87507_ (_37763_, _37582_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor _87508_ (_37764_, _37763_, _37762_);
  and _87509_ (_37765_, _37585_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _87510_ (_37766_, _37587_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor _87511_ (_37768_, _37766_, _37765_);
  and _87512_ (_37769_, _37768_, _37764_);
  nor _87513_ (_37770_, _37769_, _37607_);
  and _87514_ (_37771_, _37579_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _87515_ (_37772_, _37582_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor _87516_ (_37773_, _37772_, _37771_);
  and _87517_ (_37774_, _37585_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _87518_ (_37775_, _37587_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor _87519_ (_37776_, _37775_, _37774_);
  and _87520_ (_37777_, _37776_, _37773_);
  nor _87521_ (_37779_, _37777_, _37618_);
  nor _87522_ (_37780_, _37779_, _37770_);
  and _87523_ (_37781_, _37579_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _87524_ (_37782_, _37582_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor _87525_ (_37783_, _37782_, _37781_);
  and _87526_ (_37784_, _37585_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _87527_ (_37785_, _37587_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor _87528_ (_37786_, _37785_, _37784_);
  and _87529_ (_37787_, _37786_, _37783_);
  nor _87530_ (_37788_, _37787_, _37577_);
  and _87531_ (_37790_, _37579_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _87532_ (_37791_, _37582_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor _87533_ (_37792_, _37791_, _37790_);
  and _87534_ (_37793_, _37585_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _87535_ (_37794_, _37587_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor _87536_ (_37795_, _37794_, _37793_);
  and _87537_ (_37796_, _37795_, _37792_);
  nor _87538_ (_37797_, _37796_, _37595_);
  nor _87539_ (_37798_, _37797_, _37788_);
  and _87540_ (_37799_, _37798_, _37780_);
  and _87541_ (_37801_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and _87542_ (_37802_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _87543_ (_37803_, _37802_, _37801_);
  and _87544_ (_37804_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _87545_ (_37805_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _87546_ (_37806_, _37805_, _37804_);
  and _87547_ (_37807_, _37806_, _37803_);
  and _87548_ (_37808_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _87549_ (_37809_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _87550_ (_37810_, _37809_, _37808_);
  and _87551_ (_37812_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _87552_ (_37813_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _87553_ (_37814_, _37813_, _37812_);
  and _87554_ (_37815_, _37814_, _37810_);
  and _87555_ (_37816_, _37815_, _37807_);
  and _87556_ (_37817_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _87557_ (_37818_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _87558_ (_37819_, _37818_, _37817_);
  and _87559_ (_37820_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and _87560_ (_37821_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _87561_ (_37823_, _37821_, _37820_);
  and _87562_ (_37824_, _37823_, _37819_);
  and _87563_ (_37825_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _87564_ (_37826_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _87565_ (_37827_, _37826_, _37825_);
  and _87566_ (_37828_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and _87567_ (_37829_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _87568_ (_37830_, _37829_, _37828_);
  and _87569_ (_37831_, _37830_, _37827_);
  and _87570_ (_37832_, _37831_, _37824_);
  and _87571_ (_37834_, _37832_, _37816_);
  nand _87572_ (_37835_, _37834_, _37799_);
  or _87573_ (_37836_, _37834_, _37799_);
  and _87574_ (_37837_, _37836_, _37835_);
  and _87575_ (_37838_, _37579_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _87576_ (_37839_, _37582_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor _87577_ (_37840_, _37839_, _37838_);
  and _87578_ (_37841_, _37585_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _87579_ (_37842_, _37587_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor _87580_ (_37843_, _37842_, _37841_);
  and _87581_ (_37845_, _37843_, _37840_);
  nor _87582_ (_37846_, _37845_, _37607_);
  and _87583_ (_37847_, _37579_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _87584_ (_37848_, _37582_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor _87585_ (_37849_, _37848_, _37847_);
  and _87586_ (_37850_, _37585_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _87587_ (_37851_, _37587_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor _87588_ (_37852_, _37851_, _37850_);
  and _87589_ (_37853_, _37852_, _37849_);
  nor _87590_ (_37854_, _37853_, _37618_);
  nor _87591_ (_37856_, _37854_, _37846_);
  and _87592_ (_37857_, _37579_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _87593_ (_37858_, _37582_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor _87594_ (_37859_, _37858_, _37857_);
  and _87595_ (_37860_, _37585_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _87596_ (_37861_, _37587_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor _87597_ (_37862_, _37861_, _37860_);
  and _87598_ (_37863_, _37862_, _37859_);
  nor _87599_ (_37864_, _37863_, _37577_);
  and _87600_ (_37865_, _37579_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _87601_ (_37867_, _37582_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor _87602_ (_37868_, _37867_, _37865_);
  and _87603_ (_37869_, _37585_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _87604_ (_37870_, _37587_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor _87605_ (_37871_, _37870_, _37869_);
  and _87606_ (_37872_, _37871_, _37868_);
  nor _87607_ (_37873_, _37872_, _37595_);
  nor _87608_ (_37874_, _37873_, _37864_);
  and _87609_ (_37875_, _37874_, _37856_);
  and _87610_ (_37876_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _87611_ (_37878_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _87612_ (_37879_, _37878_, _37876_);
  and _87613_ (_37880_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and _87614_ (_37881_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _87615_ (_37882_, _37881_, _37880_);
  and _87616_ (_37883_, _37882_, _37879_);
  and _87617_ (_37884_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and _87618_ (_37885_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _87619_ (_37886_, _37885_, _37884_);
  and _87620_ (_37887_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _87621_ (_37889_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _87622_ (_37890_, _37889_, _37887_);
  and _87623_ (_37891_, _37890_, _37886_);
  and _87624_ (_37892_, _37891_, _37883_);
  and _87625_ (_37893_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and _87626_ (_37894_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _87627_ (_37895_, _37894_, _37893_);
  and _87628_ (_37896_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and _87629_ (_37897_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _87630_ (_37898_, _37897_, _37896_);
  and _87631_ (_37900_, _37898_, _37895_);
  and _87632_ (_37901_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _87633_ (_37902_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _87634_ (_37903_, _37902_, _37901_);
  and _87635_ (_37904_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and _87636_ (_37905_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _87637_ (_37906_, _37905_, _37904_);
  and _87638_ (_37907_, _37906_, _37903_);
  and _87639_ (_37908_, _37907_, _37900_);
  and _87640_ (_37909_, _37908_, _37892_);
  not _87641_ (_37911_, _37909_);
  nor _87642_ (_37912_, _37911_, _37875_);
  and _87643_ (_37913_, _37911_, _37875_);
  or _87644_ (_37914_, _37913_, _37912_);
  or _87645_ (_37915_, _37914_, _37837_);
  or _87646_ (_37916_, _37915_, _37761_);
  and _87647_ (_37917_, _37579_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _87648_ (_37918_, _37582_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor _87649_ (_37919_, _37918_, _37917_);
  and _87650_ (_37920_, _37585_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _87651_ (_37922_, _37587_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor _87652_ (_37923_, _37922_, _37920_);
  and _87653_ (_37924_, _37923_, _37919_);
  nor _87654_ (_37925_, _37924_, _37577_);
  and _87655_ (_37926_, _37579_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _87656_ (_37927_, _37582_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor _87657_ (_37928_, _37927_, _37926_);
  and _87658_ (_37929_, _37585_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _87659_ (_37930_, _37587_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor _87660_ (_37931_, _37930_, _37929_);
  and _87661_ (_37933_, _37931_, _37928_);
  nor _87662_ (_37934_, _37933_, _37618_);
  nor _87663_ (_37935_, _37934_, _37925_);
  and _87664_ (_37936_, _37579_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _87665_ (_37937_, _37582_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor _87666_ (_37938_, _37937_, _37936_);
  and _87667_ (_37939_, _37585_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _87668_ (_37940_, _37587_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor _87669_ (_37941_, _37940_, _37939_);
  and _87670_ (_37942_, _37941_, _37938_);
  nor _87671_ (_37944_, _37942_, _37607_);
  and _87672_ (_37945_, _37579_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _87673_ (_37946_, _37582_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor _87674_ (_37947_, _37946_, _37945_);
  and _87675_ (_37948_, _37585_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _87676_ (_37949_, _37587_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor _87677_ (_37950_, _37949_, _37948_);
  and _87678_ (_37951_, _37950_, _37947_);
  nor _87679_ (_37952_, _37951_, _37595_);
  nor _87680_ (_37953_, _37952_, _37944_);
  and _87681_ (_37954_, _37953_, _37935_);
  and _87682_ (_37955_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _87683_ (_37956_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _87684_ (_37957_, _37956_, _37955_);
  and _87685_ (_37958_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _87686_ (_37959_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _87687_ (_37960_, _37959_, _37958_);
  and _87688_ (_37961_, _37960_, _37957_);
  and _87689_ (_37962_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _87690_ (_37963_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor _87691_ (_37965_, _37963_, _37962_);
  and _87692_ (_37966_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _87693_ (_37967_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _87694_ (_37968_, _37967_, _37966_);
  and _87695_ (_37969_, _37968_, _37965_);
  and _87696_ (_37970_, _37969_, _37961_);
  and _87697_ (_37971_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _87698_ (_37972_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _87699_ (_37973_, _37972_, _37971_);
  and _87700_ (_37974_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _87701_ (_37976_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _87702_ (_37977_, _37976_, _37974_);
  and _87703_ (_37978_, _37977_, _37973_);
  and _87704_ (_37979_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and _87705_ (_37980_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _87706_ (_37981_, _37980_, _37979_);
  and _87707_ (_37982_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _87708_ (_37983_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _87709_ (_37984_, _37983_, _37982_);
  and _87710_ (_37985_, _37984_, _37981_);
  and _87711_ (_37987_, _37985_, _37978_);
  and _87712_ (_37988_, _37987_, _37970_);
  nand _87713_ (_37989_, _37988_, _37954_);
  or _87714_ (_37990_, _37988_, _37954_);
  and _87715_ (_37991_, _37990_, _37989_);
  and _87716_ (_37992_, _37579_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _87717_ (_37993_, _37582_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor _87718_ (_37994_, _37993_, _37992_);
  and _87719_ (_37995_, _37585_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _87720_ (_37996_, _37587_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor _87721_ (_37998_, _37996_, _37995_);
  and _87722_ (_37999_, _37998_, _37994_);
  nor _87723_ (_38000_, _37999_, _37607_);
  and _87724_ (_38001_, _37579_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _87725_ (_38002_, _37582_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor _87726_ (_38003_, _38002_, _38001_);
  and _87727_ (_38004_, _37585_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _87728_ (_38005_, _37587_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor _87729_ (_38006_, _38005_, _38004_);
  and _87730_ (_38007_, _38006_, _38003_);
  nor _87731_ (_38009_, _38007_, _37595_);
  nor _87732_ (_38010_, _38009_, _38000_);
  and _87733_ (_38011_, _37579_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _87734_ (_38012_, _37582_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor _87735_ (_38013_, _38012_, _38011_);
  and _87736_ (_38014_, _37585_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _87737_ (_38015_, _37587_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor _87738_ (_38016_, _38015_, _38014_);
  and _87739_ (_38017_, _38016_, _38013_);
  nor _87740_ (_38018_, _38017_, _37577_);
  and _87741_ (_38020_, _37579_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _87742_ (_38021_, _37582_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor _87743_ (_38022_, _38021_, _38020_);
  and _87744_ (_38023_, _37585_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _87745_ (_38024_, _37587_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor _87746_ (_38025_, _38024_, _38023_);
  and _87747_ (_38026_, _38025_, _38022_);
  nor _87748_ (_38027_, _38026_, _37618_);
  nor _87749_ (_38028_, _38027_, _38018_);
  and _87750_ (_38029_, _38028_, _38010_);
  and _87751_ (_38031_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _87752_ (_38032_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _87753_ (_38033_, _38032_, _38031_);
  and _87754_ (_38034_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _87755_ (_38035_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _87756_ (_38036_, _38035_, _38034_);
  and _87757_ (_38037_, _38036_, _38033_);
  and _87758_ (_38038_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _87759_ (_38039_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _87760_ (_38040_, _38039_, _38038_);
  and _87761_ (_38042_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _87762_ (_38043_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _87763_ (_38044_, _38043_, _38042_);
  and _87764_ (_38045_, _38044_, _38040_);
  and _87765_ (_38046_, _38045_, _38037_);
  and _87766_ (_38047_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and _87767_ (_38048_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _87768_ (_38049_, _38048_, _38047_);
  and _87769_ (_38050_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and _87770_ (_38051_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _87771_ (_38053_, _38051_, _38050_);
  and _87772_ (_38054_, _38053_, _38049_);
  and _87773_ (_38055_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _87774_ (_38056_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _87775_ (_38057_, _38056_, _38055_);
  and _87776_ (_38058_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and _87777_ (_38059_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor _87778_ (_38060_, _38059_, _38058_);
  and _87779_ (_38061_, _38060_, _38057_);
  and _87780_ (_38062_, _38061_, _38054_);
  and _87781_ (_38064_, _38062_, _38046_);
  not _87782_ (_38065_, _38064_);
  nor _87783_ (_38066_, _38065_, _38029_);
  and _87784_ (_38067_, _38065_, _38029_);
  or _87785_ (_38068_, _38067_, _38066_);
  or _87786_ (_38069_, _38068_, _37991_);
  and _87787_ (_38070_, _37579_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _87788_ (_38071_, _37582_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor _87789_ (_38072_, _38071_, _38070_);
  and _87790_ (_38073_, _37585_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _87791_ (_38075_, _37587_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor _87792_ (_38076_, _38075_, _38073_);
  and _87793_ (_38077_, _38076_, _38072_);
  nor _87794_ (_38078_, _38077_, _37607_);
  and _87795_ (_38079_, _37579_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _87796_ (_38080_, _37582_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor _87797_ (_38081_, _38080_, _38079_);
  and _87798_ (_38082_, _37585_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _87799_ (_38083_, _37587_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor _87800_ (_38084_, _38083_, _38082_);
  and _87801_ (_38086_, _38084_, _38081_);
  nor _87802_ (_38087_, _38086_, _37595_);
  nor _87803_ (_38088_, _38087_, _38078_);
  and _87804_ (_38089_, _37579_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _87805_ (_38090_, _37582_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor _87806_ (_38091_, _38090_, _38089_);
  and _87807_ (_38092_, _37585_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _87808_ (_38093_, _37587_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor _87809_ (_38094_, _38093_, _38092_);
  and _87810_ (_38095_, _38094_, _38091_);
  nor _87811_ (_38097_, _38095_, _37577_);
  and _87812_ (_38098_, _37579_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _87813_ (_38099_, _37582_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor _87814_ (_38100_, _38099_, _38098_);
  and _87815_ (_38101_, _37585_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _87816_ (_38102_, _37587_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor _87817_ (_38103_, _38102_, _38101_);
  and _87818_ (_38104_, _38103_, _38100_);
  nor _87819_ (_38105_, _38104_, _37618_);
  nor _87820_ (_38106_, _38105_, _38097_);
  and _87821_ (_38108_, _38106_, _38088_);
  and _87822_ (_38109_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and _87823_ (_38110_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _87824_ (_38111_, _38110_, _38109_);
  and _87825_ (_38112_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _87826_ (_38113_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _87827_ (_38114_, _38113_, _38112_);
  and _87828_ (_38115_, _38114_, _38111_);
  and _87829_ (_38116_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and _87830_ (_38117_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _87831_ (_38119_, _38117_, _38116_);
  and _87832_ (_38120_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and _87833_ (_38121_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _87834_ (_38122_, _38121_, _38120_);
  and _87835_ (_38123_, _38122_, _38119_);
  and _87836_ (_38124_, _38123_, _38115_);
  and _87837_ (_38125_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and _87838_ (_38126_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _87839_ (_38127_, _38126_, _38125_);
  and _87840_ (_38128_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and _87841_ (_38130_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _87842_ (_38131_, _38130_, _38128_);
  and _87843_ (_38132_, _38131_, _38127_);
  and _87844_ (_38133_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and _87845_ (_38134_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _87846_ (_38135_, _38134_, _38133_);
  and _87847_ (_38136_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _87848_ (_38137_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _87849_ (_38138_, _38137_, _38136_);
  and _87850_ (_38139_, _38138_, _38135_);
  and _87851_ (_38141_, _38139_, _38132_);
  and _87852_ (_38142_, _38141_, _38124_);
  nand _87853_ (_38143_, _38142_, _38108_);
  or _87854_ (_38144_, _38142_, _38108_);
  and _87855_ (_38145_, _38144_, _38143_);
  and _87856_ (_38146_, _37579_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _87857_ (_38147_, _37582_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor _87858_ (_38148_, _38147_, _38146_);
  and _87859_ (_38149_, _37585_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _87860_ (_38150_, _37587_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor _87861_ (_38152_, _38150_, _38149_);
  and _87862_ (_38153_, _38152_, _38148_);
  nor _87863_ (_38154_, _38153_, _37607_);
  and _87864_ (_38155_, _37579_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _87865_ (_38156_, _37582_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor _87866_ (_38157_, _38156_, _38155_);
  and _87867_ (_38158_, _37585_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _87868_ (_38159_, _37587_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor _87869_ (_38160_, _38159_, _38158_);
  and _87870_ (_38161_, _38160_, _38157_);
  nor _87871_ (_38163_, _38161_, _37618_);
  nor _87872_ (_38164_, _38163_, _38154_);
  and _87873_ (_38165_, _37579_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _87874_ (_38166_, _37582_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor _87875_ (_38167_, _38166_, _38165_);
  and _87876_ (_38168_, _37585_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _87877_ (_38169_, _37587_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor _87878_ (_38170_, _38169_, _38168_);
  and _87879_ (_38171_, _38170_, _38167_);
  nor _87880_ (_38172_, _38171_, _37577_);
  and _87881_ (_38174_, _37579_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _87882_ (_38175_, _37582_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor _87883_ (_38176_, _38175_, _38174_);
  and _87884_ (_38177_, _37585_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _87885_ (_38178_, _37587_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor _87886_ (_38179_, _38178_, _38177_);
  and _87887_ (_38180_, _38179_, _38176_);
  nor _87888_ (_38181_, _38180_, _37595_);
  nor _87889_ (_38182_, _38181_, _38172_);
  and _87890_ (_38183_, _38182_, _38164_);
  and _87891_ (_38185_, _37630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _87892_ (_38186_, _37638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _87893_ (_38187_, _38186_, _38185_);
  and _87894_ (_38188_, _37673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _87895_ (_38189_, _37655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor _87896_ (_38190_, _38189_, _38188_);
  and _87897_ (_38191_, _38190_, _38187_);
  and _87898_ (_38192_, _37650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and _87899_ (_38193_, _37675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _87900_ (_38194_, _38193_, _38192_);
  and _87901_ (_38196_, _37644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _87902_ (_38197_, _37663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _87903_ (_38198_, _38197_, _38196_);
  and _87904_ (_38199_, _38198_, _38194_);
  and _87905_ (_38200_, _38199_, _38191_);
  and _87906_ (_38201_, _37632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and _87907_ (_38202_, _37636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _87908_ (_38203_, _38202_, _38201_);
  and _87909_ (_38204_, _37648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and _87910_ (_38205_, _37667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _87911_ (_38207_, _38205_, _38204_);
  and _87912_ (_38208_, _38207_, _38203_);
  and _87913_ (_38209_, _37642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and _87914_ (_38210_, _37661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _87915_ (_38211_, _38210_, _38209_);
  and _87916_ (_38212_, _37658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _87917_ (_38213_, _37670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _87918_ (_38214_, _38213_, _38212_);
  and _87919_ (_38215_, _38214_, _38211_);
  and _87920_ (_38216_, _38215_, _38208_);
  and _87921_ (_38218_, _38216_, _38200_);
  not _87922_ (_38219_, _38218_);
  nor _87923_ (_38220_, _38219_, _38183_);
  and _87924_ (_38221_, _38219_, _38183_);
  or _87925_ (_38222_, _38221_, _38220_);
  or _87926_ (_38223_, _38222_, _38145_);
  or _87927_ (_38224_, _38223_, _38069_);
  or _87928_ (_38225_, _38224_, _37916_);
  and _87929_ (property_invalid_iram, _38225_, _37575_);
  nand _87930_ (_38226_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _87931_ (_38228_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _87932_ (_38229_, _38228_, _38226_);
  and _87933_ (_38230_, _07506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _87934_ (_38231_, _07506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _87935_ (_38232_, _38231_, _38230_);
  or _87936_ (_38233_, _38232_, _38229_);
  nor _87937_ (_38234_, _03233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _87938_ (_38235_, _03233_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _87939_ (_38236_, _38235_, _38234_);
  and _87940_ (_38237_, _03321_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _87941_ (_38239_, _03321_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _87942_ (_38240_, _38239_, _38237_);
  or _87943_ (_38241_, _38240_, _38236_);
  or _87944_ (_38242_, _38241_, _38233_);
  or _87945_ (_38243_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _87946_ (_38244_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _87947_ (_38245_, _38244_, _38243_);
  or _87948_ (_38246_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _87949_ (_38247_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _87950_ (_38248_, _38247_, _38246_);
  or _87951_ (_38250_, _38248_, _38245_);
  and _87952_ (_38251_, _07346_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _87953_ (_38252_, _07346_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _87954_ (_38253_, _38252_, _38251_);
  nand _87955_ (_38254_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _87956_ (_38255_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _87957_ (_38256_, _38255_, _38254_);
  or _87958_ (_38257_, _38256_, _38253_);
  or _87959_ (_38258_, _38257_, _38250_);
  or _87960_ (_38259_, _38258_, _38242_);
  and _87961_ (property_invalid_acc, _38259_, _37575_);
  or _87962_ (_38261_, _26542_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _87963_ (_38262_, _26542_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _87964_ (_38263_, _38262_, _38261_);
  nor _87965_ (_38264_, _27605_, _43884_);
  and _87966_ (_38265_, _28314_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _87967_ (_38266_, _27605_, _43884_);
  or _87968_ (_38267_, _38266_, _38265_);
  or _87969_ (_38268_, _38267_, _38264_);
  nor _87970_ (_38269_, _26901_, _43876_);
  and _87971_ (_38271_, _26901_, _43876_);
  nor _87972_ (_38272_, _28314_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _87973_ (_38273_, _27253_, _43880_);
  nor _87974_ (_38274_, _28666_, _43895_);
  and _87975_ (_38275_, _28666_, _43895_);
  and _87976_ (_38276_, _28997_, _38487_);
  nand _87977_ (_38277_, _30892_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _87978_ (_38278_, _30892_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _87979_ (_38279_, _38278_, _38277_);
  nor _87980_ (_38280_, _29635_, _38498_);
  or _87981_ (_38282_, _26153_, _43869_);
  nand _87982_ (_38283_, _26153_, _43869_);
  and _87983_ (_38284_, _38283_, _38282_);
  and _87984_ (_38285_, _29635_, _38498_);
  or _87985_ (_38286_, _38285_, _38284_);
  or _87986_ (_38287_, _38286_, _38280_);
  nor _87987_ (_38288_, _30264_, _38504_);
  and _87988_ (_38289_, _30264_, _38504_);
  or _87989_ (_38290_, _38289_, _38288_);
  or _87990_ (_38291_, _38290_, _38287_);
  or _87991_ (_38293_, _38291_, _38279_);
  and _87992_ (_38294_, _10868_, _38515_);
  nor _87993_ (_38295_, _10868_, _38515_);
  or _87994_ (_38296_, _38295_, _38294_);
  or _87995_ (_38297_, _38296_, _38293_);
  and _87996_ (_38298_, _29945_, _38483_);
  nor _87997_ (_38299_, _29945_, _38483_);
  or _87998_ (_38300_, _38299_, _38298_);
  nor _87999_ (_38301_, _30581_, _38479_);
  and _88000_ (_38302_, _30581_, _38479_);
  or _88001_ (_38304_, _38302_, _38301_);
  or _88002_ (_38305_, _38304_, _38300_);
  or _88003_ (_38306_, _38305_, _38297_);
  or _88004_ (_38307_, _38306_, _38276_);
  and _88005_ (_38308_, _29327_, _38493_);
  nor _88006_ (_38309_, _28997_, _38487_);
  nor _88007_ (_38310_, _29327_, _38493_);
  or _88008_ (_38311_, _38310_, _38309_);
  or _88009_ (_38312_, _38311_, _38308_);
  or _88010_ (_38313_, _38312_, _38307_);
  or _88011_ (_38315_, _38313_, _38275_);
  or _88012_ (_38316_, _38315_, _38274_);
  or _88013_ (_38317_, _38316_, _38273_);
  nor _88014_ (_38318_, _27965_, _43888_);
  nor _88015_ (_38319_, _27253_, _43880_);
  and _88016_ (_38320_, _27965_, _43888_);
  or _88017_ (_38321_, _38320_, _38319_);
  or _88018_ (_38322_, _38321_, _38318_);
  or _88019_ (_38323_, _38322_, _38317_);
  or _88020_ (_38324_, _38323_, _38272_);
  or _88021_ (_38326_, _38324_, _38271_);
  or _88022_ (_38327_, _38326_, _38269_);
  or _88023_ (_38328_, _38327_, _38268_);
  or _88024_ (_38329_, _38328_, _38263_);
  and _88025_ (_38330_, _37573_, _42963_);
  and _88026_ (property_invalid_pc, _38330_, _38329_);
  buf _88027_ (_01429_, _41755_);
  buf _88028_ (_01481_, _41755_);
  buf _88029_ (_01532_, _41755_);
  buf _88030_ (_01584_, _41755_);
  buf _88031_ (_01623_, _41755_);
  buf _88032_ (_01676_, _41755_);
  buf _88033_ (_01728_, _41755_);
  buf _88034_ (_01780_, _41755_);
  buf _88035_ (_01831_, _41755_);
  buf _88036_ (_01884_, _41755_);
  buf _88037_ (_01936_, _41755_);
  buf _88038_ (_01988_, _41755_);
  buf _88039_ (_02040_, _41755_);
  buf _88040_ (_02092_, _41755_);
  buf _88041_ (_02144_, _41755_);
  buf _88042_ (_02196_, _41755_);
  buf _88043_ (_38864_, _38761_);
  buf _88044_ (_38865_, _38762_);
  buf _88045_ (_38878_, _38761_);
  buf _88046_ (_38879_, _38762_);
  buf _88047_ (_39191_, _38781_);
  buf _88048_ (_39192_, _38783_);
  buf _88049_ (_39193_, _38784_);
  buf _88050_ (_39194_, _38785_);
  buf _88051_ (_39195_, _38786_);
  buf _88052_ (_39196_, _38787_);
  buf _88053_ (_39197_, _38789_);
  buf _88054_ (_39199_, _38790_);
  buf _88055_ (_39200_, _38791_);
  buf _88056_ (_39201_, _38792_);
  buf _88057_ (_39202_, _38793_);
  buf _88058_ (_39203_, _38795_);
  buf _88059_ (_39204_, _38796_);
  buf _88060_ (_39205_, _38797_);
  buf _88061_ (_39257_, _38781_);
  buf _88062_ (_39258_, _38783_);
  buf _88063_ (_39259_, _38784_);
  buf _88064_ (_39260_, _38785_);
  buf _88065_ (_39261_, _38786_);
  buf _88066_ (_39262_, _38787_);
  buf _88067_ (_39263_, _38789_);
  buf _88068_ (_39265_, _38790_);
  buf _88069_ (_39266_, _38791_);
  buf _88070_ (_39267_, _38792_);
  buf _88071_ (_39268_, _38793_);
  buf _88072_ (_39269_, _38795_);
  buf _88073_ (_39270_, _38796_);
  buf _88074_ (_39271_, _38797_);
  buf _88075_ (_39597_, _39563_);
  buf _88076_ (_39711_, _39563_);
  dff _88077_ (p0in_reg[0], _00002_[0], clk);
  dff _88078_ (p0in_reg[1], _00002_[1], clk);
  dff _88079_ (p0in_reg[2], _00002_[2], clk);
  dff _88080_ (p0in_reg[3], _00002_[3], clk);
  dff _88081_ (p0in_reg[4], _00002_[4], clk);
  dff _88082_ (p0in_reg[5], _00002_[5], clk);
  dff _88083_ (p0in_reg[6], _00002_[6], clk);
  dff _88084_ (p0in_reg[7], _00002_[7], clk);
  dff _88085_ (p1in_reg[0], _00003_[0], clk);
  dff _88086_ (p1in_reg[1], _00003_[1], clk);
  dff _88087_ (p1in_reg[2], _00003_[2], clk);
  dff _88088_ (p1in_reg[3], _00003_[3], clk);
  dff _88089_ (p1in_reg[4], _00003_[4], clk);
  dff _88090_ (p1in_reg[5], _00003_[5], clk);
  dff _88091_ (p1in_reg[6], _00003_[6], clk);
  dff _88092_ (p1in_reg[7], _00003_[7], clk);
  dff _88093_ (p2in_reg[0], _00004_[0], clk);
  dff _88094_ (p2in_reg[1], _00004_[1], clk);
  dff _88095_ (p2in_reg[2], _00004_[2], clk);
  dff _88096_ (p2in_reg[3], _00004_[3], clk);
  dff _88097_ (p2in_reg[4], _00004_[4], clk);
  dff _88098_ (p2in_reg[5], _00004_[5], clk);
  dff _88099_ (p2in_reg[6], _00004_[6], clk);
  dff _88100_ (p2in_reg[7], _00004_[7], clk);
  dff _88101_ (p3in_reg[0], _00005_[0], clk);
  dff _88102_ (p3in_reg[1], _00005_[1], clk);
  dff _88103_ (p3in_reg[2], _00005_[2], clk);
  dff _88104_ (p3in_reg[3], _00005_[3], clk);
  dff _88105_ (p3in_reg[4], _00005_[4], clk);
  dff _88106_ (p3in_reg[5], _00005_[5], clk);
  dff _88107_ (p3in_reg[6], _00005_[6], clk);
  dff _88108_ (p3in_reg[7], _00005_[7], clk);
  dff _88109_ (op0_cnst, _00001_, clk);
  dff _88110_ (inst_finished_r, _00000_, clk);
  dff _88111_ (\oc8051_gm_cxrom_1.cell0.data [0], _01433_, clk);
  dff _88112_ (\oc8051_gm_cxrom_1.cell0.data [1], _01437_, clk);
  dff _88113_ (\oc8051_gm_cxrom_1.cell0.data [2], _01441_, clk);
  dff _88114_ (\oc8051_gm_cxrom_1.cell0.data [3], _01445_, clk);
  dff _88115_ (\oc8051_gm_cxrom_1.cell0.data [4], _01449_, clk);
  dff _88116_ (\oc8051_gm_cxrom_1.cell0.data [5], _01453_, clk);
  dff _88117_ (\oc8051_gm_cxrom_1.cell0.data [6], _01457_, clk);
  dff _88118_ (\oc8051_gm_cxrom_1.cell0.data [7], _01426_, clk);
  dff _88119_ (\oc8051_gm_cxrom_1.cell0.valid , _01429_, clk);
  dff _88120_ (\oc8051_gm_cxrom_1.cell1.data [0], _01485_, clk);
  dff _88121_ (\oc8051_gm_cxrom_1.cell1.data [1], _01489_, clk);
  dff _88122_ (\oc8051_gm_cxrom_1.cell1.data [2], _01493_, clk);
  dff _88123_ (\oc8051_gm_cxrom_1.cell1.data [3], _01496_, clk);
  dff _88124_ (\oc8051_gm_cxrom_1.cell1.data [4], _01500_, clk);
  dff _88125_ (\oc8051_gm_cxrom_1.cell1.data [5], _01504_, clk);
  dff _88126_ (\oc8051_gm_cxrom_1.cell1.data [6], _01508_, clk);
  dff _88127_ (\oc8051_gm_cxrom_1.cell1.data [7], _01478_, clk);
  dff _88128_ (\oc8051_gm_cxrom_1.cell1.valid , _01481_, clk);
  dff _88129_ (\oc8051_gm_cxrom_1.cell10.data [0], _01940_, clk);
  dff _88130_ (\oc8051_gm_cxrom_1.cell10.data [1], _01943_, clk);
  dff _88131_ (\oc8051_gm_cxrom_1.cell10.data [2], _01947_, clk);
  dff _88132_ (\oc8051_gm_cxrom_1.cell10.data [3], _01951_, clk);
  dff _88133_ (\oc8051_gm_cxrom_1.cell10.data [4], _01955_, clk);
  dff _88134_ (\oc8051_gm_cxrom_1.cell10.data [5], _01959_, clk);
  dff _88135_ (\oc8051_gm_cxrom_1.cell10.data [6], _01963_, clk);
  dff _88136_ (\oc8051_gm_cxrom_1.cell10.data [7], _01933_, clk);
  dff _88137_ (\oc8051_gm_cxrom_1.cell10.valid , _01936_, clk);
  dff _88138_ (\oc8051_gm_cxrom_1.cell11.data [0], _01992_, clk);
  dff _88139_ (\oc8051_gm_cxrom_1.cell11.data [1], _01996_, clk);
  dff _88140_ (\oc8051_gm_cxrom_1.cell11.data [2], _01999_, clk);
  dff _88141_ (\oc8051_gm_cxrom_1.cell11.data [3], _02003_, clk);
  dff _88142_ (\oc8051_gm_cxrom_1.cell11.data [4], _02007_, clk);
  dff _88143_ (\oc8051_gm_cxrom_1.cell11.data [5], _02011_, clk);
  dff _88144_ (\oc8051_gm_cxrom_1.cell11.data [6], _02015_, clk);
  dff _88145_ (\oc8051_gm_cxrom_1.cell11.data [7], _01985_, clk);
  dff _88146_ (\oc8051_gm_cxrom_1.cell11.valid , _01988_, clk);
  dff _88147_ (\oc8051_gm_cxrom_1.cell12.data [0], _02044_, clk);
  dff _88148_ (\oc8051_gm_cxrom_1.cell12.data [1], _02048_, clk);
  dff _88149_ (\oc8051_gm_cxrom_1.cell12.data [2], _02052_, clk);
  dff _88150_ (\oc8051_gm_cxrom_1.cell12.data [3], _02055_, clk);
  dff _88151_ (\oc8051_gm_cxrom_1.cell12.data [4], _02059_, clk);
  dff _88152_ (\oc8051_gm_cxrom_1.cell12.data [5], _02063_, clk);
  dff _88153_ (\oc8051_gm_cxrom_1.cell12.data [6], _02067_, clk);
  dff _88154_ (\oc8051_gm_cxrom_1.cell12.data [7], _02037_, clk);
  dff _88155_ (\oc8051_gm_cxrom_1.cell12.valid , _02040_, clk);
  dff _88156_ (\oc8051_gm_cxrom_1.cell13.data [0], _02096_, clk);
  dff _88157_ (\oc8051_gm_cxrom_1.cell13.data [1], _02100_, clk);
  dff _88158_ (\oc8051_gm_cxrom_1.cell13.data [2], _02104_, clk);
  dff _88159_ (\oc8051_gm_cxrom_1.cell13.data [3], _02108_, clk);
  dff _88160_ (\oc8051_gm_cxrom_1.cell13.data [4], _02111_, clk);
  dff _88161_ (\oc8051_gm_cxrom_1.cell13.data [5], _02115_, clk);
  dff _88162_ (\oc8051_gm_cxrom_1.cell13.data [6], _02119_, clk);
  dff _88163_ (\oc8051_gm_cxrom_1.cell13.data [7], _02089_, clk);
  dff _88164_ (\oc8051_gm_cxrom_1.cell13.valid , _02092_, clk);
  dff _88165_ (\oc8051_gm_cxrom_1.cell14.data [0], _02148_, clk);
  dff _88166_ (\oc8051_gm_cxrom_1.cell14.data [1], _02152_, clk);
  dff _88167_ (\oc8051_gm_cxrom_1.cell14.data [2], _02156_, clk);
  dff _88168_ (\oc8051_gm_cxrom_1.cell14.data [3], _02160_, clk);
  dff _88169_ (\oc8051_gm_cxrom_1.cell14.data [4], _02164_, clk);
  dff _88170_ (\oc8051_gm_cxrom_1.cell14.data [5], _02167_, clk);
  dff _88171_ (\oc8051_gm_cxrom_1.cell14.data [6], _02171_, clk);
  dff _88172_ (\oc8051_gm_cxrom_1.cell14.data [7], _02141_, clk);
  dff _88173_ (\oc8051_gm_cxrom_1.cell14.valid , _02144_, clk);
  dff _88174_ (\oc8051_gm_cxrom_1.cell15.data [0], _02200_, clk);
  dff _88175_ (\oc8051_gm_cxrom_1.cell15.data [1], _02204_, clk);
  dff _88176_ (\oc8051_gm_cxrom_1.cell15.data [2], _02208_, clk);
  dff _88177_ (\oc8051_gm_cxrom_1.cell15.data [3], _02212_, clk);
  dff _88178_ (\oc8051_gm_cxrom_1.cell15.data [4], _02216_, clk);
  dff _88179_ (\oc8051_gm_cxrom_1.cell15.data [5], _02220_, clk);
  dff _88180_ (\oc8051_gm_cxrom_1.cell15.data [6], _02223_, clk);
  dff _88181_ (\oc8051_gm_cxrom_1.cell15.data [7], _02193_, clk);
  dff _88182_ (\oc8051_gm_cxrom_1.cell15.valid , _02196_, clk);
  dff _88183_ (\oc8051_gm_cxrom_1.cell2.data [0], _01536_, clk);
  dff _88184_ (\oc8051_gm_cxrom_1.cell2.data [1], _01540_, clk);
  dff _88185_ (\oc8051_gm_cxrom_1.cell2.data [2], _01544_, clk);
  dff _88186_ (\oc8051_gm_cxrom_1.cell2.data [3], _01548_, clk);
  dff _88187_ (\oc8051_gm_cxrom_1.cell2.data [4], _01552_, clk);
  dff _88188_ (\oc8051_gm_cxrom_1.cell2.data [5], _01556_, clk);
  dff _88189_ (\oc8051_gm_cxrom_1.cell2.data [6], _01560_, clk);
  dff _88190_ (\oc8051_gm_cxrom_1.cell2.data [7], _01529_, clk);
  dff _88191_ (\oc8051_gm_cxrom_1.cell2.valid , _01532_, clk);
  dff _88192_ (\oc8051_gm_cxrom_1.cell3.data [0], _01588_, clk);
  dff _88193_ (\oc8051_gm_cxrom_1.cell3.data [1], _01592_, clk);
  dff _88194_ (\oc8051_gm_cxrom_1.cell3.data [2], _01596_, clk);
  dff _88195_ (\oc8051_gm_cxrom_1.cell3.data [3], _01600_, clk);
  dff _88196_ (\oc8051_gm_cxrom_1.cell3.data [4], _01604_, clk);
  dff _88197_ (\oc8051_gm_cxrom_1.cell3.data [5], _01607_, clk);
  dff _88198_ (\oc8051_gm_cxrom_1.cell3.data [6], _01608_, clk);
  dff _88199_ (\oc8051_gm_cxrom_1.cell3.data [7], _01581_, clk);
  dff _88200_ (\oc8051_gm_cxrom_1.cell3.valid , _01584_, clk);
  dff _88201_ (\oc8051_gm_cxrom_1.cell4.data [0], _01627_, clk);
  dff _88202_ (\oc8051_gm_cxrom_1.cell4.data [1], _01631_, clk);
  dff _88203_ (\oc8051_gm_cxrom_1.cell4.data [2], _01635_, clk);
  dff _88204_ (\oc8051_gm_cxrom_1.cell4.data [3], _01639_, clk);
  dff _88205_ (\oc8051_gm_cxrom_1.cell4.data [4], _01643_, clk);
  dff _88206_ (\oc8051_gm_cxrom_1.cell4.data [5], _01647_, clk);
  dff _88207_ (\oc8051_gm_cxrom_1.cell4.data [6], _01651_, clk);
  dff _88208_ (\oc8051_gm_cxrom_1.cell4.data [7], _01620_, clk);
  dff _88209_ (\oc8051_gm_cxrom_1.cell4.valid , _01623_, clk);
  dff _88210_ (\oc8051_gm_cxrom_1.cell5.data [0], _01680_, clk);
  dff _88211_ (\oc8051_gm_cxrom_1.cell5.data [1], _01684_, clk);
  dff _88212_ (\oc8051_gm_cxrom_1.cell5.data [2], _01688_, clk);
  dff _88213_ (\oc8051_gm_cxrom_1.cell5.data [3], _01692_, clk);
  dff _88214_ (\oc8051_gm_cxrom_1.cell5.data [4], _01696_, clk);
  dff _88215_ (\oc8051_gm_cxrom_1.cell5.data [5], _01700_, clk);
  dff _88216_ (\oc8051_gm_cxrom_1.cell5.data [6], _01704_, clk);
  dff _88217_ (\oc8051_gm_cxrom_1.cell5.data [7], _01673_, clk);
  dff _88218_ (\oc8051_gm_cxrom_1.cell5.valid , _01676_, clk);
  dff _88219_ (\oc8051_gm_cxrom_1.cell6.data [0], _01732_, clk);
  dff _88220_ (\oc8051_gm_cxrom_1.cell6.data [1], _01736_, clk);
  dff _88221_ (\oc8051_gm_cxrom_1.cell6.data [2], _01740_, clk);
  dff _88222_ (\oc8051_gm_cxrom_1.cell6.data [3], _01744_, clk);
  dff _88223_ (\oc8051_gm_cxrom_1.cell6.data [4], _01748_, clk);
  dff _88224_ (\oc8051_gm_cxrom_1.cell6.data [5], _01752_, clk);
  dff _88225_ (\oc8051_gm_cxrom_1.cell6.data [6], _01756_, clk);
  dff _88226_ (\oc8051_gm_cxrom_1.cell6.data [7], _01725_, clk);
  dff _88227_ (\oc8051_gm_cxrom_1.cell6.valid , _01728_, clk);
  dff _88228_ (\oc8051_gm_cxrom_1.cell7.data [0], _01784_, clk);
  dff _88229_ (\oc8051_gm_cxrom_1.cell7.data [1], _01788_, clk);
  dff _88230_ (\oc8051_gm_cxrom_1.cell7.data [2], _01792_, clk);
  dff _88231_ (\oc8051_gm_cxrom_1.cell7.data [3], _01795_, clk);
  dff _88232_ (\oc8051_gm_cxrom_1.cell7.data [4], _01799_, clk);
  dff _88233_ (\oc8051_gm_cxrom_1.cell7.data [5], _01803_, clk);
  dff _88234_ (\oc8051_gm_cxrom_1.cell7.data [6], _01807_, clk);
  dff _88235_ (\oc8051_gm_cxrom_1.cell7.data [7], _01777_, clk);
  dff _88236_ (\oc8051_gm_cxrom_1.cell7.valid , _01780_, clk);
  dff _88237_ (\oc8051_gm_cxrom_1.cell8.data [0], _01835_, clk);
  dff _88238_ (\oc8051_gm_cxrom_1.cell8.data [1], _01839_, clk);
  dff _88239_ (\oc8051_gm_cxrom_1.cell8.data [2], _01843_, clk);
  dff _88240_ (\oc8051_gm_cxrom_1.cell8.data [3], _01847_, clk);
  dff _88241_ (\oc8051_gm_cxrom_1.cell8.data [4], _01851_, clk);
  dff _88242_ (\oc8051_gm_cxrom_1.cell8.data [5], _01855_, clk);
  dff _88243_ (\oc8051_gm_cxrom_1.cell8.data [6], _01859_, clk);
  dff _88244_ (\oc8051_gm_cxrom_1.cell8.data [7], _01828_, clk);
  dff _88245_ (\oc8051_gm_cxrom_1.cell8.valid , _01831_, clk);
  dff _88246_ (\oc8051_gm_cxrom_1.cell9.data [0], _01887_, clk);
  dff _88247_ (\oc8051_gm_cxrom_1.cell9.data [1], _01891_, clk);
  dff _88248_ (\oc8051_gm_cxrom_1.cell9.data [2], _01895_, clk);
  dff _88249_ (\oc8051_gm_cxrom_1.cell9.data [3], _01899_, clk);
  dff _88250_ (\oc8051_gm_cxrom_1.cell9.data [4], _01903_, clk);
  dff _88251_ (\oc8051_gm_cxrom_1.cell9.data [5], _01907_, clk);
  dff _88252_ (\oc8051_gm_cxrom_1.cell9.data [6], _01911_, clk);
  dff _88253_ (\oc8051_gm_cxrom_1.cell9.data [7], _01881_, clk);
  dff _88254_ (\oc8051_gm_cxrom_1.cell9.valid , _01884_, clk);
  dff _88255_ (\oc8051_golden_model_1.IRAM[15] [0], _40746_, clk);
  dff _88256_ (\oc8051_golden_model_1.IRAM[15] [1], _40747_, clk);
  dff _88257_ (\oc8051_golden_model_1.IRAM[15] [2], _40748_, clk);
  dff _88258_ (\oc8051_golden_model_1.IRAM[15] [3], _40749_, clk);
  dff _88259_ (\oc8051_golden_model_1.IRAM[15] [4], _40751_, clk);
  dff _88260_ (\oc8051_golden_model_1.IRAM[15] [5], _40752_, clk);
  dff _88261_ (\oc8051_golden_model_1.IRAM[15] [6], _40753_, clk);
  dff _88262_ (\oc8051_golden_model_1.IRAM[15] [7], _40514_, clk);
  dff _88263_ (\oc8051_golden_model_1.IRAM[14] [0], _40734_, clk);
  dff _88264_ (\oc8051_golden_model_1.IRAM[14] [1], _40735_, clk);
  dff _88265_ (\oc8051_golden_model_1.IRAM[14] [2], _40736_, clk);
  dff _88266_ (\oc8051_golden_model_1.IRAM[14] [3], _40737_, clk);
  dff _88267_ (\oc8051_golden_model_1.IRAM[14] [4], _40739_, clk);
  dff _88268_ (\oc8051_golden_model_1.IRAM[14] [5], _40740_, clk);
  dff _88269_ (\oc8051_golden_model_1.IRAM[14] [6], _40741_, clk);
  dff _88270_ (\oc8051_golden_model_1.IRAM[14] [7], _40742_, clk);
  dff _88271_ (\oc8051_golden_model_1.IRAM[13] [0], _40722_, clk);
  dff _88272_ (\oc8051_golden_model_1.IRAM[13] [1], _40723_, clk);
  dff _88273_ (\oc8051_golden_model_1.IRAM[13] [2], _40724_, clk);
  dff _88274_ (\oc8051_golden_model_1.IRAM[13] [3], _40725_, clk);
  dff _88275_ (\oc8051_golden_model_1.IRAM[13] [4], _40727_, clk);
  dff _88276_ (\oc8051_golden_model_1.IRAM[13] [5], _40728_, clk);
  dff _88277_ (\oc8051_golden_model_1.IRAM[13] [6], _40729_, clk);
  dff _88278_ (\oc8051_golden_model_1.IRAM[13] [7], _40730_, clk);
  dff _88279_ (\oc8051_golden_model_1.IRAM[12] [0], _40710_, clk);
  dff _88280_ (\oc8051_golden_model_1.IRAM[12] [1], _40711_, clk);
  dff _88281_ (\oc8051_golden_model_1.IRAM[12] [2], _40712_, clk);
  dff _88282_ (\oc8051_golden_model_1.IRAM[12] [3], _40713_, clk);
  dff _88283_ (\oc8051_golden_model_1.IRAM[12] [4], _40714_, clk);
  dff _88284_ (\oc8051_golden_model_1.IRAM[12] [5], _40716_, clk);
  dff _88285_ (\oc8051_golden_model_1.IRAM[12] [6], _40717_, clk);
  dff _88286_ (\oc8051_golden_model_1.IRAM[12] [7], _40718_, clk);
  dff _88287_ (\oc8051_golden_model_1.IRAM[11] [0], _40697_, clk);
  dff _88288_ (\oc8051_golden_model_1.IRAM[11] [1], _40699_, clk);
  dff _88289_ (\oc8051_golden_model_1.IRAM[11] [2], _40700_, clk);
  dff _88290_ (\oc8051_golden_model_1.IRAM[11] [3], _40701_, clk);
  dff _88291_ (\oc8051_golden_model_1.IRAM[11] [4], _40702_, clk);
  dff _88292_ (\oc8051_golden_model_1.IRAM[11] [5], _40703_, clk);
  dff _88293_ (\oc8051_golden_model_1.IRAM[11] [6], _40705_, clk);
  dff _88294_ (\oc8051_golden_model_1.IRAM[11] [7], _40706_, clk);
  dff _88295_ (\oc8051_golden_model_1.IRAM[10] [0], _40685_, clk);
  dff _88296_ (\oc8051_golden_model_1.IRAM[10] [1], _40686_, clk);
  dff _88297_ (\oc8051_golden_model_1.IRAM[10] [2], _40688_, clk);
  dff _88298_ (\oc8051_golden_model_1.IRAM[10] [3], _40689_, clk);
  dff _88299_ (\oc8051_golden_model_1.IRAM[10] [4], _40690_, clk);
  dff _88300_ (\oc8051_golden_model_1.IRAM[10] [5], _40691_, clk);
  dff _88301_ (\oc8051_golden_model_1.IRAM[10] [6], _40692_, clk);
  dff _88302_ (\oc8051_golden_model_1.IRAM[10] [7], _40694_, clk);
  dff _88303_ (\oc8051_golden_model_1.IRAM[9] [0], _40673_, clk);
  dff _88304_ (\oc8051_golden_model_1.IRAM[9] [1], _40674_, clk);
  dff _88305_ (\oc8051_golden_model_1.IRAM[9] [2], _40676_, clk);
  dff _88306_ (\oc8051_golden_model_1.IRAM[9] [3], _40677_, clk);
  dff _88307_ (\oc8051_golden_model_1.IRAM[9] [4], _40678_, clk);
  dff _88308_ (\oc8051_golden_model_1.IRAM[9] [5], _40679_, clk);
  dff _88309_ (\oc8051_golden_model_1.IRAM[9] [6], _40680_, clk);
  dff _88310_ (\oc8051_golden_model_1.IRAM[9] [7], _40682_, clk);
  dff _88311_ (\oc8051_golden_model_1.IRAM[8] [0], _40661_, clk);
  dff _88312_ (\oc8051_golden_model_1.IRAM[8] [1], _40662_, clk);
  dff _88313_ (\oc8051_golden_model_1.IRAM[8] [2], _40663_, clk);
  dff _88314_ (\oc8051_golden_model_1.IRAM[8] [3], _40665_, clk);
  dff _88315_ (\oc8051_golden_model_1.IRAM[8] [4], _40666_, clk);
  dff _88316_ (\oc8051_golden_model_1.IRAM[8] [5], _40667_, clk);
  dff _88317_ (\oc8051_golden_model_1.IRAM[8] [6], _40668_, clk);
  dff _88318_ (\oc8051_golden_model_1.IRAM[8] [7], _40669_, clk);
  dff _88319_ (\oc8051_golden_model_1.IRAM[7] [0], _40648_, clk);
  dff _88320_ (\oc8051_golden_model_1.IRAM[7] [1], _40650_, clk);
  dff _88321_ (\oc8051_golden_model_1.IRAM[7] [2], _40651_, clk);
  dff _88322_ (\oc8051_golden_model_1.IRAM[7] [3], _40652_, clk);
  dff _88323_ (\oc8051_golden_model_1.IRAM[7] [4], _40653_, clk);
  dff _88324_ (\oc8051_golden_model_1.IRAM[7] [5], _40654_, clk);
  dff _88325_ (\oc8051_golden_model_1.IRAM[7] [6], _40656_, clk);
  dff _88326_ (\oc8051_golden_model_1.IRAM[7] [7], _40657_, clk);
  dff _88327_ (\oc8051_golden_model_1.IRAM[6] [0], _40636_, clk);
  dff _88328_ (\oc8051_golden_model_1.IRAM[6] [1], _40637_, clk);
  dff _88329_ (\oc8051_golden_model_1.IRAM[6] [2], _40639_, clk);
  dff _88330_ (\oc8051_golden_model_1.IRAM[6] [3], _40640_, clk);
  dff _88331_ (\oc8051_golden_model_1.IRAM[6] [4], _40641_, clk);
  dff _88332_ (\oc8051_golden_model_1.IRAM[6] [5], _40642_, clk);
  dff _88333_ (\oc8051_golden_model_1.IRAM[6] [6], _40643_, clk);
  dff _88334_ (\oc8051_golden_model_1.IRAM[6] [7], _40645_, clk);
  dff _88335_ (\oc8051_golden_model_1.IRAM[5] [0], _40624_, clk);
  dff _88336_ (\oc8051_golden_model_1.IRAM[5] [1], _40625_, clk);
  dff _88337_ (\oc8051_golden_model_1.IRAM[5] [2], _40627_, clk);
  dff _88338_ (\oc8051_golden_model_1.IRAM[5] [3], _40628_, clk);
  dff _88339_ (\oc8051_golden_model_1.IRAM[5] [4], _40629_, clk);
  dff _88340_ (\oc8051_golden_model_1.IRAM[5] [5], _40630_, clk);
  dff _88341_ (\oc8051_golden_model_1.IRAM[5] [6], _40631_, clk);
  dff _88342_ (\oc8051_golden_model_1.IRAM[5] [7], _40633_, clk);
  dff _88343_ (\oc8051_golden_model_1.IRAM[4] [0], _40612_, clk);
  dff _88344_ (\oc8051_golden_model_1.IRAM[4] [1], _40613_, clk);
  dff _88345_ (\oc8051_golden_model_1.IRAM[4] [2], _40614_, clk);
  dff _88346_ (\oc8051_golden_model_1.IRAM[4] [3], _40616_, clk);
  dff _88347_ (\oc8051_golden_model_1.IRAM[4] [4], _40617_, clk);
  dff _88348_ (\oc8051_golden_model_1.IRAM[4] [5], _40618_, clk);
  dff _88349_ (\oc8051_golden_model_1.IRAM[4] [6], _40619_, clk);
  dff _88350_ (\oc8051_golden_model_1.IRAM[4] [7], _40620_, clk);
  dff _88351_ (\oc8051_golden_model_1.IRAM[3] [0], _40599_, clk);
  dff _88352_ (\oc8051_golden_model_1.IRAM[3] [1], _40601_, clk);
  dff _88353_ (\oc8051_golden_model_1.IRAM[3] [2], _40602_, clk);
  dff _88354_ (\oc8051_golden_model_1.IRAM[3] [3], _40603_, clk);
  dff _88355_ (\oc8051_golden_model_1.IRAM[3] [4], _40604_, clk);
  dff _88356_ (\oc8051_golden_model_1.IRAM[3] [5], _40605_, clk);
  dff _88357_ (\oc8051_golden_model_1.IRAM[3] [6], _40607_, clk);
  dff _88358_ (\oc8051_golden_model_1.IRAM[3] [7], _40608_, clk);
  dff _88359_ (\oc8051_golden_model_1.IRAM[2] [0], _40587_, clk);
  dff _88360_ (\oc8051_golden_model_1.IRAM[2] [1], _40588_, clk);
  dff _88361_ (\oc8051_golden_model_1.IRAM[2] [2], _40589_, clk);
  dff _88362_ (\oc8051_golden_model_1.IRAM[2] [3], _40591_, clk);
  dff _88363_ (\oc8051_golden_model_1.IRAM[2] [4], _40592_, clk);
  dff _88364_ (\oc8051_golden_model_1.IRAM[2] [5], _40593_, clk);
  dff _88365_ (\oc8051_golden_model_1.IRAM[2] [6], _40594_, clk);
  dff _88366_ (\oc8051_golden_model_1.IRAM[2] [7], _40595_, clk);
  dff _88367_ (\oc8051_golden_model_1.IRAM[1] [0], _40574_, clk);
  dff _88368_ (\oc8051_golden_model_1.IRAM[1] [1], _40576_, clk);
  dff _88369_ (\oc8051_golden_model_1.IRAM[1] [2], _40577_, clk);
  dff _88370_ (\oc8051_golden_model_1.IRAM[1] [3], _40578_, clk);
  dff _88371_ (\oc8051_golden_model_1.IRAM[1] [4], _40579_, clk);
  dff _88372_ (\oc8051_golden_model_1.IRAM[1] [5], _40580_, clk);
  dff _88373_ (\oc8051_golden_model_1.IRAM[1] [6], _40582_, clk);
  dff _88374_ (\oc8051_golden_model_1.IRAM[1] [7], _40583_, clk);
  dff _88375_ (\oc8051_golden_model_1.IRAM[0] [0], _40560_, clk);
  dff _88376_ (\oc8051_golden_model_1.IRAM[0] [1], _40562_, clk);
  dff _88377_ (\oc8051_golden_model_1.IRAM[0] [2], _40563_, clk);
  dff _88378_ (\oc8051_golden_model_1.IRAM[0] [3], _40565_, clk);
  dff _88379_ (\oc8051_golden_model_1.IRAM[0] [4], _40566_, clk);
  dff _88380_ (\oc8051_golden_model_1.IRAM[0] [5], _40567_, clk);
  dff _88381_ (\oc8051_golden_model_1.IRAM[0] [6], _40569_, clk);
  dff _88382_ (\oc8051_golden_model_1.IRAM[0] [7], _40570_, clk);
  dff _88383_ (\oc8051_golden_model_1.B [0], _43194_, clk);
  dff _88384_ (\oc8051_golden_model_1.B [1], _43195_, clk);
  dff _88385_ (\oc8051_golden_model_1.B [2], _43196_, clk);
  dff _88386_ (\oc8051_golden_model_1.B [3], _43198_, clk);
  dff _88387_ (\oc8051_golden_model_1.B [4], _43199_, clk);
  dff _88388_ (\oc8051_golden_model_1.B [5], _43200_, clk);
  dff _88389_ (\oc8051_golden_model_1.B [6], _43201_, clk);
  dff _88390_ (\oc8051_golden_model_1.B [7], _40515_, clk);
  dff _88391_ (\oc8051_golden_model_1.ACC [0], _43203_, clk);
  dff _88392_ (\oc8051_golden_model_1.ACC [1], _43204_, clk);
  dff _88393_ (\oc8051_golden_model_1.ACC [2], _43205_, clk);
  dff _88394_ (\oc8051_golden_model_1.ACC [3], _43206_, clk);
  dff _88395_ (\oc8051_golden_model_1.ACC [4], _43207_, clk);
  dff _88396_ (\oc8051_golden_model_1.ACC [5], _43208_, clk);
  dff _88397_ (\oc8051_golden_model_1.ACC [6], _43209_, clk);
  dff _88398_ (\oc8051_golden_model_1.ACC [7], _40516_, clk);
  dff _88399_ (\oc8051_golden_model_1.SBUF [0], _43210_, clk);
  dff _88400_ (\oc8051_golden_model_1.SBUF [1], _43211_, clk);
  dff _88401_ (\oc8051_golden_model_1.SBUF [2], _43212_, clk);
  dff _88402_ (\oc8051_golden_model_1.SBUF [3], _43213_, clk);
  dff _88403_ (\oc8051_golden_model_1.SBUF [4], _43214_, clk);
  dff _88404_ (\oc8051_golden_model_1.SBUF [5], _43217_, clk);
  dff _88405_ (\oc8051_golden_model_1.SBUF [6], _43218_, clk);
  dff _88406_ (\oc8051_golden_model_1.SBUF [7], _40517_, clk);
  dff _88407_ (\oc8051_golden_model_1.SCON [0], _43219_, clk);
  dff _88408_ (\oc8051_golden_model_1.SCON [1], _43222_, clk);
  dff _88409_ (\oc8051_golden_model_1.SCON [2], _43223_, clk);
  dff _88410_ (\oc8051_golden_model_1.SCON [3], _43224_, clk);
  dff _88411_ (\oc8051_golden_model_1.SCON [4], _43225_, clk);
  dff _88412_ (\oc8051_golden_model_1.SCON [5], _43226_, clk);
  dff _88413_ (\oc8051_golden_model_1.SCON [6], _43227_, clk);
  dff _88414_ (\oc8051_golden_model_1.SCON [7], _40518_, clk);
  dff _88415_ (\oc8051_golden_model_1.PCON [0], _43228_, clk);
  dff _88416_ (\oc8051_golden_model_1.PCON [1], _43229_, clk);
  dff _88417_ (\oc8051_golden_model_1.PCON [2], _43230_, clk);
  dff _88418_ (\oc8051_golden_model_1.PCON [3], _43231_, clk);
  dff _88419_ (\oc8051_golden_model_1.PCON [4], _43232_, clk);
  dff _88420_ (\oc8051_golden_model_1.PCON [5], _43233_, clk);
  dff _88421_ (\oc8051_golden_model_1.PCON [6], _43234_, clk);
  dff _88422_ (\oc8051_golden_model_1.PCON [7], _40520_, clk);
  dff _88423_ (\oc8051_golden_model_1.TCON [0], _43237_, clk);
  dff _88424_ (\oc8051_golden_model_1.TCON [1], _43238_, clk);
  dff _88425_ (\oc8051_golden_model_1.TCON [2], _43239_, clk);
  dff _88426_ (\oc8051_golden_model_1.TCON [3], _43242_, clk);
  dff _88427_ (\oc8051_golden_model_1.TCON [4], _43243_, clk);
  dff _88428_ (\oc8051_golden_model_1.TCON [5], _43244_, clk);
  dff _88429_ (\oc8051_golden_model_1.TCON [6], _43245_, clk);
  dff _88430_ (\oc8051_golden_model_1.TCON [7], _40521_, clk);
  dff _88431_ (\oc8051_golden_model_1.TL0 [0], _43246_, clk);
  dff _88432_ (\oc8051_golden_model_1.TL0 [1], _43247_, clk);
  dff _88433_ (\oc8051_golden_model_1.TL0 [2], _43248_, clk);
  dff _88434_ (\oc8051_golden_model_1.TL0 [3], _43249_, clk);
  dff _88435_ (\oc8051_golden_model_1.TL0 [4], _43250_, clk);
  dff _88436_ (\oc8051_golden_model_1.TL0 [5], _43251_, clk);
  dff _88437_ (\oc8051_golden_model_1.TL0 [6], _43252_, clk);
  dff _88438_ (\oc8051_golden_model_1.TL0 [7], _40522_, clk);
  dff _88439_ (\oc8051_golden_model_1.TL1 [0], _43255_, clk);
  dff _88440_ (\oc8051_golden_model_1.TL1 [1], _43256_, clk);
  dff _88441_ (\oc8051_golden_model_1.TL1 [2], _43257_, clk);
  dff _88442_ (\oc8051_golden_model_1.TL1 [3], _43258_, clk);
  dff _88443_ (\oc8051_golden_model_1.TL1 [4], _43259_, clk);
  dff _88444_ (\oc8051_golden_model_1.TL1 [5], _43262_, clk);
  dff _88445_ (\oc8051_golden_model_1.TL1 [6], _43263_, clk);
  dff _88446_ (\oc8051_golden_model_1.TL1 [7], _40523_, clk);
  dff _88447_ (\oc8051_golden_model_1.TH0 [0], _43264_, clk);
  dff _88448_ (\oc8051_golden_model_1.TH0 [1], _43265_, clk);
  dff _88449_ (\oc8051_golden_model_1.TH0 [2], _43266_, clk);
  dff _88450_ (\oc8051_golden_model_1.TH0 [3], _43267_, clk);
  dff _88451_ (\oc8051_golden_model_1.TH0 [4], _43268_, clk);
  dff _88452_ (\oc8051_golden_model_1.TH0 [5], _43269_, clk);
  dff _88453_ (\oc8051_golden_model_1.TH0 [6], _43270_, clk);
  dff _88454_ (\oc8051_golden_model_1.TH0 [7], _40524_, clk);
  dff _88455_ (\oc8051_golden_model_1.TH1 [0], _43273_, clk);
  dff _88456_ (\oc8051_golden_model_1.TH1 [1], _43274_, clk);
  dff _88457_ (\oc8051_golden_model_1.TH1 [2], _43275_, clk);
  dff _88458_ (\oc8051_golden_model_1.TH1 [3], _43276_, clk);
  dff _88459_ (\oc8051_golden_model_1.TH1 [4], _43277_, clk);
  dff _88460_ (\oc8051_golden_model_1.TH1 [5], _43278_, clk);
  dff _88461_ (\oc8051_golden_model_1.TH1 [6], _43279_, clk);
  dff _88462_ (\oc8051_golden_model_1.TH1 [7], _40526_, clk);
  dff _88463_ (\oc8051_golden_model_1.TMOD [0], _43282_, clk);
  dff _88464_ (\oc8051_golden_model_1.TMOD [1], _43283_, clk);
  dff _88465_ (\oc8051_golden_model_1.TMOD [2], _43284_, clk);
  dff _88466_ (\oc8051_golden_model_1.TMOD [3], _43285_, clk);
  dff _88467_ (\oc8051_golden_model_1.TMOD [4], _43286_, clk);
  dff _88468_ (\oc8051_golden_model_1.TMOD [5], _43287_, clk);
  dff _88469_ (\oc8051_golden_model_1.TMOD [6], _43288_, clk);
  dff _88470_ (\oc8051_golden_model_1.TMOD [7], _40527_, clk);
  dff _88471_ (\oc8051_golden_model_1.IE [0], _43291_, clk);
  dff _88472_ (\oc8051_golden_model_1.IE [1], _43292_, clk);
  dff _88473_ (\oc8051_golden_model_1.IE [2], _43293_, clk);
  dff _88474_ (\oc8051_golden_model_1.IE [3], _43294_, clk);
  dff _88475_ (\oc8051_golden_model_1.IE [4], _43295_, clk);
  dff _88476_ (\oc8051_golden_model_1.IE [5], _43296_, clk);
  dff _88477_ (\oc8051_golden_model_1.IE [6], _43297_, clk);
  dff _88478_ (\oc8051_golden_model_1.IE [7], _40528_, clk);
  dff _88479_ (\oc8051_golden_model_1.IP [0], _43300_, clk);
  dff _88480_ (\oc8051_golden_model_1.IP [1], _43301_, clk);
  dff _88481_ (\oc8051_golden_model_1.IP [2], _43302_, clk);
  dff _88482_ (\oc8051_golden_model_1.IP [3], _43303_, clk);
  dff _88483_ (\oc8051_golden_model_1.IP [4], _43304_, clk);
  dff _88484_ (\oc8051_golden_model_1.IP [5], _43305_, clk);
  dff _88485_ (\oc8051_golden_model_1.IP [6], _43306_, clk);
  dff _88486_ (\oc8051_golden_model_1.IP [7], _40529_, clk);
  dff _88487_ (\oc8051_golden_model_1.DPL [0], _43307_, clk);
  dff _88488_ (\oc8051_golden_model_1.DPL [1], _43310_, clk);
  dff _88489_ (\oc8051_golden_model_1.DPL [2], _43311_, clk);
  dff _88490_ (\oc8051_golden_model_1.DPL [3], _43312_, clk);
  dff _88491_ (\oc8051_golden_model_1.DPL [4], _43313_, clk);
  dff _88492_ (\oc8051_golden_model_1.DPL [5], _43314_, clk);
  dff _88493_ (\oc8051_golden_model_1.DPL [6], _43315_, clk);
  dff _88494_ (\oc8051_golden_model_1.DPL [7], _40530_, clk);
  dff _88495_ (\oc8051_golden_model_1.DPH [0], _43318_, clk);
  dff _88496_ (\oc8051_golden_model_1.DPH [1], _43319_, clk);
  dff _88497_ (\oc8051_golden_model_1.DPH [2], _43320_, clk);
  dff _88498_ (\oc8051_golden_model_1.DPH [3], _43321_, clk);
  dff _88499_ (\oc8051_golden_model_1.DPH [4], _43322_, clk);
  dff _88500_ (\oc8051_golden_model_1.DPH [5], _43323_, clk);
  dff _88501_ (\oc8051_golden_model_1.DPH [6], _43324_, clk);
  dff _88502_ (\oc8051_golden_model_1.DPH [7], _40532_, clk);
  dff _88503_ (\oc8051_golden_model_1.PC [0], _43327_, clk);
  dff _88504_ (\oc8051_golden_model_1.PC [1], _43328_, clk);
  dff _88505_ (\oc8051_golden_model_1.PC [2], _43329_, clk);
  dff _88506_ (\oc8051_golden_model_1.PC [3], _43330_, clk);
  dff _88507_ (\oc8051_golden_model_1.PC [4], _43331_, clk);
  dff _88508_ (\oc8051_golden_model_1.PC [5], _43334_, clk);
  dff _88509_ (\oc8051_golden_model_1.PC [6], _43335_, clk);
  dff _88510_ (\oc8051_golden_model_1.PC [7], _43336_, clk);
  dff _88511_ (\oc8051_golden_model_1.PC [8], _43337_, clk);
  dff _88512_ (\oc8051_golden_model_1.PC [9], _43338_, clk);
  dff _88513_ (\oc8051_golden_model_1.PC [10], _43339_, clk);
  dff _88514_ (\oc8051_golden_model_1.PC [11], _43340_, clk);
  dff _88515_ (\oc8051_golden_model_1.PC [12], _43341_, clk);
  dff _88516_ (\oc8051_golden_model_1.PC [13], _43342_, clk);
  dff _88517_ (\oc8051_golden_model_1.PC [14], _43343_, clk);
  dff _88518_ (\oc8051_golden_model_1.PC [15], _40533_, clk);
  dff _88519_ (\oc8051_golden_model_1.P2 [0], _43345_, clk);
  dff _88520_ (\oc8051_golden_model_1.P2 [1], _43346_, clk);
  dff _88521_ (\oc8051_golden_model_1.P2 [2], _43347_, clk);
  dff _88522_ (\oc8051_golden_model_1.P2 [3], _43350_, clk);
  dff _88523_ (\oc8051_golden_model_1.P2 [4], _43351_, clk);
  dff _88524_ (\oc8051_golden_model_1.P2 [5], _43352_, clk);
  dff _88525_ (\oc8051_golden_model_1.P2 [6], _43353_, clk);
  dff _88526_ (\oc8051_golden_model_1.P2 [7], _40534_, clk);
  dff _88527_ (\oc8051_golden_model_1.P3 [0], _43355_, clk);
  dff _88528_ (\oc8051_golden_model_1.P3 [1], _43356_, clk);
  dff _88529_ (\oc8051_golden_model_1.P3 [2], _43357_, clk);
  dff _88530_ (\oc8051_golden_model_1.P3 [3], _43358_, clk);
  dff _88531_ (\oc8051_golden_model_1.P3 [4], _43359_, clk);
  dff _88532_ (\oc8051_golden_model_1.P3 [5], _43360_, clk);
  dff _88533_ (\oc8051_golden_model_1.P3 [6], _43361_, clk);
  dff _88534_ (\oc8051_golden_model_1.P3 [7], _40535_, clk);
  dff _88535_ (\oc8051_golden_model_1.P0 [0], _43363_, clk);
  dff _88536_ (\oc8051_golden_model_1.P0 [1], _43364_, clk);
  dff _88537_ (\oc8051_golden_model_1.P0 [2], _43365_, clk);
  dff _88538_ (\oc8051_golden_model_1.P0 [3], _43366_, clk);
  dff _88539_ (\oc8051_golden_model_1.P0 [4], _43367_, clk);
  dff _88540_ (\oc8051_golden_model_1.P0 [5], _43369_, clk);
  dff _88541_ (\oc8051_golden_model_1.P0 [6], _43370_, clk);
  dff _88542_ (\oc8051_golden_model_1.P0 [7], _40536_, clk);
  dff _88543_ (\oc8051_golden_model_1.P1 [0], _43371_, clk);
  dff _88544_ (\oc8051_golden_model_1.P1 [1], _43373_, clk);
  dff _88545_ (\oc8051_golden_model_1.P1 [2], _43374_, clk);
  dff _88546_ (\oc8051_golden_model_1.P1 [3], _43375_, clk);
  dff _88547_ (\oc8051_golden_model_1.P1 [4], _43376_, clk);
  dff _88548_ (\oc8051_golden_model_1.P1 [5], _43377_, clk);
  dff _88549_ (\oc8051_golden_model_1.P1 [6], _43378_, clk);
  dff _88550_ (\oc8051_golden_model_1.P1 [7], _40538_, clk);
  dff _88551_ (\oc8051_golden_model_1.SP [0], _43379_, clk);
  dff _88552_ (\oc8051_golden_model_1.SP [1], _43380_, clk);
  dff _88553_ (\oc8051_golden_model_1.SP [2], _43381_, clk);
  dff _88554_ (\oc8051_golden_model_1.SP [3], _43382_, clk);
  dff _88555_ (\oc8051_golden_model_1.SP [4], _43383_, clk);
  dff _88556_ (\oc8051_golden_model_1.SP [5], _43384_, clk);
  dff _88557_ (\oc8051_golden_model_1.SP [6], _43385_, clk);
  dff _88558_ (\oc8051_golden_model_1.SP [7], _40539_, clk);
  dff _88559_ (\oc8051_golden_model_1.PSW [0], _43388_, clk);
  dff _88560_ (\oc8051_golden_model_1.PSW [1], _43389_, clk);
  dff _88561_ (\oc8051_golden_model_1.PSW [2], _43390_, clk);
  dff _88562_ (\oc8051_golden_model_1.PSW [3], _43393_, clk);
  dff _88563_ (\oc8051_golden_model_1.PSW [4], _43394_, clk);
  dff _88564_ (\oc8051_golden_model_1.PSW [5], _43395_, clk);
  dff _88565_ (\oc8051_golden_model_1.PSW [6], _43396_, clk);
  dff _88566_ (\oc8051_golden_model_1.PSW [7], _40540_, clk);
  dff _88567_ (\oc8051_golden_model_1.P0INREG [0], _43397_, clk);
  dff _88568_ (\oc8051_golden_model_1.P0INREG [1], _43398_, clk);
  dff _88569_ (\oc8051_golden_model_1.P0INREG [2], _43399_, clk);
  dff _88570_ (\oc8051_golden_model_1.P0INREG [3], _43400_, clk);
  dff _88571_ (\oc8051_golden_model_1.P0INREG [4], _43401_, clk);
  dff _88572_ (\oc8051_golden_model_1.P0INREG [5], _43402_, clk);
  dff _88573_ (\oc8051_golden_model_1.P0INREG [6], _43403_, clk);
  dff _88574_ (\oc8051_golden_model_1.P0INREG [7], _40541_, clk);
  dff _88575_ (\oc8051_golden_model_1.P1INREG [0], _43406_, clk);
  dff _88576_ (\oc8051_golden_model_1.P1INREG [1], _43407_, clk);
  dff _88577_ (\oc8051_golden_model_1.P1INREG [2], _43408_, clk);
  dff _88578_ (\oc8051_golden_model_1.P1INREG [3], _43409_, clk);
  dff _88579_ (\oc8051_golden_model_1.P1INREG [4], _43410_, clk);
  dff _88580_ (\oc8051_golden_model_1.P1INREG [5], _43413_, clk);
  dff _88581_ (\oc8051_golden_model_1.P1INREG [6], _43414_, clk);
  dff _88582_ (\oc8051_golden_model_1.P1INREG [7], _40542_, clk);
  dff _88583_ (\oc8051_golden_model_1.P2INREG [0], _43415_, clk);
  dff _88584_ (\oc8051_golden_model_1.P2INREG [1], _43416_, clk);
  dff _88585_ (\oc8051_golden_model_1.P2INREG [2], _43417_, clk);
  dff _88586_ (\oc8051_golden_model_1.P2INREG [3], _43418_, clk);
  dff _88587_ (\oc8051_golden_model_1.P2INREG [4], _43419_, clk);
  dff _88588_ (\oc8051_golden_model_1.P2INREG [5], _43420_, clk);
  dff _88589_ (\oc8051_golden_model_1.P2INREG [6], _43421_, clk);
  dff _88590_ (\oc8051_golden_model_1.P2INREG [7], _40544_, clk);
  dff _88591_ (\oc8051_golden_model_1.P3INREG [0], _43424_, clk);
  dff _88592_ (\oc8051_golden_model_1.P3INREG [1], _43425_, clk);
  dff _88593_ (\oc8051_golden_model_1.P3INREG [2], _43426_, clk);
  dff _88594_ (\oc8051_golden_model_1.P3INREG [3], _43427_, clk);
  dff _88595_ (\oc8051_golden_model_1.P3INREG [4], _43428_, clk);
  dff _88596_ (\oc8051_golden_model_1.P3INREG [5], _43429_, clk);
  dff _88597_ (\oc8051_golden_model_1.P3INREG [6], _43430_, clk);
  dff _88598_ (\oc8051_golden_model_1.P3INREG [7], _40545_, clk);
  dff _88599_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _03015_, clk);
  dff _88600_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _03026_, clk);
  dff _88601_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _03047_, clk);
  dff _88602_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03069_, clk);
  dff _88603_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03090_, clk);
  dff _88604_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00894_, clk);
  dff _88605_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03101_, clk);
  dff _88606_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00863_, clk);
  dff _88607_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03112_, clk);
  dff _88608_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03123_, clk);
  dff _88609_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03134_, clk);
  dff _88610_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03145_, clk);
  dff _88611_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03156_, clk);
  dff _88612_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03167_, clk);
  dff _88613_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03178_, clk);
  dff _88614_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00915_, clk);
  dff _88615_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02465_, clk);
  dff _88616_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22440_, clk);
  dff _88617_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02660_, clk);
  dff _88618_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02854_, clk);
  dff _88619_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03058_, clk);
  dff _88620_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03269_, clk);
  dff _88621_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03470_, clk);
  dff _88622_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03671_, clk);
  dff _88623_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03872_, clk);
  dff _88624_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04073_, clk);
  dff _88625_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04174_, clk);
  dff _88626_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04275_, clk);
  dff _88627_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04376_, clk);
  dff _88628_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04477_, clk);
  dff _88629_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04578_, clk);
  dff _88630_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04679_, clk);
  dff _88631_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04780_, clk);
  dff _88632_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24614_, clk);
  dff _88633_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38774_, clk);
  dff _88634_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38775_, clk);
  dff _88635_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38776_, clk);
  dff _88636_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38777_, clk);
  dff _88637_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38778_, clk);
  dff _88638_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38779_, clk);
  dff _88639_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38780_, clk);
  dff _88640_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38759_, clk);
  dff _88641_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38781_, clk);
  dff _88642_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38783_, clk);
  dff _88643_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38784_, clk);
  dff _88644_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38785_, clk);
  dff _88645_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38786_, clk);
  dff _88646_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38787_, clk);
  dff _88647_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38789_, clk);
  dff _88648_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38761_, clk);
  dff _88649_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38790_, clk);
  dff _88650_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38791_, clk);
  dff _88651_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38792_, clk);
  dff _88652_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38793_, clk);
  dff _88653_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38795_, clk);
  dff _88654_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38796_, clk);
  dff _88655_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38797_, clk);
  dff _88656_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38762_, clk);
  dff _88657_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _30491_, clk);
  dff _88658_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06012_, clk);
  dff _88659_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _30494_, clk);
  dff _88660_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _06015_, clk);
  dff _88661_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _30496_, clk);
  dff _88662_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _30498_, clk);
  dff _88663_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06018_, clk);
  dff _88664_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _30500_, clk);
  dff _88665_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _30502_, clk);
  dff _88666_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06021_, clk);
  dff _88667_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _30504_, clk);
  dff _88668_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _06024_, clk);
  dff _88669_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _30506_, clk);
  dff _88670_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _30508_, clk);
  dff _88671_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _30510_, clk);
  dff _88672_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _06027_, clk);
  dff _88673_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _30512_, clk);
  dff _88674_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _06030_, clk);
  dff _88675_ (\oc8051_top_1.oc8051_decoder1.wr , _06033_, clk);
  dff _88676_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _06092_, clk);
  dff _88677_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _06094_, clk);
  dff _88678_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _05997_, clk);
  dff _88679_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _06097_, clk);
  dff _88680_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _06100_, clk);
  dff _88681_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _06000_, clk);
  dff _88682_ (\oc8051_top_1.oc8051_decoder1.state [0], _06103_, clk);
  dff _88683_ (\oc8051_top_1.oc8051_decoder1.state [1], _06003_, clk);
  dff _88684_ (\oc8051_top_1.oc8051_decoder1.op [0], _06106_, clk);
  dff _88685_ (\oc8051_top_1.oc8051_decoder1.op [1], _06109_, clk);
  dff _88686_ (\oc8051_top_1.oc8051_decoder1.op [2], _06112_, clk);
  dff _88687_ (\oc8051_top_1.oc8051_decoder1.op [3], _06115_, clk);
  dff _88688_ (\oc8051_top_1.oc8051_decoder1.op [4], _06118_, clk);
  dff _88689_ (\oc8051_top_1.oc8051_decoder1.op [5], _06121_, clk);
  dff _88690_ (\oc8051_top_1.oc8051_decoder1.op [6], _06124_, clk);
  dff _88691_ (\oc8051_top_1.oc8051_decoder1.op [7], _06006_, clk);
  dff _88692_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _06009_, clk);
  dff _88693_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39563_, clk);
  dff _88694_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _38933_, clk);
  dff _88695_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _38934_, clk);
  dff _88696_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _38935_, clk);
  dff _88697_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _38937_, clk);
  dff _88698_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _38938_, clk);
  dff _88699_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _38939_, clk);
  dff _88700_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _38940_, clk);
  dff _88701_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _38941_, clk);
  dff _88702_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _38942_, clk);
  dff _88703_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _38943_, clk);
  dff _88704_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _38944_, clk);
  dff _88705_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _38945_, clk);
  dff _88706_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _38946_, clk);
  dff _88707_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _38948_, clk);
  dff _88708_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _38949_, clk);
  dff _88709_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _38821_, clk);
  dff _88710_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _38953_, clk);
  dff _88711_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _38954_, clk);
  dff _88712_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _38955_, clk);
  dff _88713_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _38956_, clk);
  dff _88714_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _38957_, clk);
  dff _88715_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _38958_, clk);
  dff _88716_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _38959_, clk);
  dff _88717_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _38960_, clk);
  dff _88718_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _38962_, clk);
  dff _88719_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _38963_, clk);
  dff _88720_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _38964_, clk);
  dff _88721_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _38965_, clk);
  dff _88722_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _38966_, clk);
  dff _88723_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _38967_, clk);
  dff _88724_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _38968_, clk);
  dff _88725_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38823_, clk);
  dff _88726_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39145_, clk);
  dff _88727_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39146_, clk);
  dff _88728_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39147_, clk);
  dff _88729_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39148_, clk);
  dff _88730_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39149_, clk);
  dff _88731_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39150_, clk);
  dff _88732_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39151_, clk);
  dff _88733_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39152_, clk);
  dff _88734_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39153_, clk);
  dff _88735_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39154_, clk);
  dff _88736_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39155_, clk);
  dff _88737_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39156_, clk);
  dff _88738_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39157_, clk);
  dff _88739_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39158_, clk);
  dff _88740_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39159_, clk);
  dff _88741_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39160_, clk);
  dff _88742_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39162_, clk);
  dff _88743_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39163_, clk);
  dff _88744_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39164_, clk);
  dff _88745_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39165_, clk);
  dff _88746_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39166_, clk);
  dff _88747_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39167_, clk);
  dff _88748_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39168_, clk);
  dff _88749_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39169_, clk);
  dff _88750_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39170_, clk);
  dff _88751_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39171_, clk);
  dff _88752_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39173_, clk);
  dff _88753_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39174_, clk);
  dff _88754_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39175_, clk);
  dff _88755_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39176_, clk);
  dff _88756_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39177_, clk);
  dff _88757_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _38886_, clk);
  dff _88758_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _38859_, clk);
  dff _88759_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _88760_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39178_, clk);
  dff _88761_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39179_, clk);
  dff _88762_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39180_, clk);
  dff _88763_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39181_, clk);
  dff _88764_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _38861_, clk);
  dff _88765_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39183_, clk);
  dff _88766_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39184_, clk);
  dff _88767_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39185_, clk);
  dff _88768_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39186_, clk);
  dff _88769_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39187_, clk);
  dff _88770_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39189_, clk);
  dff _88771_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39190_, clk);
  dff _88772_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _38862_, clk);
  dff _88773_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39191_, clk);
  dff _88774_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39192_, clk);
  dff _88775_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39193_, clk);
  dff _88776_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39194_, clk);
  dff _88777_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39195_, clk);
  dff _88778_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39196_, clk);
  dff _88779_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39197_, clk);
  dff _88780_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _38864_, clk);
  dff _88781_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39199_, clk);
  dff _88782_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39200_, clk);
  dff _88783_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39201_, clk);
  dff _88784_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39202_, clk);
  dff _88785_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39203_, clk);
  dff _88786_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39204_, clk);
  dff _88787_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39205_, clk);
  dff _88788_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _38865_, clk);
  dff _88789_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38866_, clk);
  dff _88790_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38867_, clk);
  dff _88791_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39206_, clk);
  dff _88792_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39207_, clk);
  dff _88793_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39208_, clk);
  dff _88794_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39210_, clk);
  dff _88795_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39211_, clk);
  dff _88796_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39212_, clk);
  dff _88797_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39213_, clk);
  dff _88798_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38868_, clk);
  dff _88799_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39214_, clk);
  dff _88800_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39215_, clk);
  dff _88801_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39216_, clk);
  dff _88802_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39217_, clk);
  dff _88803_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39218_, clk);
  dff _88804_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39219_, clk);
  dff _88805_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39221_, clk);
  dff _88806_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39222_, clk);
  dff _88807_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39223_, clk);
  dff _88808_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39224_, clk);
  dff _88809_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39225_, clk);
  dff _88810_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39226_, clk);
  dff _88811_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39227_, clk);
  dff _88812_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39228_, clk);
  dff _88813_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39229_, clk);
  dff _88814_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _38870_, clk);
  dff _88815_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39230_, clk);
  dff _88816_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39232_, clk);
  dff _88817_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39233_, clk);
  dff _88818_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39234_, clk);
  dff _88819_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39235_, clk);
  dff _88820_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39236_, clk);
  dff _88821_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39237_, clk);
  dff _88822_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39238_, clk);
  dff _88823_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39239_, clk);
  dff _88824_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39240_, clk);
  dff _88825_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39241_, clk);
  dff _88826_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39243_, clk);
  dff _88827_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39244_, clk);
  dff _88828_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39245_, clk);
  dff _88829_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39246_, clk);
  dff _88830_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _38871_, clk);
  dff _88831_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _38872_, clk);
  dff _88832_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38875_, clk);
  dff _88833_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _38873_, clk);
  dff _88834_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39247_, clk);
  dff _88835_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39248_, clk);
  dff _88836_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39249_, clk);
  dff _88837_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39250_, clk);
  dff _88838_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39251_, clk);
  dff _88839_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39252_, clk);
  dff _88840_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39254_, clk);
  dff _88841_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _38876_, clk);
  dff _88842_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39255_, clk);
  dff _88843_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39256_, clk);
  dff _88844_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _38877_, clk);
  dff _88845_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39257_, clk);
  dff _88846_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39258_, clk);
  dff _88847_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39259_, clk);
  dff _88848_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39260_, clk);
  dff _88849_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39261_, clk);
  dff _88850_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39262_, clk);
  dff _88851_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39263_, clk);
  dff _88852_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _38878_, clk);
  dff _88853_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39265_, clk);
  dff _88854_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39266_, clk);
  dff _88855_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39267_, clk);
  dff _88856_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39268_, clk);
  dff _88857_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39269_, clk);
  dff _88858_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39270_, clk);
  dff _88859_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39271_, clk);
  dff _88860_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _38879_, clk);
  dff _88861_ (\oc8051_top_1.oc8051_memory_interface1.reti , _38880_, clk);
  dff _88862_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39272_, clk);
  dff _88863_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39273_, clk);
  dff _88864_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39274_, clk);
  dff _88865_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39275_, clk);
  dff _88866_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39276_, clk);
  dff _88867_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39277_, clk);
  dff _88868_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39278_, clk);
  dff _88869_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _38882_, clk);
  dff _88870_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _38883_, clk);
  dff _88871_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _38884_, clk);
  dff _88872_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39279_, clk);
  dff _88873_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39280_, clk);
  dff _88874_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39281_, clk);
  dff _88875_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _38885_, clk);
  dff _88876_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39282_, clk);
  dff _88877_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39283_, clk);
  dff _88878_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39284_, clk);
  dff _88879_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39286_, clk);
  dff _88880_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39287_, clk);
  dff _88881_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39288_, clk);
  dff _88882_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39289_, clk);
  dff _88883_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39290_, clk);
  dff _88884_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39291_, clk);
  dff _88885_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39292_, clk);
  dff _88886_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39293_, clk);
  dff _88887_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39294_, clk);
  dff _88888_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39295_, clk);
  dff _88889_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39297_, clk);
  dff _88890_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39298_, clk);
  dff _88891_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39299_, clk);
  dff _88892_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39300_, clk);
  dff _88893_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39301_, clk);
  dff _88894_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39302_, clk);
  dff _88895_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39303_, clk);
  dff _88896_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39304_, clk);
  dff _88897_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39305_, clk);
  dff _88898_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39306_, clk);
  dff _88899_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39308_, clk);
  dff _88900_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39309_, clk);
  dff _88901_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39310_, clk);
  dff _88902_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39311_, clk);
  dff _88903_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39312_, clk);
  dff _88904_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39313_, clk);
  dff _88905_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39314_, clk);
  dff _88906_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39315_, clk);
  dff _88907_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _38887_, clk);
  dff _88908_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39316_, clk);
  dff _88909_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39317_, clk);
  dff _88910_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39319_, clk);
  dff _88911_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39320_, clk);
  dff _88912_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39321_, clk);
  dff _88913_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39322_, clk);
  dff _88914_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39323_, clk);
  dff _88915_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _38889_, clk);
  dff _88916_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _38890_, clk);
  dff _88917_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _38891_, clk);
  dff _88918_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39324_, clk);
  dff _88919_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39325_, clk);
  dff _88920_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39326_, clk);
  dff _88921_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39327_, clk);
  dff _88922_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39328_, clk);
  dff _88923_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39330_, clk);
  dff _88924_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39331_, clk);
  dff _88925_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39332_, clk);
  dff _88926_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39333_, clk);
  dff _88927_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39334_, clk);
  dff _88928_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39335_, clk);
  dff _88929_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39336_, clk);
  dff _88930_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39337_, clk);
  dff _88931_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39338_, clk);
  dff _88932_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39339_, clk);
  dff _88933_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _38892_, clk);
  dff _88934_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _38893_, clk);
  dff _88935_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _38894_, clk);
  dff _88936_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _38895_, clk);
  dff _88937_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39341_, clk);
  dff _88938_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39342_, clk);
  dff _88939_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39343_, clk);
  dff _88940_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39344_, clk);
  dff _88941_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39345_, clk);
  dff _88942_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39346_, clk);
  dff _88943_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39347_, clk);
  dff _88944_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39348_, clk);
  dff _88945_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39349_, clk);
  dff _88946_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39350_, clk);
  dff _88947_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39352_, clk);
  dff _88948_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39353_, clk);
  dff _88949_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39354_, clk);
  dff _88950_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39355_, clk);
  dff _88951_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39356_, clk);
  dff _88952_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _38896_, clk);
  dff _88953_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _38897_, clk);
  dff _88954_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _39709_, clk);
  dff _88955_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _39728_, clk);
  dff _88956_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _39729_, clk);
  dff _88957_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _39730_, clk);
  dff _88958_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _39731_, clk);
  dff _88959_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _39732_, clk);
  dff _88960_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _39733_, clk);
  dff _88961_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _39734_, clk);
  dff _88962_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _39710_, clk);
  dff _88963_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _39711_, clk);
  dff _88964_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _39735_, clk);
  dff _88965_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _39736_, clk);
  dff _88966_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _39712_, clk);
  dff _88967_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _43774_, clk);
  dff _88968_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _43778_, clk);
  dff _88969_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _43782_, clk);
  dff _88970_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _43785_, clk);
  dff _88971_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _43788_, clk);
  dff _88972_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _43792_, clk);
  dff _88973_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _43796_, clk);
  dff _88974_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _42826_, clk);
  dff _88975_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _43745_, clk);
  dff _88976_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _43749_, clk);
  dff _88977_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _43753_, clk);
  dff _88978_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _43757_, clk);
  dff _88979_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _43761_, clk);
  dff _88980_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _43765_, clk);
  dff _88981_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _43767_, clk);
  dff _88982_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _43769_, clk);
  dff _88983_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _43713_, clk);
  dff _88984_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _43717_, clk);
  dff _88985_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _43721_, clk);
  dff _88986_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _43725_, clk);
  dff _88987_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _43729_, clk);
  dff _88988_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _43733_, clk);
  dff _88989_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _43737_, clk);
  dff _88990_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _43740_, clk);
  dff _88991_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _43082_, clk);
  dff _88992_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _43088_, clk);
  dff _88993_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _43094_, clk);
  dff _88994_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _43100_, clk);
  dff _88995_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _43106_, clk);
  dff _88996_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _43112_, clk);
  dff _88997_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _43118_, clk);
  dff _88998_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _43121_, clk);
  dff _88999_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _43129_, clk);
  dff _89000_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _43133_, clk);
  dff _89001_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _43137_, clk);
  dff _89002_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _43141_, clk);
  dff _89003_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _43145_, clk);
  dff _89004_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _43149_, clk);
  dff _89005_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _43153_, clk);
  dff _89006_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _43156_, clk);
  dff _89007_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _43164_, clk);
  dff _89008_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _43168_, clk);
  dff _89009_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _43172_, clk);
  dff _89010_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _43176_, clk);
  dff _89011_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _43180_, clk);
  dff _89012_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _43184_, clk);
  dff _89013_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _43188_, clk);
  dff _89014_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _43191_, clk);
  dff _89015_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _43387_, clk);
  dff _89016_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _43405_, clk);
  dff _89017_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _43423_, clk);
  dff _89018_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _43434_, clk);
  dff _89019_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _43438_, clk);
  dff _89020_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _43442_, clk);
  dff _89021_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _43446_, clk);
  dff _89022_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _43449_, clk);
  dff _89023_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _43216_, clk);
  dff _89024_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _43236_, clk);
  dff _89025_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _43254_, clk);
  dff _89026_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _43272_, clk);
  dff _89027_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _43290_, clk);
  dff _89028_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _43309_, clk);
  dff _89029_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _43326_, clk);
  dff _89030_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _43344_, clk);
  dff _89031_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _43584_, clk);
  dff _89032_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _43588_, clk);
  dff _89033_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _43592_, clk);
  dff _89034_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _43596_, clk);
  dff _89035_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _43600_, clk);
  dff _89036_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _43604_, clk);
  dff _89037_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _43608_, clk);
  dff _89038_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _43611_, clk);
  dff _89039_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _43552_, clk);
  dff _89040_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _43556_, clk);
  dff _89041_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _43560_, clk);
  dff _89042_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _43564_, clk);
  dff _89043_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _43568_, clk);
  dff _89044_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _43572_, clk);
  dff _89045_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _43576_, clk);
  dff _89046_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _43579_, clk);
  dff _89047_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _43517_, clk);
  dff _89048_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _43521_, clk);
  dff _89049_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _43525_, clk);
  dff _89050_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _43529_, clk);
  dff _89051_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _43533_, clk);
  dff _89052_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _43537_, clk);
  dff _89053_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _43541_, clk);
  dff _89054_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _43544_, clk);
  dff _89055_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _43485_, clk);
  dff _89056_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _43489_, clk);
  dff _89057_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _43493_, clk);
  dff _89058_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _43497_, clk);
  dff _89059_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _43501_, clk);
  dff _89060_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _43505_, clk);
  dff _89061_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _43509_, clk);
  dff _89062_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _43512_, clk);
  dff _89063_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _43454_, clk);
  dff _89064_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _43458_, clk);
  dff _89065_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _43462_, clk);
  dff _89066_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _43465_, clk);
  dff _89067_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _43469_, clk);
  dff _89068_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _43473_, clk);
  dff _89069_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _43477_, clk);
  dff _89070_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _43480_, clk);
  dff _89071_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _43616_, clk);
  dff _89072_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _43620_, clk);
  dff _89073_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _43624_, clk);
  dff _89074_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _43628_, clk);
  dff _89075_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _43632_, clk);
  dff _89076_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _43636_, clk);
  dff _89077_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _43640_, clk);
  dff _89078_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _43643_, clk);
  dff _89079_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _43681_, clk);
  dff _89080_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _43685_, clk);
  dff _89081_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _43689_, clk);
  dff _89082_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _43693_, clk);
  dff _89083_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _43697_, clk);
  dff _89084_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _43701_, clk);
  dff _89085_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _43705_, clk);
  dff _89086_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _43708_, clk);
  dff _89087_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _43648_, clk);
  dff _89088_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _43652_, clk);
  dff _89089_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _43656_, clk);
  dff _89090_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _43660_, clk);
  dff _89091_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _43664_, clk);
  dff _89092_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _43668_, clk);
  dff _89093_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _43672_, clk);
  dff _89094_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _43675_, clk);
  dff _89095_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _01407_, clk);
  dff _89096_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _01409_, clk);
  dff _89097_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _01411_, clk);
  dff _89098_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _01413_, clk);
  dff _89099_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _01415_, clk);
  dff _89100_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _01416_, clk);
  dff _89101_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _01418_, clk);
  dff _89102_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _42815_, clk);
  dff _89103_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _89104_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _89105_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _89106_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _89107_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _89108_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _89109_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _89110_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _89111_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _89112_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _89113_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _89114_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _89115_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _89116_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _89117_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _89118_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _89119_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _89120_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _89121_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _89122_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _89123_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _89124_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _89125_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _89126_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _89127_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _89128_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _89129_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _89130_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _89131_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _89132_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _89133_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _89134_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _89135_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _89136_ (\oc8051_top_1.oc8051_sfr1.bit_out , _39594_, clk);
  dff _89137_ (\oc8051_top_1.oc8051_sfr1.wait_data , _39595_, clk);
  dff _89138_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39659_, clk);
  dff _89139_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39660_, clk);
  dff _89140_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39661_, clk);
  dff _89141_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39662_, clk);
  dff _89142_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39663_, clk);
  dff _89143_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39664_, clk);
  dff _89144_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39665_, clk);
  dff _89145_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39596_, clk);
  dff _89146_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39597_, clk);
  dff _89147_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _24171_, clk);
  dff _89148_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _24183_, clk);
  dff _89149_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _24195_, clk);
  dff _89150_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _24207_, clk);
  dff _89151_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _24219_, clk);
  dff _89152_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _24230_, clk);
  dff _89153_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _24242_, clk);
  dff _89154_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _22320_, clk);
  dff _89155_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08932_, clk);
  dff _89156_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08943_, clk);
  dff _89157_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08954_, clk);
  dff _89158_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08965_, clk);
  dff _89159_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08976_, clk);
  dff _89160_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08987_, clk);
  dff _89161_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08998_, clk);
  dff _89162_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06696_, clk);
  dff _89163_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13599_, clk);
  dff _89164_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13608_, clk);
  dff _89165_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13617_, clk);
  dff _89166_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13627_, clk);
  dff _89167_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13636_, clk);
  dff _89168_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13646_, clk);
  dff _89169_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13656_, clk);
  dff _89170_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12702_, clk);
  dff _89171_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13665_, clk);
  dff _89172_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13675_, clk);
  dff _89173_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13684_, clk);
  dff _89174_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13694_, clk);
  dff _89175_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13704_, clk);
  dff _89176_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13713_, clk);
  dff _89177_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13722_, clk);
  dff _89178_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12723_, clk);
  dff _89179_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0, clk);
  dff _89180_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0, clk);
  dff _89181_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _89182_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _41755_, clk);
  dff _89183_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _42678_, clk);
  dff _89184_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _42680_, clk);
  dff _89185_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42682_, clk);
  dff _89186_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _42684_, clk);
  dff _89187_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _42686_, clk);
  dff _89188_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _42688_, clk);
  dff _89189_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42690_, clk);
  dff _89190_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _41754_, clk);
  dff _89191_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _42692_, clk);
  dff _89192_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _41752_, clk);
  dff _89193_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _41750_, clk);
  dff _89194_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _42694_, clk);
  dff _89195_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _42696_, clk);
  dff _89196_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _41748_, clk);
  dff _89197_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _42698_, clk);
  dff _89198_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _42700_, clk);
  dff _89199_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _41746_, clk);
  dff _89200_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _42702_, clk);
  dff _89201_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _41744_, clk);
  dff _89202_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _42704_, clk);
  dff _89203_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _41743_, clk);
  dff _89204_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _41711_, clk);
  dff _89205_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _41709_, clk);
  dff _89206_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _41707_, clk);
  dff _89207_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _41705_, clk);
  dff _89208_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _42706_, clk);
  dff _89209_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _42708_, clk);
  dff _89210_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _42709_, clk);
  dff _89211_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _41702_, clk);
  dff _89212_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _42711_, clk);
  dff _89213_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _42713_, clk);
  dff _89214_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _42715_, clk);
  dff _89215_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _42717_, clk);
  dff _89216_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _42719_, clk);
  dff _89217_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _42721_, clk);
  dff _89218_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _42723_, clk);
  dff _89219_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _41701_, clk);
  dff _89220_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _42725_, clk);
  dff _89221_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _42727_, clk);
  dff _89222_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _42729_, clk);
  dff _89223_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _42731_, clk);
  dff _89224_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _42733_, clk);
  dff _89225_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _42735_, clk);
  dff _89226_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _42737_, clk);
  dff _89227_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _41698_, clk);
  dff _89228_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _41155_, clk);
  dff _89229_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _41157_, clk);
  dff _89230_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _41158_, clk);
  dff _89231_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _41160_, clk);
  dff _89232_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _41162_, clk);
  dff _89233_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _41164_, clk);
  dff _89234_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _41165_, clk);
  dff _89235_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35499_, clk);
  dff _89236_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _41167_, clk);
  dff _89237_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _41169_, clk);
  dff _89238_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _41171_, clk);
  dff _89239_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _41172_, clk);
  dff _89240_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _41174_, clk);
  dff _89241_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _41176_, clk);
  dff _89242_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _41178_, clk);
  dff _89243_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35522_, clk);
  dff _89244_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _41179_, clk);
  dff _89245_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _41181_, clk);
  dff _89246_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _41183_, clk);
  dff _89247_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _41185_, clk);
  dff _89248_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _41186_, clk);
  dff _89249_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _41188_, clk);
  dff _89250_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _41190_, clk);
  dff _89251_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35545_, clk);
  dff _89252_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _41192_, clk);
  dff _89253_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _41193_, clk);
  dff _89254_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _41195_, clk);
  dff _89255_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _41197_, clk);
  dff _89256_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _41198_, clk);
  dff _89257_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _41200_, clk);
  dff _89258_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _41202_, clk);
  dff _89259_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35568_, clk);
  dff _89260_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _21487_, clk);
  dff _89261_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _21499_, clk);
  dff _89262_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _21511_, clk);
  dff _89263_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _21523_, clk);
  dff _89264_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _21535_, clk);
  dff _89265_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _21547_, clk);
  dff _89266_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _16559_, clk);
  dff _89267_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09542_, clk);
  dff _89268_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10690_, clk);
  dff _89269_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10701_, clk);
  dff _89270_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10712_, clk);
  dff _89271_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10723_, clk);
  dff _89272_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10734_, clk);
  dff _89273_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10745_, clk);
  dff _89274_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10756_, clk);
  dff _89275_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09563_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0988 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0988 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0988 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0988 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0988 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0988 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0988 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0989 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0990 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0991 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0992 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0993 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0995 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0996 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1011 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1011 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1011 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1011 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1011 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1011 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1011 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1018 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1019 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.n1027 [0]);
  buf(\oc8051_golden_model_1.n1027 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1027 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1027 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1027 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1027 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1043 , \oc8051_golden_model_1.n1044 [0]);
  buf(\oc8051_golden_model_1.n1044 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1044 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1044 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1044 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1044 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1044 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1044 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1137 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1137 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1137 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1137 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1139 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1139 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1141 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1141 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1142 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1142 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1143 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1144 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1144 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1145 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1145 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1146 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1194 , \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n1239 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1240 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1240 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1240 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1240 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1240 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1240 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1240 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1241 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1241 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1241 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1241 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1241 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1241 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1241 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1241 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1242 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1242 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1242 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1242 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1242 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1242 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1242 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1242 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1243 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1244 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1244 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1244 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1247 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1247 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1247 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1247 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1247 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1247 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1247 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1248 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1248 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1248 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1248 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1248 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1248 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1248 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1249 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1251 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1252 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1253 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1255 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1256 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1264 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1264 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1280 , \oc8051_golden_model_1.n1281 [0]);
  buf(\oc8051_golden_model_1.n1281 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1281 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1281 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1281 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1281 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1281 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1281 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1323 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1323 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1323 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1323 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1323 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1323 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1323 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1323 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1323 [8], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1323 [9], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1323 [10], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1323 [11], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1323 [12], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1323 [13], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1323 [14], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1323 [15], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1325 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1325 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1325 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1325 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1325 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1325 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1325 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1328 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1329 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1330 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1331 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1332 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1340 , \oc8051_golden_model_1.n1341 [0]);
  buf(\oc8051_golden_model_1.n1341 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1341 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1341 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1341 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1341 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1341 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1343 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1347 [8], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1349 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1349 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1349 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1349 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1350 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1354 [4], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1356 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1356 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1356 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1356 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1356 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1356 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1356 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1356 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1356 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1364 , \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1365 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1365 [2], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1365 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1365 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1365 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1365 [6], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1365 [7], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.n1382 [2]);
  buf(\oc8051_golden_model_1.n1366 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.n1382 [6]);
  buf(\oc8051_golden_model_1.n1366 [6], \oc8051_golden_model_1.n1382 [7]);
  buf(\oc8051_golden_model_1.n1381 , \oc8051_golden_model_1.n1382 [0]);
  buf(\oc8051_golden_model_1.n1382 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1382 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1382 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1382 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1404 [8], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1405 , \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1410 [4], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1411 , \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1419 , \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1420 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1420 [2], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1420 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1420 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1420 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1420 [6], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1420 [7], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1421 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1421 [1], \oc8051_golden_model_1.n1437 [2]);
  buf(\oc8051_golden_model_1.n1421 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1421 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1421 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1421 [5], \oc8051_golden_model_1.n1437 [6]);
  buf(\oc8051_golden_model_1.n1421 [6], \oc8051_golden_model_1.n1437 [7]);
  buf(\oc8051_golden_model_1.n1436 , \oc8051_golden_model_1.n1437 [0]);
  buf(\oc8051_golden_model_1.n1437 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1437 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1437 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1437 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1439 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1439 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1439 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1439 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1439 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1439 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1439 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1439 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1439 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1441 [8], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1442 , \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1443 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1443 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1443 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1443 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1444 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1444 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1444 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1444 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1446 [4], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1447 , \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1448 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n1448 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n1448 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n1448 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n1448 [4], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n1448 [5], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n1448 [6], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n1448 [7], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1448 [8], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n1455 , \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1456 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1456 [2], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1456 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1456 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1456 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1456 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1456 [7], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1457 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.n1473 [2]);
  buf(\oc8051_golden_model_1.n1457 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1457 [6], \oc8051_golden_model_1.n1473 [7]);
  buf(\oc8051_golden_model_1.n1472 , \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [0], \oc8051_golden_model_1.n1487 [0]);
  buf(\oc8051_golden_model_1.n1473 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1473 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1473 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1473 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1473 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1476 [8], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1477 , \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1484 , \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1485 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1485 [2], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1485 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1485 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1485 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1485 [6], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1485 [7], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1486 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1486 [1], \oc8051_golden_model_1.n1487 [2]);
  buf(\oc8051_golden_model_1.n1486 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1486 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1486 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1486 [5], \oc8051_golden_model_1.n1487 [6]);
  buf(\oc8051_golden_model_1.n1486 [6], \oc8051_golden_model_1.n1487 [7]);
  buf(\oc8051_golden_model_1.n1487 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1487 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1487 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1487 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1489 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1489 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1489 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1489 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1489 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1489 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1489 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1489 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1489 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1491 [8], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1493 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1495 [4], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1496 , \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1497 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1497 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1497 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1497 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1497 [4], \oc8051_golden_model_1.n2751 );
  buf(\oc8051_golden_model_1.n1497 [5], \oc8051_golden_model_1.n2750 );
  buf(\oc8051_golden_model_1.n1497 [6], \oc8051_golden_model_1.n2749 );
  buf(\oc8051_golden_model_1.n1497 [7], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1497 [8], \oc8051_golden_model_1.n2748 );
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1521 , \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1522 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1524 [4], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1526 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1527 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1527 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1527 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1527 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1527 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1527 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1527 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1528 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1528 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1530 [8], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1531 , \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1538 , \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1539 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1539 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1539 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1539 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1539 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1539 [6], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1539 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1540 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1540 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1540 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1540 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1540 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1540 [5], \oc8051_golden_model_1.n1541 [6]);
  buf(\oc8051_golden_model_1.n1540 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1541 [0], \oc8051_golden_model_1.n1544 [0]);
  buf(\oc8051_golden_model_1.n1541 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1541 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1541 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1541 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1541 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1541 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1543 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1543 [1], \oc8051_golden_model_1.n1544 [2]);
  buf(\oc8051_golden_model_1.n1543 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1543 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1543 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1543 [5], \oc8051_golden_model_1.n1544 [6]);
  buf(\oc8051_golden_model_1.n1543 [6], \oc8051_golden_model_1.n1544 [7]);
  buf(\oc8051_golden_model_1.n1544 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1544 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1544 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1547 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1547 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1548 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1548 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1548 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1549 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1549 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1549 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1549 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1549 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1549 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1549 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1549 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1550 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1550 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1550 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1550 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1550 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1550 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1550 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1550 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1551 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1552 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1553 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1555 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1556 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1557 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1559 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1566 , \oc8051_golden_model_1.n1567 [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1568 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1571 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1571 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1573 [8], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1575 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1575 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1575 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1577 [4], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1585 , \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1586 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1586 [2], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1586 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1586 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1586 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1586 [6], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1586 [7], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1587 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.n1603 [2]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.n1603 [6]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.n1603 [7]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1603 [0]);
  buf(\oc8051_golden_model_1.n1603 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1603 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1603 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1603 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [8], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1608 , \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1610 [4], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1611 , \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1618 , \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1619 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1619 [2], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1619 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1619 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1619 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1619 [6], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1619 [7], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1620 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1620 [1], \oc8051_golden_model_1.n1636 [2]);
  buf(\oc8051_golden_model_1.n1620 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1620 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1620 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1620 [5], \oc8051_golden_model_1.n1636 [6]);
  buf(\oc8051_golden_model_1.n1620 [6], \oc8051_golden_model_1.n1636 [7]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1636 [0]);
  buf(\oc8051_golden_model_1.n1636 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1636 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1636 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1636 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [8], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1641 , \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1643 [4], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1644 , \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1651 , \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1652 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1652 [2], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1652 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1652 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1652 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1652 [6], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1652 [7], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1653 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1653 [1], \oc8051_golden_model_1.n1669 [2]);
  buf(\oc8051_golden_model_1.n1653 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1653 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1653 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1653 [5], \oc8051_golden_model_1.n1669 [6]);
  buf(\oc8051_golden_model_1.n1653 [6], \oc8051_golden_model_1.n1669 [7]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1669 [0]);
  buf(\oc8051_golden_model_1.n1669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [8], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1674 , \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1676 [4], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1677 , \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1684 , \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1685 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1685 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1685 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1685 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1685 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1685 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1685 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1686 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1686 [1], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1686 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1686 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1686 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1686 [5], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1686 [6], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1701 , \oc8051_golden_model_1.n1702 [0]);
  buf(\oc8051_golden_model_1.n1702 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1702 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1702 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1702 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1727 [1], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1727 [2], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1727 [3], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1727 [4], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1727 [5], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1727 [6], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1727 [7], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1728 [0], \oc8051_golden_model_1.n1729 [1]);
  buf(\oc8051_golden_model_1.n1728 [1], \oc8051_golden_model_1.n1729 [2]);
  buf(\oc8051_golden_model_1.n1728 [2], \oc8051_golden_model_1.n1729 [3]);
  buf(\oc8051_golden_model_1.n1728 [3], \oc8051_golden_model_1.n1729 [4]);
  buf(\oc8051_golden_model_1.n1728 [4], \oc8051_golden_model_1.n1729 [5]);
  buf(\oc8051_golden_model_1.n1728 [5], \oc8051_golden_model_1.n1729 [6]);
  buf(\oc8051_golden_model_1.n1728 [6], \oc8051_golden_model_1.n1729 [7]);
  buf(\oc8051_golden_model_1.n1729 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1784 , \oc8051_golden_model_1.n1785 [0]);
  buf(\oc8051_golden_model_1.n1785 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1785 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1785 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1785 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1785 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1785 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1785 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1801 , \oc8051_golden_model_1.n1802 [0]);
  buf(\oc8051_golden_model_1.n1802 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1802 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1802 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1802 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1802 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1802 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1802 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1818 , \oc8051_golden_model_1.n1819 [0]);
  buf(\oc8051_golden_model_1.n1819 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1819 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1819 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1819 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1819 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1819 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1819 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1835 , \oc8051_golden_model_1.n1836 [0]);
  buf(\oc8051_golden_model_1.n1836 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1836 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1836 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1836 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1836 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1836 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1836 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1859 [1], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1859 [2], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1859 [3], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1859 [4], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1859 [5], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1859 [6], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1859 [7], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1860 [0], \oc8051_golden_model_1.n1861 [1]);
  buf(\oc8051_golden_model_1.n1860 [1], \oc8051_golden_model_1.n1861 [2]);
  buf(\oc8051_golden_model_1.n1860 [2], \oc8051_golden_model_1.n1861 [3]);
  buf(\oc8051_golden_model_1.n1860 [3], \oc8051_golden_model_1.n1861 [4]);
  buf(\oc8051_golden_model_1.n1860 [4], \oc8051_golden_model_1.n1861 [5]);
  buf(\oc8051_golden_model_1.n1860 [5], \oc8051_golden_model_1.n1861 [6]);
  buf(\oc8051_golden_model_1.n1860 [6], \oc8051_golden_model_1.n1861 [7]);
  buf(\oc8051_golden_model_1.n1861 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n1916 , \oc8051_golden_model_1.n1917 [0]);
  buf(\oc8051_golden_model_1.n1917 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1917 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1917 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1917 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1917 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1917 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1917 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1933 , \oc8051_golden_model_1.n1934 [0]);
  buf(\oc8051_golden_model_1.n1934 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1934 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1934 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1934 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1934 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1934 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1934 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1950 , \oc8051_golden_model_1.n1951 [0]);
  buf(\oc8051_golden_model_1.n1951 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1951 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1951 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1951 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1951 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1951 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1951 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1967 , \oc8051_golden_model_1.n1968 [0]);
  buf(\oc8051_golden_model_1.n1968 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1968 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1968 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1968 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1968 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1968 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1968 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2065 , \oc8051_golden_model_1.n2066 [0]);
  buf(\oc8051_golden_model_1.n2066 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2066 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2066 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2066 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2066 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2066 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2066 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2082 , \oc8051_golden_model_1.n2083 [0]);
  buf(\oc8051_golden_model_1.n2083 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2083 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2083 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2083 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2083 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2083 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2083 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2099 , \oc8051_golden_model_1.n2100 [0]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2100 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2116 , \oc8051_golden_model_1.n2117 [0]);
  buf(\oc8051_golden_model_1.n2117 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2117 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2117 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2117 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2117 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2117 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2117 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2121 , \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2122 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2122 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2122 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2122 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2122 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2122 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2122 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2123 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2123 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2123 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2123 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2123 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2123 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2123 [7], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2124 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2124 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2124 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2124 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2124 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2124 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2124 [6], \oc8051_golden_model_1.n2125 [7]);
  buf(\oc8051_golden_model_1.n2125 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2125 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2125 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2125 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2125 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2125 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2125 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2140 , \oc8051_golden_model_1.n2141 [0]);
  buf(\oc8051_golden_model_1.n2141 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2141 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2141 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2141 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2141 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2141 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2180 , \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2181 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2181 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2181 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2181 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2181 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2181 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2181 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2181 [7], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2182 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2182 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2182 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2182 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2182 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2182 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2182 [6], \oc8051_golden_model_1.n2183 [7]);
  buf(\oc8051_golden_model_1.n2183 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2183 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2183 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2183 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2183 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2183 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2183 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2190 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2190 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2190 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2190 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2191 , \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2192 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2192 [2], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2192 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2192 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2192 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2192 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2192 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2193 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2193 [1], \oc8051_golden_model_1.n2209 [2]);
  buf(\oc8051_golden_model_1.n2193 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2193 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2193 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2193 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2193 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2208 , \oc8051_golden_model_1.n2209 [0]);
  buf(\oc8051_golden_model_1.n2209 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2209 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2209 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2209 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2209 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2209 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2421 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2421 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2424 , \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2426 , \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2432 , \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2433 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2433 [2], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2433 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2433 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2433 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2433 [6], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2433 [7], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2434 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2434 [1], \oc8051_golden_model_1.n2450 [2]);
  buf(\oc8051_golden_model_1.n2434 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2434 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2434 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2434 [5], \oc8051_golden_model_1.n2450 [6]);
  buf(\oc8051_golden_model_1.n2434 [6], \oc8051_golden_model_1.n2450 [7]);
  buf(\oc8051_golden_model_1.n2449 , \oc8051_golden_model_1.n2450 [0]);
  buf(\oc8051_golden_model_1.n2450 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2450 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2450 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2450 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 , \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2456 , \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2462 , \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2463 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2463 [2], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2463 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2463 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2463 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2463 [6], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2463 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2464 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2464 [1], \oc8051_golden_model_1.n2480 [2]);
  buf(\oc8051_golden_model_1.n2464 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2464 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2464 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2464 [5], \oc8051_golden_model_1.n2480 [6]);
  buf(\oc8051_golden_model_1.n2464 [6], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2479 , \oc8051_golden_model_1.n2480 [0]);
  buf(\oc8051_golden_model_1.n2480 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2480 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2480 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2480 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 , \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2486 , \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2492 , \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2493 [2], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2493 [6], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2493 [7], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2494 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2494 [1], \oc8051_golden_model_1.n2510 [2]);
  buf(\oc8051_golden_model_1.n2494 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2494 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2494 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2494 [5], \oc8051_golden_model_1.n2510 [6]);
  buf(\oc8051_golden_model_1.n2494 [6], \oc8051_golden_model_1.n2510 [7]);
  buf(\oc8051_golden_model_1.n2509 , \oc8051_golden_model_1.n2510 [0]);
  buf(\oc8051_golden_model_1.n2510 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2510 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2510 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2510 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 , \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2516 , \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2523 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2523 [2], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2523 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2523 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2523 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2523 [6], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2523 [7], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2524 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2524 [1], \oc8051_golden_model_1.n2540 [2]);
  buf(\oc8051_golden_model_1.n2524 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2524 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2524 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2524 [5], \oc8051_golden_model_1.n2540 [6]);
  buf(\oc8051_golden_model_1.n2524 [6], \oc8051_golden_model_1.n2540 [7]);
  buf(\oc8051_golden_model_1.n2539 , \oc8051_golden_model_1.n2540 [0]);
  buf(\oc8051_golden_model_1.n2540 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2540 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2540 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2540 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2545 [7]);
  buf(\oc8051_golden_model_1.n2545 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2545 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2545 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2545 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2545 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2545 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2545 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2546 [7], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2547 [6], \oc8051_golden_model_1.n2548 [7]);
  buf(\oc8051_golden_model_1.n2548 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2548 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2548 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2552 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2552 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2552 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2552 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2552 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2552 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2552 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2552 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2552 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2552 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2558 , \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2559 [2], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2559 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2559 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.n2576 [2]);
  buf(\oc8051_golden_model_1.n2560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2560 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2575 , \oc8051_golden_model_1.n2576 [0]);
  buf(\oc8051_golden_model_1.n2576 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2576 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2576 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2576 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2576 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2576 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2579 , \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [7], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2581 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2581 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2581 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2581 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2581 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2581 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2581 [6], \oc8051_golden_model_1.n2582 [7]);
  buf(\oc8051_golden_model_1.n2582 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2582 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2582 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2582 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2582 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2582 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2582 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2614 , \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2615 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2615 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2615 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2615 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2615 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2615 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2615 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2615 [7], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2616 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2616 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2616 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2616 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2616 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2616 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2616 [6], \oc8051_golden_model_1.n2617 [7]);
  buf(\oc8051_golden_model_1.n2617 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2617 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2617 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2617 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2617 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2617 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2617 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2622 , \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2623 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2623 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2623 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2623 [7], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2624 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2624 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2624 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2624 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2624 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2624 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2624 [6], \oc8051_golden_model_1.n2625 [7]);
  buf(\oc8051_golden_model_1.n2625 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2625 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2625 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2625 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2625 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2625 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2625 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2630 , \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2631 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2631 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2631 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2631 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2631 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2631 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2631 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2631 [7], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2632 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2632 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2632 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2632 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2632 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2632 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2632 [6], \oc8051_golden_model_1.n2633 [7]);
  buf(\oc8051_golden_model_1.n2633 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2633 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2633 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2633 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2633 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2633 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2633 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2638 , \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2639 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2639 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2639 [7], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2640 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2640 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2640 [6], \oc8051_golden_model_1.n2641 [7]);
  buf(\oc8051_golden_model_1.n2641 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2641 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2641 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2641 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2641 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2641 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2641 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2646 , \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2647 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2647 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2647 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2647 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2647 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2647 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2647 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2647 [7], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2648 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2648 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2648 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2648 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2648 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2648 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2648 [6], \oc8051_golden_model_1.n2649 [7]);
  buf(\oc8051_golden_model_1.n2649 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2649 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2649 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2649 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2649 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2649 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2649 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2674 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2674 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2674 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2674 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2674 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2674 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2674 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2675 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2675 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2675 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2675 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2675 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2675 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2675 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2676 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2676 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2676 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2676 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2676 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2676 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2676 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2676 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2677 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2677 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2677 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2677 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2678 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2678 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2678 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2678 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2678 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2678 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2678 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2679 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2680 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2681 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2682 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2683 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2684 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2685 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2686 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2693 , \oc8051_golden_model_1.n2694 [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2715 [0], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2715 [1], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2715 [2], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2715 [3], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2715 [4], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2715 [5], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2715 [6], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2731 [1], \oc8051_golden_model_1.n2893 [1]);
  buf(\oc8051_golden_model_1.n2731 [2], \oc8051_golden_model_1.n2893 [2]);
  buf(\oc8051_golden_model_1.n2731 [3], \oc8051_golden_model_1.n2893 [3]);
  buf(\oc8051_golden_model_1.n2731 [4], \oc8051_golden_model_1.n2893 [4]);
  buf(\oc8051_golden_model_1.n2731 [5], \oc8051_golden_model_1.n2893 [5]);
  buf(\oc8051_golden_model_1.n2731 [6], \oc8051_golden_model_1.n2893 [6]);
  buf(\oc8051_golden_model_1.n2731 [7], \oc8051_golden_model_1.n2893 [7]);
  buf(\oc8051_golden_model_1.n2732 , \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2733 , \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2734 , \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2735 , \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2736 , \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2737 , \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2738 , \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2739 , \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2746 , \oc8051_golden_model_1.n2747 [0]);
  buf(\oc8051_golden_model_1.n2747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2747 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2747 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2747 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2762 , \oc8051_golden_model_1.n2763 [0]);
  buf(\oc8051_golden_model_1.n2763 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2763 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2763 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2763 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2763 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2763 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2763 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2795 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2795 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2795 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2795 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2795 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2795 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2795 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2795 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2796 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2796 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2796 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2796 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2796 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2796 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2796 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2797 [0], \oc8051_golden_model_1.n2893 [0]);
  buf(\oc8051_golden_model_1.n2797 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2797 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2797 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2797 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2797 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2797 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2797 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 , \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2818 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2818 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2818 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2818 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2818 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2818 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2818 [6], \oc8051_golden_model_1.n2834 [7]);
  buf(\oc8051_golden_model_1.n2833 , \oc8051_golden_model_1.n2834 [0]);
  buf(\oc8051_golden_model_1.n2834 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2834 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2834 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2834 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2834 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2834 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.n2848 );
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.n2847 );
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.n2846 );
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.n2845 );
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2838 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2839 [0], \oc8051_golden_model_1.n2840 [4]);
  buf(\oc8051_golden_model_1.n2839 [1], \oc8051_golden_model_1.n2840 [5]);
  buf(\oc8051_golden_model_1.n2839 [2], \oc8051_golden_model_1.n2840 [6]);
  buf(\oc8051_golden_model_1.n2839 [3], \oc8051_golden_model_1.n2840 [7]);
  buf(\oc8051_golden_model_1.n2840 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2840 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2840 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2840 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2841 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2842 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2843 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2844 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2855 , \oc8051_golden_model_1.n2856 [0]);
  buf(\oc8051_golden_model_1.n2856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2874 , \oc8051_golden_model_1.n2875 [0]);
  buf(\oc8051_golden_model_1.n2875 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2875 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2875 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2875 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2875 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2875 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2875 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2891 , \oc8051_golden_model_1.n2892 [0]);
  buf(\oc8051_golden_model_1.n2892 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2892 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2892 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2892 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2892 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2892 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2892 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(ie_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(ie_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(ie_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(ie_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(ie_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(ie_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(ie_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(ie_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
