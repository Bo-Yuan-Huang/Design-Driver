
module oc8051_gm_top(clk, rst, word_in, xram_data_in, RD_IRAM_0_ABSTR_ADDR, RD_IRAM_1_ABSTR_ADDR, RD_ROM_1_ABSTR_ADDR, RD_ROM_2_ABSTR_ADDR, ACC_abstr, P2_abstr, P0_abstr, P1_abstr, P3_abstr, SP_abstr, PC_abstr, B_abstr, DPL_abstr, PSW_abstr, DPH_abstr, XRAM_DATA_OUT_abstr, XRAM_ADDR_abstr, WR_COND_ABSTR_IRAM_0, WR_ADDR_ABSTR_IRAM_0, WR_DATA_ABSTR_IRAM_0, WR_COND_ABSTR_IRAM_1, WR_ADDR_ABSTR_IRAM_1, WR_DATA_ABSTR_IRAM_1, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_xram_addr, property_invalid_xram_data_out);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire [7:0] _00006_;
  wire [7:0] _00007_;
  wire _00008_;
  wire _00009_;
  wire [7:0] _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire [7:0] _12609_;
  wire [7:0] _12610_;
  wire _12611_;
  wire [7:0] _12612_;
  wire [7:0] _12613_;
  wire [7:0] _12614_;
  wire [7:0] _12615_;
  wire [7:0] _12616_;
  wire [7:0] _12617_;
  wire [7:0] _12618_;
  wire [7:0] _12619_;
  wire [7:0] _12620_;
  wire [7:0] _12621_;
  wire [7:0] _12622_;
  wire [15:0] _12623_;
  wire [7:0] _12624_;
  wire [7:0] _12625_;
  wire [7:0] _12626_;
  wire [7:0] _12627_;
  wire [7:0] _12628_;
  wire [7:0] _12629_;
  wire [7:0] _12630_;
  wire [7:0] _12631_;
  wire [7:0] _12632_;
  wire [7:0] _12633_;
  wire [15:0] _12634_;
  wire [7:0] _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire [7:0] _12662_;
  wire [7:0] _12663_;
  wire [7:0] _12664_;
  wire [7:0] _12665_;
  wire [7:0] _12666_;
  wire [7:0] _12667_;
  wire [7:0] _12668_;
  wire [7:0] _12669_;
  wire [7:0] _12670_;
  wire [7:0] _12671_;
  wire [7:0] _12672_;
  wire [7:0] _12673_;
  wire [7:0] _12674_;
  wire [7:0] _12675_;
  wire [7:0] _12676_;
  wire [7:0] _12677_;
  wire [2:0] _12678_;
  wire [2:0] _12679_;
  wire [1:0] _12680_;
  wire [7:0] _12681_;
  wire _12682_;
  wire [1:0] _12683_;
  wire [1:0] _12684_;
  wire [2:0] _12685_;
  wire [2:0] _12686_;
  wire [1:0] _12687_;
  wire [3:0] _12688_;
  wire [1:0] _12689_;
  wire _12690_;
  wire _12691_;
  wire [15:0] _12692_;
  wire [15:0] _12693_;
  wire _12694_;
  wire _12695_;
  wire [4:0] _12696_;
  wire [7:0] _12697_;
  wire [7:0] _12698_;
  wire [7:0] _12699_;
  wire _12700_;
  wire _12701_;
  wire [7:0] _12702_;
  wire [15:0] _12703_;
  wire [15:0] _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire [7:0] _12708_;
  wire [2:0] _12709_;
  wire [7:0] _12710_;
  wire [7:0] _12711_;
  wire _12712_;
  wire [7:0] _12713_;
  wire _12714_;
  wire _12715_;
  wire [3:0] _12716_;
  wire [31:0] _12717_;
  wire [31:0] _12718_;
  wire [7:0] _12719_;
  wire _12720_;
  wire _12721_;
  wire [15:0] _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire [15:0] _12726_;
  wire _12727_;
  wire _12728_;
  wire [7:0] _12729_;
  wire _12730_;
  wire [2:0] _12731_;
  wire _12732_;
  wire _12733_;
  wire [7:0] _12734_;
  wire _12735_;
  input [7:0] ACC_abstr;
  wire [7:0] ACC_gm;
  input [7:0] B_abstr;
  wire [7:0] B_gm;
  input [7:0] DPH_abstr;
  wire [7:0] DPH_gm;
  input [7:0] DPL_abstr;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IE_gm_next;
  wire [7:0] IP_gm;
  wire [7:0] IP_gm_next;
  input [7:0] P0_abstr;
  wire [7:0] P0_gm;
  input [7:0] P1_abstr;
  wire [7:0] P1_gm;
  input [7:0] P2_abstr;
  wire [7:0] P2_gm;
  input [7:0] P3_abstr;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PCON_gm_next;
  input [15:0] PC_abstr;
  input [7:0] PSW_abstr;
  wire [7:0] PSW_gm;
  input [7:0] RD_IRAM_0_ABSTR_ADDR;
  input [7:0] RD_IRAM_1_ABSTR_ADDR;
  input [15:0] RD_ROM_1_ABSTR_ADDR;
  input [15:0] RD_ROM_2_ABSTR_ADDR;
  wire [7:0] SBUF_gm;
  wire [7:0] SBUF_gm_next;
  wire [7:0] SCON_gm;
  wire [7:0] SCON_gm_next;
  input [7:0] SP_abstr;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TCON_gm_next;
  wire [7:0] TH0_gm;
  wire [7:0] TH0_gm_next;
  wire [7:0] TH1_gm;
  wire [7:0] TH1_gm_next;
  wire [7:0] TL0_gm;
  wire [7:0] TL0_gm_next;
  wire [7:0] TL1_gm;
  wire [7:0] TL1_gm_next;
  wire [7:0] TMOD_gm;
  wire [7:0] TMOD_gm_next;
  input [3:0] WR_ADDR_ABSTR_IRAM_0;
  input [3:0] WR_ADDR_ABSTR_IRAM_1;
  input WR_COND_ABSTR_IRAM_0;
  input WR_COND_ABSTR_IRAM_1;
  input [7:0] WR_DATA_ABSTR_IRAM_0;
  input [7:0] WR_DATA_ABSTR_IRAM_1;
  input [15:0] XRAM_ADDR_abstr;
  input [7:0] XRAM_DATA_OUT_abstr;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire eq_state_1;
  wire eq_state_2;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_1 ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_2 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_abstr ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.B_49 ;
  wire [7:0] \oc8051_golden_model_1.B_abstr ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPH_49 ;
  wire [7:0] \oc8051_golden_model_1.DPH_abstr ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.DPL_49 ;
  wire [7:0] \oc8051_golden_model_1.DPL_abstr ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IE_next ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IP_next ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0_49 ;
  wire [7:0] \oc8051_golden_model_1.P0_abstr ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1_49 ;
  wire [7:0] \oc8051_golden_model_1.P1_abstr ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2_49 ;
  wire [7:0] \oc8051_golden_model_1.P2_abstr ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3_49 ;
  wire [7:0] \oc8051_golden_model_1.P3_abstr ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [7:0] \oc8051_golden_model_1.PCON_next ;
  wire [15:0] \oc8051_golden_model_1.PC_abstr ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_abstr ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_1_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_2_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SBUF_next ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SCON_next ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.SP_49 ;
  wire [7:0] \oc8051_golden_model_1.SP_abstr ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TCON_next ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH0_next ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TH1_next ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL0_next ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TL1_next ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire [7:0] \oc8051_golden_model_1.TMOD_next ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_0_IRAM ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_1_IRAM ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 ;
  wire [3:0] \oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 ;
  wire \oc8051_golden_model_1.WR_COND_ABSTR_IRAM_0 ;
  wire \oc8051_golden_model_1.WR_COND_ABSTR_IRAM_1 ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_0_IRAM ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_1_IRAM ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_abstr ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_IN ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_abstr ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0004 ;
  wire [7:0] \oc8051_golden_model_1.n0006 ;
  wire [3:0] \oc8051_golden_model_1.n0010 ;
  wire [7:0] \oc8051_golden_model_1.n0085 ;
  wire [3:0] \oc8051_golden_model_1.n0086 ;
  wire [3:0] \oc8051_golden_model_1.n0088 ;
  wire [7:0] \oc8051_golden_model_1.n0090 ;
  wire [3:0] \oc8051_golden_model_1.n0091 ;
  wire [7:0] \oc8051_golden_model_1.n0093 ;
  wire [3:0] \oc8051_golden_model_1.n0094 ;
  wire [7:0] \oc8051_golden_model_1.n0096 ;
  wire [3:0] \oc8051_golden_model_1.n0097 ;
  wire [7:0] \oc8051_golden_model_1.n0099 ;
  wire [3:0] \oc8051_golden_model_1.n0100 ;
  wire [7:0] \oc8051_golden_model_1.n0102 ;
  wire [3:0] \oc8051_golden_model_1.n0103 ;
  wire [7:0] \oc8051_golden_model_1.n0105 ;
  wire [3:0] \oc8051_golden_model_1.n0106 ;
  wire [6:0] \oc8051_golden_model_1.n0170 ;
  wire \oc8051_golden_model_1.n0185 ;
  wire [7:0] \oc8051_golden_model_1.n0186 ;
  wire \oc8051_golden_model_1.n0236 ;
  wire [7:0] \oc8051_golden_model_1.n0237 ;
  wire [3:0] \oc8051_golden_model_1.n0277 ;
  wire [3:0] \oc8051_golden_model_1.n0278 ;
  wire [7:0] \oc8051_golden_model_1.n0279 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_i ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_i ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire \oc8051_top_1.wbd_ack_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_i ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  output property_invalid_xram_addr;
  output property_invalid_xram_data_out;
  wire property_valid_psw_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  wire [15:0] rd_rom_1_addr;
  wire [15:0] rd_rom_2_addr;
  input rst;
  wire this_op_cnst_r;
  wire wbd_ack_i;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_i;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  input [7:0] xram_data_in;
  wire [7:0] xram_data_in_model;
  wire [7:0] xram_data_in_reg;
  not (_05610_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_05611_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05610_);
  and (_05612_, _05611_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05613_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05610_);
  and (_05614_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05610_);
  nor (_05615_, _05614_, _05613_);
  and (_05616_, _05615_, _05612_);
  not (_05617_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_05618_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _05617_);
  not (_05619_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_05621_, _05619_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nor (_05622_, _05621_, _05618_);
  nand (_05623_, _05622_, _05616_);
  not (_12493_, rst);
  or (_05624_, _05616_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_05625_, _05624_, _12493_);
  and (_06348_, _05625_, _05623_);
  nor (_05626_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_05627_, _05626_);
  and (_05628_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_05629_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  nor (_05630_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_05631_, _05630_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05632_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_05633_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_05634_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_05635_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_05636_, _05635_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_05637_, _05636_, _05634_);
  nor (_05638_, _05637_, _05633_);
  nor (_05639_, _05638_, _05632_);
  and (_05640_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_05641_, _05640_, _05634_);
  and (_05642_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_05643_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05644_, _05643_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_05645_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_05646_, _05645_, _05642_);
  and (_05647_, _05646_, _05639_);
  not (_05648_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_05649_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05648_);
  or (_05650_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  not (_05651_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_05652_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _05651_);
  and (_05653_, _05652_, _05650_);
  or (_05654_, _05653_, _05649_);
  nand (_05655_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05648_);
  or (_05656_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_05657_, _05656_, _05654_);
  nand (_05658_, _05630_, _05634_);
  or (_05659_, _05658_, _05657_);
  or (_05660_, _05636_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_05661_, _05660_);
  and (_05662_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_05663_, _05640_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05664_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_05665_, _05664_, _05662_);
  and (_05666_, _05665_, _05659_);
  and (_05667_, _05666_, _05647_);
  not (_05668_, _05667_);
  or (_05669_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_05670_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or (_05671_, _05651_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_05672_, _05671_, _05670_);
  or (_05673_, _05672_, _05649_);
  or (_05674_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_05675_, _05674_, _05673_);
  or (_05676_, _05675_, _05669_);
  and (_05677_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_05678_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_05679_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_05680_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_05681_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _05680_);
  nor (_05682_, _05681_, _05679_);
  nor (_05683_, _05682_, _05678_);
  and (_05684_, _05683_, _05676_);
  nand (_05685_, _05684_, _05626_);
  not (_05686_, _05618_);
  or (_05687_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_05688_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _05651_);
  and (_05689_, _05688_, _05687_);
  or (_05690_, _05689_, _05649_);
  or (_05691_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_05692_, _05691_, _05690_);
  or (_05693_, _05692_, _05669_);
  nand (_05694_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not (_05695_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_05696_, _05681_, _05695_);
  and (_05697_, _05696_, _05694_);
  and (_05698_, _05697_, _05693_);
  or (_05699_, _05698_, _05686_);
  not (_05700_, _05621_);
  or (_05701_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_05702_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _05651_);
  and (_05703_, _05702_, _05701_);
  or (_05704_, _05703_, _05649_);
  or (_05705_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_05706_, _05705_, _05704_);
  or (_05707_, _05706_, _05669_);
  nand (_05708_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not (_05709_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_05710_, _05681_, _05709_);
  and (_05711_, _05710_, _05708_);
  and (_05712_, _05711_, _05707_);
  or (_05713_, _05712_, _05700_);
  and (_05714_, _05713_, _05699_);
  or (_05715_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_05716_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _05651_);
  and (_05717_, _05716_, _05715_);
  or (_05718_, _05717_, _05649_);
  or (_05719_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_05720_, _05719_, _05718_);
  or (_05721_, _05720_, _05669_);
  nand (_05722_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not (_05723_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_05724_, _05681_, _05723_);
  and (_05725_, _05724_, _05722_);
  nand (_05726_, _05725_, _05721_);
  or (_05727_, _05726_, _05617_);
  nand (_05728_, _05727_, _05622_);
  nand (_05729_, _05728_, _05714_);
  and (_05730_, _05729_, _05685_);
  and (_05731_, _05730_, _05668_);
  or (_05732_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  or (_05733_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _05651_);
  and (_05734_, _05733_, _05732_);
  or (_05735_, _05734_, _05649_);
  or (_05736_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_05737_, _05736_, _05735_);
  or (_05738_, _05737_, _05669_);
  and (_05739_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_05740_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05741_, _05681_, _05740_);
  nor (_05742_, _05741_, _05739_);
  and (_05743_, _05742_, _05738_);
  nand (_05744_, _05743_, _05626_);
  or (_05745_, _05657_, _05669_);
  nand (_05746_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_05747_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_05748_, _05681_, _05747_);
  and (_05749_, _05748_, _05746_);
  and (_05750_, _05749_, _05745_);
  or (_05751_, _05750_, _05686_);
  or (_05752_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_05753_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _05651_);
  and (_05754_, _05753_, _05752_);
  or (_05755_, _05754_, _05649_);
  or (_05756_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_05757_, _05756_, _05755_);
  or (_05758_, _05757_, _05669_);
  nand (_05759_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_05760_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_05761_, _05681_, _05760_);
  and (_05762_, _05761_, _05759_);
  and (_05763_, _05762_, _05758_);
  or (_05764_, _05763_, _05700_);
  and (_05765_, _05764_, _05751_);
  or (_05766_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_05767_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _05651_);
  and (_05768_, _05767_, _05766_);
  or (_05769_, _05768_, _05649_);
  or (_05770_, _05655_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_05771_, _05770_, _05769_);
  or (_05772_, _05771_, _05669_);
  nand (_05773_, _05677_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not (_05774_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_05775_, _05681_, _05774_);
  and (_05776_, _05775_, _05773_);
  nand (_05777_, _05776_, _05772_);
  or (_05778_, _05777_, _05617_);
  nand (_05779_, _05778_, _05622_);
  nand (_05780_, _05779_, _05765_);
  and (_05781_, _05780_, _05744_);
  not (_05782_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_05783_, _05637_, _05782_);
  nand (_05784_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_05785_, _05784_, _05783_);
  nand (_05786_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nand (_05787_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_05788_, _05787_, _05786_);
  and (_05789_, _05788_, _05785_);
  or (_05790_, _05706_, _05658_);
  nand (_05791_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nand (_05792_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_05793_, _05792_, _05791_);
  and (_05794_, _05793_, _05790_);
  and (_05795_, _05794_, _05789_);
  not (_05796_, _05795_);
  and (_05797_, _05796_, _05781_);
  and (_05798_, _05797_, _05731_);
  and (_05799_, _05668_, _05781_);
  not (_05800_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_05801_, _05637_, _05800_);
  and (_05802_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_05803_, _05802_, _05801_);
  and (_05804_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_05805_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_05806_, _05805_, _05804_);
  and (_05807_, _05806_, _05803_);
  or (_05808_, _05692_, _05658_);
  and (_05809_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_05810_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05811_, _05810_, _05809_);
  and (_05812_, _05811_, _05808_);
  and (_05813_, _05812_, _05807_);
  not (_05814_, _05813_);
  and (_05815_, _05814_, _05730_);
  nand (_05816_, _05815_, _05799_);
  and (_05817_, _05814_, _05781_);
  or (_05818_, _05817_, _05731_);
  and (_05819_, _05818_, _05816_);
  and (_05820_, _05819_, _05798_);
  not (_05821_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_05822_, _05637_, _05821_);
  and (_05823_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_05824_, _05823_, _05822_);
  and (_05825_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_05826_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_05827_, _05826_, _05825_);
  and (_05828_, _05827_, _05824_);
  or (_05829_, _05658_, _05737_);
  and (_05830_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_05831_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05832_, _05831_, _05830_);
  and (_05833_, _05832_, _05829_);
  and (_05834_, _05833_, _05828_);
  or (_05835_, _05834_, _05816_);
  not (_05836_, _05834_);
  and (_05837_, _05836_, _05781_);
  not (_05838_, _05837_);
  nand (_05839_, _05838_, _05816_);
  and (_05840_, _05839_, _05835_);
  nand (_05841_, _05840_, _05815_);
  or (_05842_, _05837_, _05815_);
  and (_05843_, _05842_, _05841_);
  nand (_05844_, _05843_, _05820_);
  not (_05845_, _05844_);
  not (_05846_, _05835_);
  and (_05847_, _05840_, _05815_);
  nand (_05848_, _05729_, _05685_);
  or (_05849_, _05834_, _05848_);
  nand (_05850_, _05780_, _05744_);
  and (_05851_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_05852_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_05853_, _05637_, _05852_);
  nor (_05854_, _05853_, _05851_);
  and (_05855_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_05856_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_05857_, _05856_, _05855_);
  and (_05858_, _05857_, _05854_);
  nor (_05859_, _05675_, _05658_);
  not (_05860_, _05859_);
  and (_05861_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_05862_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_05863_, _05862_, _05861_);
  and (_05864_, _05863_, _05860_);
  and (_05865_, _05864_, _05858_);
  or (_05866_, _05865_, _05850_);
  or (_05867_, _05866_, _05849_);
  nand (_05868_, _05866_, _05849_);
  and (_05869_, _05868_, _05867_);
  nand (_05870_, _05869_, _05847_);
  or (_05871_, _05869_, _05847_);
  and (_05872_, _05871_, _05870_);
  nand (_05873_, _05872_, _05846_);
  or (_05874_, _05872_, _05846_);
  and (_05875_, _05874_, _05873_);
  nand (_05876_, _05875_, _05845_);
  or (_05877_, _05875_, _05845_);
  nand (_05878_, _05877_, _05876_);
  not (_05879_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_05880_, _05637_, _05879_);
  nand (_05881_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_05882_, _05881_, _05880_);
  nand (_05883_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nand (_05884_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_05885_, _05884_, _05883_);
  and (_05886_, _05885_, _05882_);
  or (_05887_, _05720_, _05658_);
  nand (_05888_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand (_05889_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_05890_, _05889_, _05888_);
  and (_05891_, _05890_, _05887_);
  nand (_05892_, _05891_, _05886_);
  and (_05893_, _05892_, _05730_);
  nand (_05894_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand (_05895_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_05896_, _05895_, _05894_);
  not (_05897_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_05898_, _05637_, _05897_);
  nand (_05899_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_05900_, _05899_, _05898_);
  and (_05901_, _05900_, _05896_);
  or (_05902_, _05658_, _05757_);
  nand (_05903_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand (_05904_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_05905_, _05904_, _05903_);
  and (_05906_, _05905_, _05902_);
  nand (_05907_, _05906_, _05901_);
  and (_05908_, _05907_, _05781_);
  and (_05909_, _05908_, _05893_);
  not (_05910_, _05909_);
  and (_05911_, _05892_, _05781_);
  not (_05912_, _05911_);
  and (_05913_, _05907_, _05730_);
  and (_05914_, _05913_, _05912_);
  nand (_05915_, _05914_, _05797_);
  nand (_05916_, _05915_, _05910_);
  not (_05917_, _05798_);
  and (_05918_, _05796_, _05730_);
  or (_05919_, _05918_, _05799_);
  and (_05920_, _05919_, _05917_);
  and (_05921_, _05920_, _05916_);
  not (_05922_, _05820_);
  or (_05923_, _05819_, _05798_);
  and (_05924_, _05923_, _05922_);
  and (_05925_, _05924_, _05921_);
  or (_05926_, _05843_, _05820_);
  and (_05927_, _05926_, _05844_);
  nand (_05928_, _05927_, _05925_);
  not (_05929_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_05930_, _05637_, _05929_);
  and (_05931_, _05631_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_05932_, _05931_, _05930_);
  and (_05933_, _05661_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_05934_, _05644_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_05935_, _05934_, _05933_);
  and (_05936_, _05935_, _05932_);
  nor (_05937_, _05658_, _05771_);
  and (_05938_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_05939_, _05663_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_05940_, _05939_, _05938_);
  not (_05941_, _05940_);
  nor (_05942_, _05941_, _05937_);
  and (_05943_, _05942_, _05936_);
  not (_05944_, _05943_);
  and (_05945_, _05944_, _05730_);
  and (_05946_, _05945_, _05911_);
  or (_05947_, _05908_, _05893_);
  and (_05948_, _05947_, _05910_);
  and (_05949_, _05948_, _05946_);
  or (_05950_, _05914_, _05797_);
  and (_05951_, _05950_, _05915_);
  nand (_05952_, _05951_, _05949_);
  not (_05953_, _05952_);
  nand (_05954_, _05920_, _05916_);
  or (_05955_, _05920_, _05916_);
  and (_05956_, _05955_, _05954_);
  nand (_05957_, _05956_, _05953_);
  nand (_05958_, _05924_, _05921_);
  or (_05959_, _05924_, _05921_);
  nand (_05960_, _05959_, _05958_);
  or (_05961_, _05960_, _05957_);
  or (_05962_, _05927_, _05925_);
  nand (_05963_, _05962_, _05928_);
  or (_05964_, _05963_, _05961_);
  and (_05965_, _05964_, _05928_);
  or (_05966_, _05965_, _05878_);
  nand (_05967_, _05966_, _05876_);
  not (_05968_, _05865_);
  and (_05969_, _05968_, _05730_);
  and (_05970_, _05969_, _05838_);
  and (_05971_, _05873_, _05870_);
  not (_05972_, _05971_);
  nand (_05973_, _05972_, _05970_);
  or (_05974_, _05972_, _05970_);
  and (_05975_, _05974_, _05973_);
  nand (_05976_, _05975_, _05967_);
  and (_05977_, _05973_, _05867_);
  nand (_05978_, _05977_, _05976_);
  or (_05979_, _05978_, _05629_);
  nand (_05980_, _05978_, _05629_);
  and (_05981_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_05982_, _05975_, _05967_);
  and (_05983_, _05982_, _05976_);
  nand (_05984_, _05983_, _05981_);
  nand (_05985_, _05984_, _05980_);
  nand (_05986_, _05985_, _05979_);
  and (_05987_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_05988_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_05989_, _05988_, _05987_);
  not (_05990_, _05989_);
  nor (_05991_, _05990_, _05986_);
  and (_05992_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_05993_, _05965_, _05878_);
  and (_05994_, _05993_, _05966_);
  nand (_05995_, _05994_, _05992_);
  or (_05996_, _05994_, _05992_);
  nand (_05997_, _05996_, _05995_);
  and (_05998_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand (_05999_, _05963_, _05961_);
  and (_06000_, _05999_, _05964_);
  nand (_06001_, _06000_, _05998_);
  or (_06002_, _06000_, _05998_);
  nand (_06003_, _06002_, _06001_);
  and (_06004_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand (_06005_, _05960_, _05957_);
  and (_06006_, _06005_, _05961_);
  nand (_06007_, _06006_, _06004_);
  or (_06008_, _06006_, _06004_);
  nand (_06009_, _06008_, _06007_);
  and (_06010_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_06011_, _05956_, _05953_);
  and (_06012_, _06011_, _05957_);
  nand (_06013_, _06012_, _06010_);
  and (_06014_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_06015_, _05951_, _05949_);
  and (_06016_, _06015_, _05952_);
  nand (_06017_, _06016_, _06014_);
  and (_06018_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_06019_, _05948_, _05946_);
  or (_06020_, _05948_, _05946_);
  and (_06021_, _06020_, _06019_);
  and (_06022_, _06021_, _06018_);
  not (_06023_, _06022_);
  or (_06024_, _06016_, _06014_);
  nand (_06025_, _06024_, _06017_);
  or (_06026_, _06025_, _06023_);
  and (_06027_, _06026_, _06017_);
  or (_06028_, _06012_, _06010_);
  nand (_06029_, _06028_, _06013_);
  or (_06030_, _06029_, _06027_);
  and (_06031_, _06030_, _06013_);
  or (_06032_, _06031_, _06009_);
  and (_06033_, _06032_, _06007_);
  or (_06034_, _06033_, _06003_);
  and (_06035_, _06034_, _06001_);
  or (_06036_, _06035_, _05997_);
  nand (_06037_, _06036_, _05995_);
  and (_06038_, _05980_, _05979_);
  or (_06039_, _05983_, _05981_);
  and (_06040_, _06039_, _05984_);
  and (_06041_, _06040_, _06038_);
  and (_06042_, _05989_, _06041_);
  and (_06043_, _06042_, _06037_);
  or (_06044_, _06043_, _05991_);
  and (_06045_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_06046_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_06047_, _06046_, _06045_);
  and (_06048_, _06047_, _06044_);
  nand (_06049_, _06048_, _05628_);
  and (_06050_, _05627_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_06051_, _06050_, _06049_);
  or (_06052_, _06049_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_06053_, _06052_, _06051_);
  and (_06542_, _06053_, _12493_);
  nor (_06054_, _05616_, _05619_);
  and (_06055_, _05616_, _05619_);
  or (_06056_, _06055_, _06054_);
  and (_02732_, _06056_, _12493_);
  and (_06057_, _05944_, _05781_);
  and (_02918_, _06057_, _12493_);
  nor (_06058_, _05945_, _05911_);
  nor (_06059_, _06058_, _05946_);
  and (_03102_, _06059_, _12493_);
  nor (_06060_, _06021_, _06018_);
  nor (_06061_, _06060_, _06022_);
  and (_03276_, _06061_, _12493_);
  and (_06062_, _06025_, _06023_);
  not (_06063_, _06062_);
  and (_06064_, _06063_, _06026_);
  and (_03449_, _06064_, _12493_);
  and (_06065_, _06029_, _06027_);
  not (_06066_, _06065_);
  and (_06068_, _06066_, _06030_);
  and (_03619_, _06068_, _12493_);
  and (_06071_, _06031_, _06009_);
  not (_06073_, _06071_);
  and (_06075_, _06073_, _06032_);
  and (_03811_, _06075_, _12493_);
  and (_06077_, _06033_, _06003_);
  not (_06078_, _06077_);
  and (_06079_, _06078_, _06034_);
  and (_04009_, _06079_, _12493_);
  and (_06080_, _06035_, _05997_);
  not (_06081_, _06080_);
  and (_06082_, _06081_, _06036_);
  and (_04153_, _06082_, _12493_);
  and (_06083_, _06040_, _06037_);
  nor (_06084_, _06040_, _06037_);
  nor (_06085_, _06084_, _06083_);
  and (_04221_, _06085_, _12493_);
  not (_06086_, _06083_);
  and (_06087_, _06086_, _05984_);
  and (_06088_, _06087_, _06038_);
  nor (_06089_, _06087_, _06038_);
  or (_06090_, _06089_, _06088_);
  and (_04268_, _06090_, _12493_);
  nand (_06091_, _06083_, _06038_);
  and (_06092_, _06091_, _05986_);
  not (_06093_, _06092_);
  nand (_06094_, _06093_, _05987_);
  or (_06095_, _06093_, _05987_);
  and (_06096_, _06095_, _06094_);
  and (_04356_, _06096_, _12493_);
  not (_06097_, _05988_);
  and (_06098_, _06097_, _06094_);
  nor (_06099_, _06098_, _06044_);
  and (_04433_, _06099_, _12493_);
  nand (_06100_, _06045_, _06044_);
  or (_06101_, _06045_, _06044_);
  and (_06102_, _06101_, _06100_);
  and (_04509_, _06102_, _12493_);
  not (_06103_, _06046_);
  and (_06104_, _06103_, _06100_);
  nor (_06105_, _06104_, _06048_);
  and (_04610_, _06105_, _12493_);
  or (_06106_, _06048_, _05628_);
  and (_06107_, _06106_, _06049_);
  and (_04711_, _06107_, _12493_);
  and (_06108_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05610_);
  nor (_06109_, _06108_, _05611_);
  not (_06110_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_06111_, _05613_, _06110_);
  and (_06112_, _06111_, _06109_);
  and (_06113_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_06114_, _06113_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_06115_, _06113_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_06116_, _06115_, _06114_);
  and (_01016_, _06116_, _12493_);
  and (_01047_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _12493_);
  nor (_06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_06118_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_06119_, _06118_);
  nand (_06120_, _06117_, _05865_);
  and (_06121_, _06120_, _06119_);
  not (_06122_, _06121_);
  or (_06123_, _05777_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_06124_, _05763_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_06125_, _06124_, _06123_);
  or (_06126_, _06125_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_06127_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_06128_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_06129_, _05750_, _06128_);
  nand (_06130_, _05743_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_06131_, _06130_, _06129_);
  or (_06132_, _06131_, _06127_);
  and (_06133_, _06132_, _06126_);
  or (_06134_, _06133_, _06122_);
  and (_06135_, _06117_, _05834_);
  nor (_06137_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor (_06138_, _06137_, _06135_);
  and (_06139_, _05725_, _05721_);
  or (_06140_, _06139_, _06128_);
  and (_06141_, _06140_, _06127_);
  not (_06142_, _06141_);
  nand (_06143_, _05712_, _06128_);
  nand (_06144_, _05698_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_06145_, _06144_, _06143_);
  or (_06146_, _06145_, _06127_);
  and (_06147_, _06146_, _06142_);
  not (_06148_, _06147_);
  and (_06149_, _06148_, _06138_);
  not (_06150_, _06133_);
  or (_06151_, _06150_, _06121_);
  and (_06152_, _06151_, _06134_);
  nand (_06153_, _06152_, _06149_);
  and (_06154_, _06153_, _06134_);
  nor (_06155_, _06148_, _06138_);
  nor (_06156_, _06155_, _06149_);
  and (_06157_, _06156_, _06152_);
  nand (_06158_, _06117_, _05813_);
  nor (_06159_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_06160_, _06159_);
  and (_06161_, _06160_, _06158_);
  not (_06162_, _06161_);
  and (_06163_, _05777_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_06164_, _06163_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_06165_, _05763_, _06128_);
  nand (_06166_, _05750_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_06167_, _06166_, _06165_);
  or (_06168_, _06167_, _06127_);
  and (_06169_, _06168_, _06164_);
  or (_06170_, _06169_, _06162_);
  or (_06171_, _05726_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_06172_, _05712_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_06173_, _06172_, _06171_);
  and (_06174_, _06173_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_06175_, _06174_);
  nor (_06176_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_06177_, _06176_);
  nand (_06178_, _06117_, _05667_);
  and (_06179_, _06178_, _06177_);
  nand (_06180_, _06179_, _06175_);
  nand (_06181_, _06169_, _06162_);
  and (_06182_, _06170_, _06181_);
  not (_06183_, _06182_);
  or (_06184_, _06183_, _06180_);
  nand (_06185_, _06184_, _06170_);
  and (_06186_, _06125_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_06187_, _06186_);
  nand (_06188_, _06117_, _05795_);
  nor (_06189_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_06190_, _06189_);
  and (_06191_, _06190_, _06188_);
  nand (_06192_, _06191_, _06187_);
  or (_06193_, _06191_, _06187_);
  nand (_06194_, _06193_, _06192_);
  or (_06195_, _06140_, _06127_);
  nor (_06196_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_06197_, _06196_);
  not (_06198_, _06117_);
  or (_06199_, _06198_, _05907_);
  and (_06200_, _06199_, _06197_);
  nand (_06201_, _06200_, _06195_);
  and (_06202_, _06163_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_06203_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_06204_, _06203_);
  or (_06205_, _06198_, _05892_);
  nand (_06206_, _06205_, _06204_);
  and (_06207_, _06206_, _06202_);
  or (_06208_, _06200_, _06195_);
  nand (_06209_, _06208_, _06201_);
  or (_06210_, _06209_, _06207_);
  and (_06211_, _06210_, _06201_);
  or (_06212_, _06211_, _06194_);
  nand (_06213_, _06212_, _06192_);
  or (_06214_, _06179_, _06175_);
  and (_06215_, _06214_, _06180_);
  and (_06216_, _06182_, _06215_);
  and (_06217_, _06216_, _06213_);
  or (_06218_, _06217_, _06185_);
  nand (_06219_, _06218_, _06157_);
  nand (_06220_, _06219_, _06154_);
  and (_06221_, _05684_, _05743_);
  nor (_06222_, _06221_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_06223_, _06167_, _06131_);
  and (_06224_, _05698_, _06128_);
  and (_06225_, _05684_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_06226_, _06225_, _06224_);
  nor (_06227_, _06226_, _06145_);
  and (_06228_, _06227_, _06223_);
  nor (_06229_, _06228_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_06230_, _06229_, _06222_);
  nor (_06231_, _06173_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_06232_, _06226_, _06127_);
  nor (_06233_, _06232_, _06231_);
  not (_06234_, _06233_);
  and (_06235_, _06234_, _06230_);
  and (_06236_, _06235_, _06220_);
  nor (_06237_, _06236_, _06122_);
  not (_06238_, _06236_);
  and (_06239_, _06218_, _06156_);
  nor (_06240_, _06239_, _06149_);
  and (_06241_, _06240_, _06152_);
  nor (_06242_, _06240_, _06152_);
  nor (_06243_, _06242_, _06241_);
  nor (_06244_, _06243_, _06238_);
  nor (_06245_, _06244_, _06237_);
  and (_06246_, _06245_, _06233_);
  nor (_06247_, _06245_, _06233_);
  nor (_06248_, _06218_, _06156_);
  nor (_06249_, _06248_, _06239_);
  nor (_06250_, _06249_, _06238_);
  nor (_06251_, _06236_, _06138_);
  nor (_06252_, _06251_, _06250_);
  and (_06253_, _06252_, _06150_);
  nor (_06254_, _06253_, _06247_);
  nor (_06255_, _06254_, _06246_);
  nor (_06256_, _06247_, _06246_);
  nor (_06257_, _06252_, _06150_);
  nor (_06258_, _06257_, _06253_);
  and (_06259_, _06258_, _06256_);
  or (_06260_, _06236_, _06162_);
  and (_06261_, _06215_, _06213_);
  not (_06262_, _06261_);
  and (_06263_, _06262_, _06180_);
  nand (_06264_, _06263_, _06182_);
  or (_06265_, _06263_, _06182_);
  nand (_06266_, _06265_, _06264_);
  nand (_06267_, _06266_, _06236_);
  and (_06268_, _06267_, _06260_);
  nor (_06269_, _06268_, _06147_);
  not (_06270_, _06169_);
  nor (_06271_, _06215_, _06213_);
  nor (_06272_, _06271_, _06261_);
  or (_06273_, _06272_, _06238_);
  or (_06274_, _06236_, _06179_);
  and (_06275_, _06274_, _06273_);
  and (_06276_, _06275_, _06270_);
  and (_06277_, _06268_, _06147_);
  or (_06278_, _06277_, _06269_);
  not (_06279_, _06278_);
  and (_06280_, _06279_, _06276_);
  nor (_06281_, _06280_, _06269_);
  and (_06282_, _06211_, _06194_);
  not (_06283_, _06282_);
  and (_06284_, _06283_, _06212_);
  or (_06285_, _06284_, _06238_);
  or (_06286_, _06236_, _06191_);
  and (_06287_, _06286_, _06285_);
  nor (_06288_, _06287_, _06175_);
  not (_06289_, _06288_);
  or (_06290_, _06236_, _06206_);
  not (_06291_, _06202_);
  and (_06292_, _06206_, _06291_);
  nor (_06293_, _06206_, _06291_);
  nor (_06294_, _06293_, _06292_);
  nand (_06295_, _06236_, _06294_);
  nand (_06296_, _06295_, _06290_);
  nand (_06297_, _06296_, _06195_);
  or (_06298_, _06296_, _06195_);
  nand (_06299_, _06298_, _06297_);
  nor (_06300_, _06117_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_06301_, _06117_, _05943_);
  nor (_06302_, _06301_, _06300_);
  nor (_06303_, _06302_, _06291_);
  or (_06304_, _06303_, _06299_);
  and (_06305_, _06304_, _06297_);
  and (_06306_, _06209_, _06207_);
  not (_06307_, _06306_);
  and (_06309_, _06307_, _06210_);
  or (_06311_, _06309_, _06238_);
  or (_06313_, _06236_, _06200_);
  and (_06315_, _06313_, _06311_);
  nand (_06317_, _06315_, _06187_);
  or (_06319_, _06315_, _06187_);
  nand (_06321_, _06319_, _06317_);
  or (_06322_, _06321_, _06305_);
  and (_06323_, _06287_, _06175_);
  not (_06324_, _06323_);
  and (_06325_, _06324_, _06317_);
  nand (_06326_, _06325_, _06322_);
  and (_06327_, _06326_, _06289_);
  not (_06328_, _06276_);
  or (_06329_, _06275_, _06270_);
  and (_06330_, _06329_, _06328_);
  and (_06331_, _06279_, _06330_);
  nand (_06332_, _06331_, _06327_);
  nand (_06333_, _06332_, _06281_);
  and (_06334_, _06333_, _06259_);
  or (_06335_, _06334_, _06255_);
  and (_06336_, _06335_, _06230_);
  or (_06337_, _06336_, _06245_);
  and (_06338_, _06333_, _06258_);
  nor (_06339_, _06338_, _06253_);
  nand (_06340_, _06339_, _06256_);
  or (_06341_, _06339_, _06256_);
  nand (_06342_, _06341_, _06340_);
  nand (_06343_, _06342_, _06336_);
  nand (_06344_, _06343_, _06337_);
  and (_01068_, _06344_, _12493_);
  and (_02971_, _06336_, _12493_);
  and (_02980_, _06236_, _12493_);
  and (_02999_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _12493_);
  and (_03017_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _12493_);
  and (_03035_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _12493_);
  or (_06345_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_06346_, _06113_, rst);
  and (_03044_, _06346_, _06345_);
  not (_06347_, _06302_);
  and (_06349_, _06336_, _06202_);
  nor (_06350_, _06349_, _06347_);
  and (_06351_, _06349_, _06347_);
  or (_06352_, _06351_, _06350_);
  and (_03055_, _06352_, _12493_);
  nand (_06353_, _06335_, _06230_);
  and (_06354_, _06303_, _06299_);
  not (_06355_, _06354_);
  and (_06356_, _06355_, _06304_);
  or (_06357_, _06356_, _06353_);
  or (_06358_, _06336_, _06296_);
  and (_06359_, _06358_, _06357_);
  and (_03065_, _06359_, _12493_);
  not (_06360_, _06322_);
  and (_06361_, _06321_, _06305_);
  nor (_06362_, _06361_, _06360_);
  or (_06363_, _06362_, _06353_);
  or (_06364_, _06336_, _06315_);
  and (_06365_, _06364_, _06363_);
  and (_03074_, _06365_, _12493_);
  or (_06366_, _06323_, _06288_);
  and (_06367_, _06322_, _06317_);
  or (_06368_, _06367_, _06366_);
  nand (_06369_, _06367_, _06366_);
  nand (_06370_, _06369_, _06368_);
  nand (_06371_, _06370_, _06336_);
  or (_06372_, _06336_, _06287_);
  and (_06373_, _06372_, _06371_);
  and (_03083_, _06373_, _12493_);
  nand (_06374_, _06330_, _06327_);
  or (_06375_, _06330_, _06327_);
  nand (_06376_, _06375_, _06374_);
  nand (_06377_, _06376_, _06336_);
  or (_06378_, _06336_, _06275_);
  and (_06379_, _06378_, _06377_);
  and (_03093_, _06379_, _12493_);
  and (_06380_, _06374_, _06328_);
  nand (_06381_, _06278_, _06380_);
  or (_06382_, _06278_, _06380_);
  nand (_06383_, _06382_, _06381_);
  nand (_06384_, _06383_, _06336_);
  nand (_06385_, _06353_, _06268_);
  and (_06386_, _06385_, _06384_);
  and (_03103_, _06386_, _12493_);
  nor (_06387_, _06333_, _06258_);
  or (_06388_, _06387_, _06338_);
  nand (_06389_, _06388_, _06336_);
  or (_06390_, _06336_, _06252_);
  and (_06391_, _06390_, _06389_);
  and (_03113_, _06391_, _12493_);
  and (_06392_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06393_, _06392_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_06394_, _06393_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_06395_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_06396_, _06395_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_06397_, _06396_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_06398_, _06397_);
  not (_06399_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06400_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05610_);
  and (_06401_, _06400_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_06402_, _06401_, _06399_);
  not (_06403_, _06402_);
  nor (_06404_, _06396_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_06405_, _06404_, _06403_);
  and (_06406_, _06405_, _06398_);
  not (_06407_, _06406_);
  and (_06408_, _06401_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_06409_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_06410_, _06400_, _06409_);
  and (_06411_, _06410_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06412_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_06413_, _06412_, _06408_);
  not (_06414_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_06415_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05610_);
  and (_06416_, _06415_, _06399_);
  and (_06417_, _06416_, _06414_);
  and (_06418_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_06419_, _06410_, _06399_);
  and (_06420_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_06421_, _06420_, _06418_);
  and (_06422_, _06421_, _06413_);
  and (_06423_, _06422_, _06407_);
  nor (_06424_, _06395_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_06425_, _06424_);
  nor (_06426_, _06403_, _06396_);
  and (_06427_, _06426_, _06425_);
  not (_06428_, _06427_);
  and (_06429_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_06430_, _06429_, _06408_);
  and (_06431_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_06432_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_06433_, _06432_, _06431_);
  and (_06434_, _06433_, _06430_);
  and (_06435_, _06434_, _06428_);
  nor (_06436_, _06435_, _06423_);
  not (_06437_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_06438_, _06397_, _06437_);
  and (_06439_, _06397_, _06437_);
  nor (_06440_, _06439_, _06438_);
  nor (_06441_, _06440_, _06403_);
  not (_06442_, _06441_);
  and (_06443_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_06444_, _06443_);
  not (_06445_, _06408_);
  and (_06446_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_06447_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_06448_, _06447_, _06446_);
  and (_06449_, _06448_, _06445_);
  and (_06450_, _06449_, _06444_);
  and (_06451_, _06450_, _06442_);
  not (_06452_, _06451_);
  and (_06453_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_06454_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_06455_, _06454_, _06453_);
  not (_06456_, _06394_);
  nor (_06457_, _06393_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_06458_, _06457_, _06403_);
  and (_06459_, _06458_, _06456_);
  or (_06460_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06461_, _06460_, _05610_);
  nor (_06462_, _06461_, _06400_);
  and (_06463_, _06462_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_06464_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_06465_, _06464_, _06463_);
  not (_06466_, _06465_);
  nor (_06467_, _06466_, _06459_);
  and (_06468_, _06467_, _06455_);
  not (_06469_, _06468_);
  and (_06470_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_06471_, _06470_);
  and (_06472_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_06473_, _06472_, _06408_);
  and (_06474_, _06473_, _06471_);
  nor (_06475_, _06394_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_06476_, _06475_);
  nor (_06477_, _06403_, _06395_);
  and (_06478_, _06477_, _06476_);
  and (_06479_, _06462_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_06480_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_06481_, _06480_, _06479_);
  not (_06482_, _06481_);
  nor (_06483_, _06482_, _06478_);
  and (_06484_, _06483_, _06474_);
  nor (_06485_, _06484_, _06469_);
  and (_06486_, _06485_, _06452_);
  and (_06487_, _06486_, _06436_);
  and (_06488_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_06489_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_06490_, _06489_, _06488_);
  and (_06491_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_06492_, _06491_);
  not (_06493_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06494_, _06402_, _06493_);
  and (_06495_, _06462_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_06496_, _06495_, _06494_);
  and (_06497_, _06496_, _06492_);
  and (_06498_, _06497_, _06490_);
  nor (_06499_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_06500_, _06499_, _06392_);
  and (_06501_, _06500_, _06402_);
  and (_06502_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_06503_, _06502_, _06501_);
  and (_06504_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_06505_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_06506_, _06462_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_06507_, _06506_, _06505_);
  nor (_06508_, _06507_, _06504_);
  and (_06509_, _06508_, _06503_);
  nor (_06510_, _06392_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_06511_, _06510_, _06393_);
  and (_06512_, _06511_, _06402_);
  and (_06513_, _06417_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_06514_, _06513_, _06512_);
  and (_06515_, _06411_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_06516_, _06419_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_06517_, _06462_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_06518_, _06517_, _06516_);
  nor (_06519_, _06518_, _06515_);
  and (_06520_, _06519_, _06514_);
  and (_06521_, _06520_, _06509_);
  and (_06522_, _06521_, _06498_);
  nand (_06523_, _06522_, _06487_);
  nand (_06524_, _06344_, _06112_);
  nand (_06525_, _06053_, _05616_);
  not (_06526_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06527_, _05611_, _06526_);
  and (_06528_, _06527_, _05615_);
  not (_06529_, _06528_);
  nor (_06530_, _05865_, _05684_);
  and (_06531_, _05865_, _05684_);
  nor (_06532_, _06531_, _06530_);
  not (_06533_, _05743_);
  nor (_06534_, _05834_, _06533_);
  nor (_06535_, _05834_, _05743_);
  and (_06536_, _05834_, _05743_);
  nor (_06537_, _06536_, _06535_);
  not (_06538_, _05698_);
  nor (_06539_, _05813_, _06538_);
  nor (_06540_, _05813_, _05698_);
  and (_06541_, _05813_, _05698_);
  nor (_06543_, _06541_, _06540_);
  not (_06544_, _05750_);
  and (_06545_, _05667_, _06544_);
  nor (_06546_, _06545_, _06543_);
  nor (_06547_, _06546_, _06539_);
  nor (_06548_, _06547_, _06537_);
  nor (_06549_, _06548_, _06534_);
  and (_06550_, _06547_, _06537_);
  nor (_06551_, _06550_, _06548_);
  not (_06552_, _06551_);
  and (_06553_, _06545_, _06543_);
  nor (_06554_, _06553_, _06546_);
  not (_06555_, _06554_);
  nor (_06556_, _05667_, _05750_);
  and (_06557_, _05667_, _05750_);
  nor (_06558_, _06557_, _06556_);
  not (_06559_, _06558_);
  and (_06560_, _05795_, _05712_);
  nor (_06561_, _05795_, _05712_);
  nor (_06562_, _06561_, _06560_);
  not (_06563_, _05763_);
  and (_06564_, _05907_, _06563_);
  nor (_06565_, _05907_, _06563_);
  nor (_06566_, _06565_, _06564_);
  and (_06567_, _05892_, _05726_);
  nor (_06568_, _05892_, _05726_);
  nor (_06569_, _06568_, _06567_);
  and (_06570_, _05943_, _05777_);
  nor (_06571_, _06570_, _06569_);
  and (_06572_, _05892_, _06139_);
  nor (_06573_, _06572_, _06571_);
  nor (_06574_, _06573_, _06566_);
  and (_06575_, _05907_, _05763_);
  nor (_06576_, _06575_, _06574_);
  nor (_06577_, _06576_, _06562_);
  and (_06578_, _06576_, _06562_);
  nor (_06579_, _06578_, _06577_);
  not (_06580_, _06579_);
  and (_06581_, _06573_, _06566_);
  nor (_06582_, _06581_, _06574_);
  not (_06583_, _06582_);
  and (_06584_, _06570_, _06569_);
  nor (_06585_, _06584_, _06571_);
  not (_06586_, _06585_);
  not (_06587_, _05777_);
  nor (_06588_, _05943_, _06587_);
  and (_06589_, _05943_, _06587_);
  nor (_06590_, _06589_, _06588_);
  nor (_06591_, _05655_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_06592_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_06593_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_06594_, _06593_, _05672_);
  nor (_06595_, _06594_, _06592_);
  nor (_06596_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_06597_, _06596_, _05653_);
  not (_06598_, _06597_);
  not (_06599_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_06600_, _06599_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_06601_, _06600_, _05734_);
  not (_06602_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_06603_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _06602_);
  and (_06604_, _06603_, _05689_);
  nor (_06605_, _06604_, _06601_);
  and (_06606_, _06605_, _06598_);
  and (_06607_, _06606_, _06595_);
  and (_06608_, _06593_, _05703_);
  nor (_06609_, _06608_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_06610_, _06603_, _05717_);
  not (_06611_, _06610_);
  and (_06612_, _06600_, _05754_);
  and (_06613_, _06596_, _05768_);
  nor (_06614_, _06613_, _06612_);
  and (_06615_, _06614_, _06611_);
  and (_06616_, _06615_, _06609_);
  nor (_06617_, _06616_, _06607_);
  nor (_06618_, _06617_, _05649_);
  nor (_06619_, _06618_, _06591_);
  and (_06620_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_06621_, _06620_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_06622_, _06621_);
  and (_06623_, _06622_, _06619_);
  and (_06624_, _06622_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_06625_, _06624_, _06623_);
  nor (_06626_, _06625_, _06590_);
  and (_06627_, _06626_, _06586_);
  and (_06628_, _06627_, _06583_);
  and (_06629_, _06628_, _06580_);
  not (_06630_, _05712_);
  or (_06631_, _05795_, _06630_);
  and (_06632_, _05795_, _06630_);
  or (_06633_, _06576_, _06632_);
  and (_06634_, _06633_, _06631_);
  or (_06635_, _06634_, _06629_);
  and (_06636_, _06635_, _06559_);
  and (_06637_, _06636_, _06555_);
  and (_06638_, _06637_, _06552_);
  nor (_06639_, _06638_, _06549_);
  nor (_06640_, _06639_, _06532_);
  and (_06641_, _06639_, _06532_);
  nor (_06642_, _06641_, _06640_);
  nor (_06643_, _06642_, _06529_);
  not (_06644_, _06643_);
  not (_06645_, _06532_);
  not (_06646_, _06566_);
  and (_06647_, _06588_, _06569_);
  nor (_06648_, _06647_, _06567_);
  nor (_06649_, _06648_, _06646_);
  nor (_06650_, _06649_, _06564_);
  nor (_06651_, _06650_, _06562_);
  and (_06652_, _06650_, _06562_);
  nor (_06653_, _06652_, _06651_);
  not (_06654_, _06590_);
  nor (_06655_, _06625_, _06654_);
  and (_06656_, _06655_, _06569_);
  and (_06657_, _06648_, _06646_);
  nor (_06658_, _06657_, _06649_);
  and (_06659_, _06658_, _06656_);
  not (_06660_, _06659_);
  nor (_06661_, _06660_, _06653_);
  nor (_06662_, _06650_, _06560_);
  or (_06663_, _06662_, _06561_);
  or (_06664_, _06663_, _06661_);
  and (_06665_, _06664_, _06558_);
  and (_06666_, _06665_, _06543_);
  not (_06667_, _06537_);
  and (_06668_, _06556_, _06543_);
  nor (_06669_, _06668_, _06540_);
  nor (_06670_, _06669_, _06667_);
  and (_06671_, _06669_, _06667_);
  nor (_06672_, _06671_, _06670_);
  and (_06673_, _06672_, _06666_);
  nor (_06674_, _06670_, _06535_);
  not (_06675_, _06674_);
  nor (_06676_, _06675_, _06673_);
  and (_06677_, _06676_, _06645_);
  nor (_06678_, _06676_, _06645_);
  not (_06679_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_06680_, _06108_, _06679_);
  and (_06681_, _06680_, _05615_);
  not (_06682_, _06681_);
  or (_06683_, _06682_, _06678_);
  nor (_06684_, _06683_, _06677_);
  and (_06685_, _05614_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06686_, _06685_, _06527_);
  not (_06687_, _05892_);
  nor (_06688_, _05943_, _06687_);
  and (_06689_, _06688_, _05907_);
  and (_06690_, _06689_, _05796_);
  and (_06691_, _06690_, _05668_);
  and (_06692_, _06691_, _05814_);
  and (_06693_, _06692_, _05836_);
  and (_06694_, _06693_, _06625_);
  not (_06695_, _06625_);
  and (_06696_, _05834_, _05813_);
  nor (_06697_, _05907_, _05892_);
  and (_06698_, _06697_, _05943_);
  and (_06699_, _06698_, _05795_);
  and (_06700_, _06699_, _05667_);
  and (_06701_, _06700_, _06696_);
  and (_06702_, _06701_, _06695_);
  nor (_06703_, _06702_, _06694_);
  and (_06704_, _06703_, _05865_);
  nor (_06705_, _06703_, _05865_);
  nor (_06706_, _06705_, _06704_);
  and (_06707_, _06706_, _06686_);
  not (_06708_, _05684_);
  nor (_06709_, _06625_, _06708_);
  not (_06710_, _06709_);
  and (_06711_, _06625_, _05865_);
  and (_06712_, _06685_, _05612_);
  not (_06713_, _06712_);
  nor (_06714_, _06713_, _06711_);
  and (_06715_, _06714_, _06710_);
  nor (_06716_, _06715_, _06707_);
  and (_06717_, _06680_, _06111_);
  not (_06718_, _06717_);
  not (_06719_, _06696_);
  nor (_06720_, _06697_, _05795_);
  and (_06721_, _06720_, _06717_);
  and (_06722_, _06721_, _05668_);
  nor (_06723_, _06722_, _06719_);
  nor (_06724_, _06696_, _05865_);
  nor (_06725_, _06724_, _06721_);
  and (_06726_, _06725_, _06625_);
  nor (_06727_, _06726_, _06723_);
  and (_06728_, _06727_, _05865_);
  nor (_06729_, _06727_, _05865_);
  nor (_06730_, _06729_, _06728_);
  nor (_06731_, _06730_, _06718_);
  not (_06732_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06733_, _05614_, _06732_);
  and (_06734_, _06733_, _06109_);
  and (_06735_, _06734_, _06532_);
  and (_06736_, _06733_, _06680_);
  not (_06737_, _06736_);
  nor (_06738_, _06737_, _06531_);
  or (_06739_, _06738_, _06735_);
  not (_06740_, _06739_);
  and (_06741_, _06685_, _06680_);
  not (_06742_, _06741_);
  nor (_06743_, _06742_, _06625_);
  not (_06744_, _06743_);
  and (_06745_, _06109_, _05615_);
  not (_06746_, _06745_);
  nor (_06747_, _06746_, _05865_);
  and (_06748_, _06733_, _05611_);
  not (_06749_, _06748_);
  nor (_06750_, _06749_, _05834_);
  and (_06751_, _06685_, _06109_);
  and (_06752_, _06751_, _05944_);
  or (_06753_, _06752_, _06750_);
  nor (_06754_, _06753_, _06747_);
  and (_06755_, _06111_, _05612_);
  and (_06756_, _06755_, _06530_);
  and (_06757_, _06527_, _06111_);
  and (_06758_, _06757_, _05865_);
  nor (_06759_, _06758_, _06756_);
  and (_06760_, _06759_, _06754_);
  and (_06761_, _06760_, _06744_);
  and (_06762_, _06761_, _06740_);
  not (_06763_, _06762_);
  nor (_06764_, _06763_, _06731_);
  and (_06765_, _06764_, _06716_);
  not (_06766_, _06765_);
  nor (_06767_, _06766_, _06684_);
  and (_06768_, _06767_, _06644_);
  and (_06769_, _06768_, _06525_);
  and (_06770_, _06769_, _06524_);
  not (_06771_, _06770_);
  or (_06772_, _06771_, _06523_);
  not (_06773_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_06774_, \oc8051_top_1.oc8051_decoder1.wr , _05610_);
  not (_06775_, _06774_);
  nor (_06776_, _06775_, _06416_);
  and (_06777_, _06776_, _06773_);
  not (_06778_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_06779_, _06523_, _06778_);
  and (_06780_, _06779_, _06777_);
  and (_06781_, _06780_, _06772_);
  nor (_06782_, _06776_, _06778_);
  nor (_06783_, _06678_, _06530_);
  nor (_06784_, _06783_, _06682_);
  not (_06785_, _06784_);
  and (_06786_, _05865_, _06708_);
  nor (_06787_, _06786_, _06640_);
  nor (_06788_, _06787_, _06529_);
  and (_06789_, _06723_, _06625_);
  nor (_06790_, _06789_, _06711_);
  not (_06791_, _06723_);
  nor (_06792_, _06625_, _05865_);
  and (_06793_, _06792_, _06791_);
  nor (_06794_, _06793_, _06718_);
  and (_06795_, _06794_, _06790_);
  not (_06796_, _06795_);
  and (_06797_, _06621_, _06619_);
  and (_06798_, _06733_, _06527_);
  and (_06799_, _06755_, _06619_);
  nor (_06800_, _06799_, _06798_);
  nor (_06801_, _06800_, _06797_);
  not (_06802_, _06801_);
  nor (_06803_, _06746_, _06625_);
  not (_06804_, _06803_);
  and (_06805_, _06733_, _05612_);
  not (_06806_, _06805_);
  nor (_06807_, _06806_, _05865_);
  not (_06808_, _06807_);
  nor (_06809_, _06742_, _05943_);
  nor (_06810_, _06809_, _06721_);
  and (_06811_, _06810_, _06808_);
  and (_06812_, _06811_, _06804_);
  nor (_06813_, _06624_, _06619_);
  not (_06814_, _06734_);
  nor (_06815_, _06814_, _06623_);
  nor (_06816_, _06815_, _06736_);
  nor (_06817_, _06816_, _06813_);
  not (_06818_, _06624_);
  and (_06819_, _06757_, _06818_);
  and (_06820_, _06751_, _06624_);
  nor (_06821_, _06820_, _06819_);
  nor (_06822_, _06821_, _06623_);
  nor (_06823_, _06822_, _06817_);
  and (_06824_, _06823_, _06812_);
  and (_06825_, _06824_, _06802_);
  and (_06826_, _06825_, _06796_);
  not (_06827_, _06826_);
  nor (_06828_, _06827_, _06788_);
  and (_06829_, _06828_, _06785_);
  not (_06830_, _06498_);
  nor (_06831_, _06520_, _06509_);
  and (_06832_, _06831_, _06830_);
  and (_06833_, _06832_, _06487_);
  nand (_06834_, _06833_, _06829_);
  and (_06835_, _06776_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_06836_, _06833_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_06837_, _06836_, _06835_);
  and (_06838_, _06837_, _06834_);
  or (_06839_, _06838_, _06782_);
  or (_06840_, _06839_, _06781_);
  and (_05577_, _06840_, _12493_);
  nand (_06841_, _06352_, _06112_);
  and (_06842_, _06085_, _05616_);
  and (_06843_, _06625_, _06654_);
  nor (_06844_, _06843_, _06655_);
  not (_06845_, _06844_);
  nor (_06846_, _06681_, _06528_);
  nor (_06847_, _06846_, _06845_);
  not (_06848_, _06847_);
  nor (_06849_, _06806_, _06625_);
  not (_06850_, _06849_);
  nor (_06851_, _06814_, _06588_);
  nor (_06852_, _06851_, _06736_);
  or (_06853_, _06852_, _06589_);
  and (_06854_, _06755_, _06588_);
  not (_06855_, _06854_);
  and (_06856_, _06686_, _05943_);
  not (_06857_, _06856_);
  and (_06858_, _06712_, _05777_);
  and (_06859_, _06757_, _05943_);
  nor (_06860_, _06859_, _06858_);
  and (_06861_, _06860_, _06857_);
  and (_06862_, _06861_, _06855_);
  and (_06863_, _06685_, _06679_);
  and (_06864_, _06863_, _05892_);
  not (_06865_, _06864_);
  and (_06866_, _06798_, _05968_);
  nor (_06867_, _06745_, _06717_);
  nor (_06868_, _06867_, _05943_);
  nor (_06869_, _06868_, _06866_);
  and (_06870_, _06869_, _06865_);
  and (_06871_, _06870_, _06862_);
  and (_06872_, _06871_, _06853_);
  and (_06873_, _06872_, _06850_);
  and (_06874_, _06873_, _06848_);
  not (_06875_, _06874_);
  nor (_06876_, _06875_, _06842_);
  and (_06877_, _06876_, _06841_);
  not (_06878_, _06877_);
  or (_06879_, _06878_, _06523_);
  not (_06880_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_06881_, _06523_, _06880_);
  and (_06882_, _06881_, _06777_);
  and (_06883_, _06882_, _06879_);
  nor (_06884_, _06776_, _06880_);
  not (_06885_, _06829_);
  or (_06886_, _06885_, _06523_);
  and (_06887_, _06881_, _06835_);
  and (_06888_, _06887_, _06886_);
  or (_06889_, _06888_, _06884_);
  or (_06890_, _06889_, _06883_);
  and (_05578_, _06890_, _12493_);
  and (_06891_, _06090_, _05616_);
  not (_06892_, _06891_);
  nand (_06893_, _06359_, _06112_);
  nor (_06894_, _06588_, _06569_);
  or (_06895_, _06894_, _06647_);
  and (_06896_, _06895_, _06655_);
  nor (_06897_, _06895_, _06655_);
  or (_06898_, _06897_, _06896_);
  and (_06899_, _06898_, _06681_);
  nor (_06900_, _06626_, _06586_);
  nor (_06901_, _06900_, _06627_);
  nor (_06902_, _06901_, _06529_);
  not (_06903_, _06902_);
  nor (_06904_, _06720_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_06905_, _06904_, _05892_);
  nor (_06906_, _06904_, _05892_);
  nor (_06907_, _06906_, _06905_);
  nor (_06908_, _06907_, _06718_);
  not (_06909_, _06908_);
  and (_06910_, _06734_, _06569_);
  nor (_06911_, _06737_, _06568_);
  not (_06912_, _06911_);
  and (_06913_, _06755_, _06567_);
  and (_06914_, _06757_, _06687_);
  nor (_06915_, _06914_, _06913_);
  nand (_06916_, _06915_, _06912_);
  nor (_06917_, _06916_, _06910_);
  nor (_06918_, _06749_, _05943_);
  not (_06919_, _06918_);
  and (_06920_, _06745_, _05892_);
  and (_06921_, _06863_, _05907_);
  nor (_06922_, _06921_, _06920_);
  and (_06923_, _06922_, _06919_);
  and (_06924_, _06923_, _06917_);
  and (_06925_, _06924_, _06909_);
  and (_06926_, _06925_, _06903_);
  and (_06927_, _06712_, _05726_);
  and (_06928_, _05943_, _06687_);
  nor (_06929_, _06928_, _06688_);
  not (_06930_, _06929_);
  nor (_06931_, _06930_, _06625_);
  and (_06932_, _06930_, _06625_);
  nor (_06933_, _06932_, _06931_);
  and (_06934_, _06933_, _06686_);
  nor (_06935_, _06934_, _06927_);
  nand (_06936_, _06935_, _06926_);
  nor (_06937_, _06936_, _06899_);
  and (_06938_, _06937_, _06893_);
  and (_06939_, _06938_, _06892_);
  not (_06940_, _06939_);
  or (_06941_, _06940_, _06523_);
  not (_06942_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_06943_, _06523_, _06942_);
  and (_06944_, _06943_, _06777_);
  and (_06945_, _06944_, _06941_);
  nor (_06946_, _06776_, _06942_);
  and (_06947_, _06521_, _06830_);
  and (_06948_, _06947_, _06487_);
  or (_06949_, _06948_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_06950_, _06949_, _06835_);
  nand (_06951_, _06948_, _06829_);
  and (_06952_, _06951_, _06950_);
  or (_06953_, _06952_, _06946_);
  or (_06954_, _06953_, _06945_);
  and (_05579_, _06954_, _12493_);
  nand (_06955_, _06096_, _05616_);
  nand (_06956_, _06365_, _06112_);
  nor (_06957_, _06713_, _05763_);
  not (_06958_, _05907_);
  and (_06959_, _06928_, _06695_);
  and (_06960_, _06688_, _06625_);
  nor (_06961_, _06960_, _06959_);
  nor (_06962_, _06961_, _06958_);
  not (_06963_, _06686_);
  and (_06964_, _06961_, _06958_);
  or (_06965_, _06964_, _06963_);
  nor (_06966_, _06965_, _06962_);
  nor (_06967_, _06966_, _06957_);
  nor (_06968_, _06627_, _06583_);
  nor (_06969_, _06968_, _06628_);
  nor (_06970_, _06969_, _06529_);
  and (_06971_, _06734_, _06566_);
  nor (_06972_, _06737_, _06565_);
  not (_06973_, _06972_);
  and (_06974_, _06755_, _06564_);
  and (_06975_, _06757_, _06958_);
  nor (_06976_, _06975_, _06974_);
  nand (_06977_, _06976_, _06973_);
  nor (_06978_, _06977_, _06971_);
  and (_06979_, _06748_, _05892_);
  not (_06980_, _06979_);
  and (_06981_, _06745_, _05907_);
  not (_06982_, _06863_);
  nor (_06983_, _06982_, _05795_);
  nor (_06984_, _06983_, _06981_);
  and (_06985_, _06984_, _06980_);
  and (_06986_, _06985_, _06978_);
  not (_06987_, _06986_);
  nor (_06988_, _06987_, _06970_);
  nor (_06989_, _06658_, _06656_);
  nor (_06990_, _06989_, _06682_);
  and (_06991_, _06990_, _06660_);
  and (_06992_, _06697_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06993_, _06906_, _06958_);
  nor (_06994_, _06993_, _06992_);
  nor (_06995_, _06994_, _06718_);
  nor (_06996_, _06995_, _06991_);
  and (_06997_, _06996_, _06988_);
  and (_06998_, _06997_, _06967_);
  and (_06999_, _06998_, _06956_);
  and (_07000_, _06999_, _06955_);
  not (_07001_, _07000_);
  or (_07002_, _07001_, _06523_);
  not (_07003_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_07004_, _06523_, _07003_);
  and (_07005_, _07004_, _06777_);
  and (_07006_, _07005_, _07002_);
  nor (_07007_, _06776_, _07003_);
  nand (_07008_, _06520_, _06487_);
  nor (_07009_, _06509_, _06498_);
  or (_07010_, _07009_, _07008_);
  and (_07011_, _07010_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_07012_, _06509_);
  and (_07013_, _06520_, _07012_);
  and (_07014_, _07013_, _06498_);
  and (_07015_, _07014_, _06885_);
  and (_07016_, _06521_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_07017_, _07016_, _07015_);
  and (_07018_, _07017_, _06487_);
  or (_07019_, _07018_, _07011_);
  and (_07020_, _07019_, _06835_);
  or (_07021_, _07020_, _07007_);
  or (_07022_, _07021_, _07006_);
  and (_05580_, _07022_, _12493_);
  nand (_07023_, _06099_, _05616_);
  nand (_07024_, _06373_, _06112_);
  and (_07025_, _06660_, _06653_);
  or (_07026_, _07025_, _06682_);
  nor (_07027_, _07026_, _06661_);
  not (_07028_, _07027_);
  nor (_07029_, _06628_, _06580_);
  nor (_07030_, _07029_, _06629_);
  nor (_07031_, _07030_, _06529_);
  and (_07032_, _06755_, _06561_);
  and (_07033_, _06757_, _05795_);
  nor (_07034_, _07033_, _07032_);
  nor (_07035_, _06746_, _05795_);
  not (_07036_, _07035_);
  nor (_07037_, _06982_, _05667_);
  and (_07038_, _06748_, _05907_);
  nor (_07039_, _07038_, _07037_);
  and (_07040_, _07039_, _07036_);
  nand (_07041_, _07040_, _07034_);
  nor (_07042_, _07041_, _07031_);
  nor (_07043_, _06713_, _05712_);
  nor (_07044_, _06698_, _06625_);
  nor (_07045_, _06689_, _06695_);
  nor (_07046_, _07045_, _07044_);
  and (_07047_, _07046_, _05796_);
  nor (_07048_, _07046_, _05796_);
  or (_07049_, _07048_, _06963_);
  nor (_07050_, _07049_, _07047_);
  nor (_07051_, _07050_, _07043_);
  nor (_07052_, _06737_, _06560_);
  and (_07053_, _06734_, _06562_);
  nor (_07054_, _07053_, _07052_);
  not (_07055_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_07056_, _06697_, _07055_);
  nor (_07057_, _07056_, _05796_);
  or (_07058_, _07057_, _06718_);
  or (_07059_, _07058_, _06720_);
  and (_07060_, _07059_, _07054_);
  and (_07061_, _07060_, _07051_);
  and (_07062_, _07061_, _07042_);
  and (_07063_, _07062_, _07028_);
  and (_07064_, _07063_, _07024_);
  nand (_07065_, _07064_, _07023_);
  or (_07066_, _07065_, _06523_);
  not (_07067_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_07068_, _06523_, _07067_);
  and (_07069_, _07068_, _06777_);
  and (_07070_, _07069_, _07066_);
  nor (_07071_, _06776_, _07067_);
  and (_07072_, _07008_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_07073_, _07009_, _06520_);
  not (_07074_, _07073_);
  nor (_07075_, _07074_, _06829_);
  not (_07076_, _06520_);
  or (_07077_, _07009_, _07076_);
  nor (_07078_, _07077_, _07067_);
  or (_07079_, _07078_, _07075_);
  and (_07080_, _07079_, _06487_);
  or (_07081_, _07080_, _07072_);
  and (_07082_, _07081_, _06835_);
  or (_07083_, _07082_, _07071_);
  or (_07084_, _07083_, _07070_);
  and (_05581_, _07084_, _12493_);
  nand (_07085_, _06379_, _06112_);
  nand (_07086_, _06102_, _05616_);
  nor (_07087_, _06635_, _06558_);
  and (_07088_, _06635_, _06558_);
  nor (_07089_, _07088_, _07087_);
  and (_07090_, _07089_, _06528_);
  not (_07091_, _07090_);
  nor (_07092_, _06664_, _06558_);
  nor (_07093_, _07092_, _06665_);
  and (_07094_, _07093_, _06681_);
  and (_07095_, _06625_, _05668_);
  nor (_07096_, _06625_, _05750_);
  or (_07097_, _07096_, _07095_);
  and (_07098_, _07097_, _06712_);
  and (_07099_, _06690_, _06625_);
  and (_07100_, _06699_, _06695_);
  nor (_07101_, _07100_, _07099_);
  nor (_07102_, _07101_, _05667_);
  not (_07103_, _07102_);
  and (_07104_, _07101_, _05667_);
  nor (_07105_, _07104_, _06963_);
  and (_07106_, _07105_, _07103_);
  nor (_07107_, _07106_, _07098_);
  nor (_07108_, _06721_, _05668_);
  not (_07109_, _07108_);
  nor (_07110_, _06722_, _06718_);
  and (_07111_, _07110_, _07109_);
  not (_07112_, _07111_);
  and (_07113_, _06734_, _06558_);
  nor (_07114_, _06737_, _06557_);
  not (_07115_, _07114_);
  and (_07116_, _06755_, _06556_);
  and (_07117_, _06757_, _05667_);
  nor (_07118_, _07117_, _07116_);
  nand (_07119_, _07118_, _07115_);
  nor (_07120_, _07119_, _07113_);
  nor (_07121_, _06982_, _05813_);
  not (_07122_, _07121_);
  nor (_07123_, _06746_, _05667_);
  nor (_07124_, _06749_, _05795_);
  nor (_07125_, _07124_, _07123_);
  and (_07126_, _07125_, _07122_);
  and (_07127_, _07126_, _07120_);
  and (_07128_, _07127_, _07112_);
  and (_07129_, _07128_, _07107_);
  not (_07130_, _07129_);
  nor (_07131_, _07130_, _07094_);
  and (_07132_, _07131_, _07091_);
  and (_07133_, _07132_, _07086_);
  and (_07134_, _07133_, _07085_);
  not (_07135_, _07134_);
  or (_07136_, _07135_, _06523_);
  not (_07137_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_07138_, _06523_, _07137_);
  and (_07139_, _07138_, _06777_);
  and (_07140_, _07139_, _07136_);
  nor (_07141_, _06776_, _07137_);
  not (_07142_, _06487_);
  and (_07143_, _06509_, _06498_);
  and (_07144_, _07143_, _07076_);
  nor (_07145_, _07143_, _07076_);
  nor (_07146_, _07145_, _07144_);
  or (_07147_, _07146_, _07142_);
  and (_07148_, _07147_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_07149_, _07144_);
  nor (_07150_, _07149_, _06829_);
  and (_07151_, _07145_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_07152_, _07151_, _07150_);
  and (_07153_, _07152_, _06487_);
  or (_07154_, _07153_, _07148_);
  and (_07155_, _07154_, _06835_);
  or (_07156_, _07155_, _07141_);
  or (_07157_, _07156_, _07140_);
  and (_05582_, _07157_, _12493_);
  nand (_07158_, _06105_, _05616_);
  nand (_07159_, _06386_, _06112_);
  nor (_07160_, _06636_, _06555_);
  nor (_07161_, _07160_, _06637_);
  nor (_07162_, _07161_, _06529_);
  not (_07163_, _07162_);
  nor (_07164_, _06556_, _06543_);
  or (_07165_, _07164_, _06668_);
  and (_07166_, _07165_, _06665_);
  nor (_07167_, _07165_, _06665_);
  or (_07168_, _07167_, _07166_);
  and (_07169_, _07168_, _06681_);
  nor (_07170_, _06691_, _06695_);
  nor (_07171_, _06700_, _06625_);
  nor (_07172_, _07171_, _07170_);
  nor (_07173_, _07172_, _05814_);
  not (_07174_, _07173_);
  and (_07175_, _07172_, _05814_);
  nor (_07176_, _07175_, _06963_);
  and (_07177_, _07176_, _07174_);
  nor (_07178_, _06625_, _05698_);
  and (_07179_, _06625_, _05814_);
  nor (_07180_, _07179_, _07178_);
  nor (_07181_, _07180_, _06713_);
  nor (_07182_, _06737_, _06541_);
  and (_07183_, _06734_, _06543_);
  nor (_07184_, _07183_, _07182_);
  not (_07185_, _07184_);
  nor (_07186_, _07185_, _07181_);
  not (_07187_, _07186_);
  nor (_07188_, _07187_, _07177_);
  nor (_07189_, _06722_, _05814_);
  not (_07190_, _06726_);
  and (_07191_, _07190_, _07189_);
  nor (_07192_, _06726_, _06722_);
  nor (_07193_, _07192_, _05813_);
  nor (_07194_, _07193_, _07191_);
  nor (_07195_, _07194_, _06718_);
  and (_07196_, _06755_, _06540_);
  and (_07197_, _06757_, _05813_);
  nor (_07198_, _07197_, _07196_);
  nor (_07199_, _06982_, _05834_);
  not (_07200_, _07199_);
  nor (_07201_, _06746_, _05813_);
  nor (_07202_, _06749_, _05667_);
  nor (_07203_, _07202_, _07201_);
  and (_07204_, _07203_, _07200_);
  and (_07205_, _07204_, _07198_);
  not (_07206_, _07205_);
  nor (_07207_, _07206_, _07195_);
  and (_07208_, _07207_, _07188_);
  not (_07209_, _07208_);
  nor (_07210_, _07209_, _07169_);
  and (_07211_, _07210_, _07163_);
  and (_07212_, _07211_, _07159_);
  nand (_07213_, _07212_, _07158_);
  or (_07214_, _07213_, _06523_);
  not (_07215_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_07216_, _06523_, _07215_);
  and (_07217_, _07216_, _06777_);
  and (_07218_, _07217_, _07214_);
  nor (_07219_, _06776_, _07215_);
  and (_07220_, _07076_, _06509_);
  nor (_07221_, _07220_, _07013_);
  or (_07222_, _07221_, _07142_);
  and (_07223_, _07222_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_07224_, _06509_, _06830_);
  and (_07225_, _07224_, _07076_);
  not (_07226_, _07225_);
  nor (_07227_, _07226_, _06829_);
  or (_07228_, _07144_, _07013_);
  and (_07229_, _07228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_07230_, _07229_, _07227_);
  and (_07231_, _07230_, _06487_);
  or (_07232_, _07231_, _07223_);
  and (_07233_, _07232_, _06835_);
  or (_07234_, _07233_, _07219_);
  or (_07235_, _07234_, _07218_);
  and (_05583_, _07235_, _12493_);
  nand (_07236_, _06391_, _06112_);
  nand (_07237_, _06107_, _05616_);
  nor (_07238_, _06637_, _06552_);
  nor (_07239_, _07238_, _06638_);
  nor (_07240_, _07239_, _06529_);
  not (_07241_, _07240_);
  nor (_07242_, _06672_, _06666_);
  not (_07243_, _07242_);
  nor (_07244_, _06682_, _06673_);
  and (_07245_, _07244_, _07243_);
  and (_07246_, _06625_, _05836_);
  nor (_07247_, _06625_, _05743_);
  or (_07248_, _07247_, _07246_);
  and (_07249_, _07248_, _06712_);
  nor (_07250_, _06625_, _05814_);
  nand (_07251_, _07250_, _06700_);
  nand (_07252_, _06692_, _06625_);
  and (_07253_, _07252_, _07251_);
  nor (_07254_, _07253_, _05834_);
  not (_07255_, _07254_);
  and (_07256_, _07253_, _05834_);
  nor (_07257_, _07256_, _06963_);
  and (_07258_, _07257_, _07255_);
  nor (_07259_, _07258_, _07249_);
  nor (_07260_, _07191_, _05834_);
  and (_07261_, _07191_, _05834_);
  nor (_07262_, _07261_, _07260_);
  nor (_07263_, _07262_, _06718_);
  nor (_07264_, _06737_, _06536_);
  and (_07265_, _06734_, _06537_);
  nor (_07266_, _07265_, _07264_);
  and (_07267_, _06755_, _06535_);
  and (_07268_, _06757_, _05834_);
  nor (_07269_, _07268_, _07267_);
  nor (_07270_, _06746_, _05834_);
  not (_07271_, _07270_);
  nor (_07272_, _06982_, _05865_);
  nor (_07273_, _06749_, _05813_);
  nor (_07274_, _07273_, _07272_);
  and (_07275_, _07274_, _07271_);
  and (_07276_, _07275_, _07269_);
  and (_07277_, _07276_, _07266_);
  not (_07278_, _07277_);
  nor (_07279_, _07278_, _07263_);
  and (_07280_, _07279_, _07259_);
  not (_07281_, _07280_);
  nor (_07282_, _07281_, _07245_);
  and (_07283_, _07282_, _07241_);
  and (_07284_, _07283_, _07237_);
  and (_07285_, _07284_, _07236_);
  not (_07286_, _07285_);
  or (_07287_, _07286_, _06523_);
  not (_07288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_07289_, _06523_, _07288_);
  and (_07290_, _07289_, _06777_);
  and (_07291_, _07290_, _07287_);
  nor (_07292_, _06776_, _07288_);
  not (_07293_, _06832_);
  nand (_07294_, _07293_, _06487_);
  and (_07295_, _07294_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_07296_, _06831_, _06498_);
  not (_07297_, _07296_);
  nor (_07298_, _07297_, _06829_);
  nor (_07299_, _06831_, _07288_);
  or (_07300_, _07299_, _07298_);
  and (_07301_, _07300_, _06487_);
  or (_07302_, _07301_, _07295_);
  and (_07303_, _07302_, _06835_);
  or (_07304_, _07303_, _07292_);
  or (_07305_, _07304_, _07291_);
  and (_05584_, _07305_, _12493_);
  and (_07306_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_07307_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_07308_, _07307_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_07309_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_07310_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_07311_, _07310_, _07309_);
  and (_07312_, _07307_, _05610_);
  and (_07313_, _07312_, _07311_);
  not (_07314_, _07313_);
  and (_07315_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_07316_, _07315_);
  not (_07317_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_07318_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_07319_, _07318_);
  not (_07320_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not (_07321_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_07322_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07323_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _07322_);
  nand (_07324_, _07323_, _07321_);
  or (_07325_, _07324_, _07320_);
  not (_07326_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  not (_07327_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_07328_, _07327_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_07329_, _07328_, _07321_);
  or (_07331_, _07329_, _07326_);
  and (_07332_, _07331_, _07325_);
  nor (_07334_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_07335_, _07334_, _07321_);
  nand (_07337_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_07338_, _07334_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_07340_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_07341_, _07340_, _07337_);
  and (_07342_, _07334_, _07321_);
  nand (_07343_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_07344_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07345_, _07344_, _07321_);
  nand (_07346_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_07347_, _07346_, _07343_);
  and (_07348_, _07347_, _07341_);
  nand (_07349_, _07348_, _07332_);
  nand (_07350_, _07349_, _07319_);
  nand (_07351_, _07350_, _07317_);
  nor (_07352_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07317_);
  nor (_07353_, _07352_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_07354_, _07353_, _07351_);
  and (_07355_, _07354_, _07316_);
  or (_07356_, _07355_, _07314_);
  and (_07357_, _07311_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_07358_, _07357_, _07314_);
  not (_07359_, _07358_);
  and (_07360_, _07359_, _07356_);
  and (_07361_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_07362_, _07361_);
  not (_07363_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_07364_, _07329_, _07363_);
  not (_07365_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_07366_, _07324_, _07365_);
  and (_07367_, _07366_, _07364_);
  nand (_07368_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_07369_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_07370_, _07369_, _07368_);
  nand (_07371_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_07372_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_07373_, _07372_, _07371_);
  and (_07374_, _07373_, _07370_);
  and (_07375_, _07374_, _07367_);
  or (_07376_, _07375_, _07318_);
  nand (_07377_, _07376_, _07317_);
  nor (_07378_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _07317_);
  nor (_07379_, _07378_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_07380_, _07379_, _07377_);
  and (_07381_, _07380_, _07362_);
  or (_07382_, _07381_, _07314_);
  and (_07383_, _07311_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_07384_, _07383_, _07314_);
  not (_07385_, _07384_);
  and (_07386_, _07385_, _07382_);
  and (_07387_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_07388_, _07387_);
  not (_07389_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_07390_, _07324_, _07389_);
  not (_07391_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_07392_, _07329_, _07391_);
  and (_07393_, _07392_, _07390_);
  nand (_07394_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_07395_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_07396_, _07395_, _07394_);
  nand (_07397_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_07398_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_07399_, _07398_, _07397_);
  and (_07400_, _07399_, _07396_);
  nand (_07401_, _07400_, _07393_);
  nand (_07402_, _07401_, _07319_);
  nand (_07403_, _07402_, _07317_);
  nor (_07404_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07317_);
  nor (_07405_, _07404_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_07406_, _07405_, _07403_);
  and (_07407_, _07406_, _07388_);
  or (_07408_, _07407_, _07314_);
  and (_07409_, _07311_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_07410_, _07409_, _07314_);
  not (_07411_, _07410_);
  and (_07412_, _07411_, _07408_);
  and (_07413_, _07412_, _07386_);
  and (_07414_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_07415_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_07416_, _07415_, _07414_);
  not (_07417_, _07324_);
  and (_07418_, _07417_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_07419_, _07418_, _07416_);
  not (_07420_, _07329_);
  and (_07421_, _07420_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_07422_, _07421_, _07318_);
  and (_07423_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_07424_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_07425_, _07424_, _07423_);
  or (_07426_, _07425_, _07422_);
  or (_07427_, _07426_, _07419_);
  or (_07428_, _07427_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_07429_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07317_);
  nor (_07430_, _07429_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_07431_, _07430_, _07428_);
  and (_07432_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_07433_, _07432_, _07431_);
  nand (_07434_, _07433_, _07313_);
  and (_07435_, _07311_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_07436_, _07435_, _07314_);
  not (_07437_, _07436_);
  and (_07438_, _07437_, _07434_);
  not (_07439_, _07438_);
  and (_07440_, _07439_, _07413_);
  and (_07441_, _07440_, _07360_);
  and (_07442_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not (_07443_, _07442_);
  nand (_07444_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not (_07445_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_07446_, _07329_, _07445_);
  and (_07447_, _07446_, _07444_);
  nand (_07448_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  not (_07449_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_07450_, _07324_, _07449_);
  and (_07451_, _07450_, _07448_);
  and (_07452_, _07451_, _07447_);
  nand (_07453_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_07454_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_07455_, _07454_, _07453_);
  and (_07456_, _07455_, _07452_);
  or (_07457_, _07456_, _07318_);
  nand (_07458_, _07457_, _07317_);
  nor (_07459_, _07317_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nor (_07460_, _07459_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_07461_, _07460_, _07458_);
  and (_07462_, _07461_, _07443_);
  or (_07463_, _07462_, _07314_);
  and (_07464_, _07311_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_07465_, _07464_, _07314_);
  not (_07466_, _07465_);
  and (_07467_, _07466_, _07463_);
  and (_07468_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_07469_, _07468_);
  nand (_07470_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not (_07471_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_07472_, _07329_, _07471_);
  and (_07473_, _07472_, _07470_);
  nand (_07474_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not (_07475_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_07476_, _07324_, _07475_);
  and (_07477_, _07476_, _07474_);
  and (_07478_, _07477_, _07473_);
  nand (_07479_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_07480_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_07481_, _07480_, _07479_);
  and (_07482_, _07481_, _07478_);
  or (_07483_, _07482_, _07318_);
  nand (_07484_, _07483_, _07317_);
  nor (_07485_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07317_);
  nor (_07486_, _07485_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_07487_, _07486_, _07484_);
  and (_07488_, _07487_, _07469_);
  or (_07489_, _07488_, _07314_);
  and (_07490_, _07311_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_07491_, _07490_, _07314_);
  not (_07492_, _07491_);
  and (_07493_, _07492_, _07489_);
  and (_07494_, _07493_, _07467_);
  and (_07495_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_07496_, _07495_);
  nand (_07497_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_07498_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_07499_, _07324_, _07498_);
  and (_07500_, _07499_, _07497_);
  nand (_07501_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_07502_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_07503_, _07502_, _07501_);
  nand (_07504_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not (_07505_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_07506_, _07329_, _07505_);
  and (_07507_, _07506_, _07504_);
  and (_07508_, _07507_, _07503_);
  nand (_07509_, _07508_, _07500_);
  and (_07510_, _07509_, _07319_);
  or (_07511_, _07510_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_07512_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07317_);
  nor (_07513_, _07512_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_07514_, _07513_, _07511_);
  and (_07515_, _07514_, _07496_);
  or (_07516_, _07515_, _07314_);
  and (_07517_, _07311_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_07518_, _07517_, _07314_);
  not (_07519_, _07518_);
  and (_07520_, _07519_, _07516_);
  not (_07521_, _07520_);
  and (_07522_, _07521_, _07494_);
  and (_07523_, _07522_, _07441_);
  nand (_07524_, _07492_, _07489_);
  and (_07525_, _07524_, _07467_);
  and (_07526_, _07525_, _07521_);
  and (_07527_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_07528_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_07529_, _07528_, _07527_);
  not (_07530_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_07531_, _07324_, _07530_);
  and (_07532_, _07531_, _07319_);
  and (_07533_, _07532_, _07529_);
  and (_07534_, _07420_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_07535_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_07536_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_07537_, _07536_, _07535_);
  not (_07538_, _07537_);
  nor (_07539_, _07538_, _07534_);
  nand (_07540_, _07539_, _07533_);
  or (_07541_, _07540_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_07542_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07317_);
  nor (_07543_, _07542_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_07544_, _07543_, _07541_);
  and (_07545_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_07546_, _07545_, _07544_);
  nand (_07547_, _07546_, _07313_);
  and (_07548_, _07311_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_07549_, _07548_, _07314_);
  not (_07550_, _07549_);
  and (_07551_, _07550_, _07547_);
  not (_07552_, _07386_);
  and (_07553_, _07412_, _07552_);
  and (_07554_, _07553_, _07439_);
  and (_07555_, _07554_, _07551_);
  and (_07556_, _07555_, _07526_);
  nor (_07557_, _07556_, _07523_);
  and (_07558_, _07438_, _07360_);
  and (_07559_, _07558_, _07413_);
  not (_07560_, _07551_);
  nand (_07561_, _07466_, _07463_);
  and (_07562_, _07520_, _07524_);
  and (_07563_, _07562_, _07561_);
  and (_07564_, _07563_, _07560_);
  and (_07565_, _07564_, _07559_);
  and (_07566_, _07493_, _07561_);
  and (_07567_, _07566_, _07521_);
  nor (_07568_, _07438_, _07386_);
  and (_07569_, _07560_, _07412_);
  and (_07570_, _07569_, _07568_);
  and (_07571_, _07570_, _07567_);
  and (_07572_, _07520_, _07494_);
  and (_07573_, _07572_, _07554_);
  nor (_07574_, _07573_, _07571_);
  not (_07575_, _07574_);
  nor (_07576_, _07575_, _07565_);
  and (_07577_, _07576_, _07557_);
  not (_07578_, _07554_);
  and (_07579_, _07525_, _07520_);
  and (_07580_, _07579_, _07560_);
  nor (_07581_, _07580_, _07522_);
  nor (_07582_, _07581_, _07578_);
  and (_07583_, _07563_, _07554_);
  and (_07584_, _07566_, _07520_);
  and (_07585_, _07584_, _07570_);
  nor (_07586_, _07585_, _07583_);
  not (_07587_, _07586_);
  and (_07588_, _07551_, _07520_);
  and (_07589_, _07588_, _07566_);
  and (_07590_, _07589_, _07554_);
  or (_07591_, _07590_, _07587_);
  nor (_07592_, _07591_, _07582_);
  and (_07593_, _07592_, _07577_);
  nor (_07594_, _07520_, _07493_);
  and (_07595_, _07594_, _07561_);
  and (_07596_, _07595_, _07555_);
  and (_07597_, _07562_, _07555_);
  and (_07598_, _07597_, _07467_);
  nor (_07599_, _07598_, _07596_);
  and (_07600_, _07567_, _07551_);
  not (_07601_, _07360_);
  and (_07602_, _07440_, _07601_);
  and (_07603_, _07602_, _07600_);
  not (_07604_, _07603_);
  and (_07605_, _07526_, _07560_);
  and (_07606_, _07605_, _07602_);
  and (_07607_, _07584_, _07560_);
  and (_07608_, _07602_, _07607_);
  nor (_07609_, _07608_, _07606_);
  and (_07610_, _07609_, _07604_);
  and (_07611_, _07610_, _07599_);
  and (_07612_, _07611_, _07593_);
  nor (_07613_, _07612_, _07308_);
  not (_07614_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_07615_, _05610_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_07616_, _07615_, _07614_);
  and (_07617_, _07616_, _07526_);
  and (_07618_, _07617_, _07559_);
  and (_07619_, _07523_, _07615_);
  and (_07620_, _07619_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_07621_, _07620_, _07618_);
  nor (_07622_, _07621_, _07613_);
  nor (_07623_, _07622_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_07624_, _07623_, _07306_);
  and (_07625_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_07626_, _07567_, _07555_);
  not (_07627_, _07626_);
  and (_07628_, _07438_, _07601_);
  and (_07629_, _07628_, _07553_);
  and (_07630_, _07595_, _07551_);
  and (_07631_, _07630_, _07629_);
  and (_07632_, _07566_, _07560_);
  and (_07633_, _07632_, _07629_);
  nor (_07634_, _07633_, _07631_);
  and (_07635_, _07634_, _07627_);
  and (_07636_, _07563_, _07559_);
  and (_07637_, _07526_, _07551_);
  and (_07638_, _07637_, _07440_);
  nor (_07639_, _07638_, _07636_);
  not (_07640_, _07523_);
  and (_07641_, _07588_, _07494_);
  and (_07642_, _07641_, _07629_);
  not (_07643_, _07412_);
  and (_07644_, _07600_, _07643_);
  nor (_07645_, _07644_, _07642_);
  and (_07646_, _07645_, _07640_);
  and (_07647_, _07646_, _07639_);
  not (_07648_, _07629_);
  nor (_07649_, _07648_, _07581_);
  not (_07650_, _07649_);
  and (_07651_, _07559_, _07522_);
  and (_07652_, _07651_, _07551_);
  not (_07653_, _07559_);
  and (_07654_, _07560_, _07522_);
  and (_07655_, _07572_, _07560_);
  nor (_07656_, _07655_, _07654_);
  nor (_07657_, _07656_, _07653_);
  nor (_07658_, _07657_, _07652_);
  and (_07659_, _07658_, _07650_);
  and (_07660_, _07659_, _07647_);
  and (_07661_, _07660_, _07635_);
  and (_07662_, _07588_, _07525_);
  and (_07663_, _07662_, _07440_);
  not (_07664_, _07663_);
  and (_07665_, _07655_, _07629_);
  and (_07666_, _07567_, _07560_);
  and (_07667_, _07666_, _07559_);
  nor (_07668_, _07667_, _07665_);
  and (_07669_, _07668_, _07664_);
  and (_07670_, _07605_, _07441_);
  and (_07671_, _07629_, _07564_);
  nor (_07672_, _07671_, _07670_);
  and (_07673_, _07672_, _07669_);
  and (_07674_, _07662_, _07629_);
  and (_07675_, _07600_, _07559_);
  nor (_07676_, _07675_, _07674_);
  and (_07677_, _07666_, _07441_);
  and (_07678_, _07563_, _07551_);
  and (_07679_, _07678_, _07441_);
  nor (_07680_, _07679_, _07677_);
  and (_07681_, _07680_, _07676_);
  and (_07682_, _07681_, _07673_);
  and (_07683_, _07589_, _07441_);
  and (_07684_, _07580_, _07440_);
  nor (_07685_, _07684_, _07683_);
  and (_07686_, _07629_, _07637_);
  and (_07687_, _07678_, _07629_);
  nor (_07688_, _07687_, _07686_);
  and (_07689_, _07688_, _07685_);
  and (_07690_, _07564_, _07441_);
  and (_07691_, _07600_, _07441_);
  nor (_07692_, _07691_, _07690_);
  and (_07693_, _07607_, _07441_);
  and (_07694_, _07629_, _07589_);
  nor (_07695_, _07694_, _07693_);
  and (_07696_, _07695_, _07692_);
  and (_07697_, _07696_, _07689_);
  and (_07698_, _07697_, _07682_);
  and (_07699_, _07698_, _07661_);
  nor (_07700_, _07699_, _07308_);
  and (_07701_, _07615_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_07702_, _07701_, _07523_);
  not (_07703_, _07702_);
  and (_07704_, _07559_, _07525_);
  and (_07705_, _07704_, _07616_);
  not (_07706_, _07616_);
  nor (_07707_, _07560_, _07520_);
  and (_07708_, _07707_, _07494_);
  nand (_07709_, _07559_, _07708_);
  nand (_07710_, _07655_, _07559_);
  and (_07711_, _07710_, _07709_);
  nor (_07712_, _07711_, _07706_);
  nor (_07713_, _07712_, _07705_);
  and (_07714_, _07713_, _07703_);
  not (_07715_, _07714_);
  nor (_07716_, _07715_, _07700_);
  nor (_07717_, _07716_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_07718_, _07717_, _07625_);
  nor (_07719_, _07718_, _07624_);
  and (_07720_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_07721_, _07558_, _07553_);
  and (_07722_, _07721_, _07589_);
  and (_07723_, _07721_, _07600_);
  nor (_07724_, _07723_, _07722_);
  and (_07725_, _07724_, _07610_);
  nor (_07726_, _07725_, _07308_);
  not (_07727_, _07308_);
  nor (_07728_, _07724_, _07727_);
  nor (_07729_, _07728_, _07705_);
  not (_07730_, _07729_);
  nor (_07731_, _07730_, _07726_);
  nor (_07732_, _07731_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_07733_, _07732_, _07720_);
  and (_07734_, _07733_, _12493_);
  and (_05585_, _07734_, _07719_);
  and (_07735_, _06435_, _06423_);
  not (_07736_, _06484_);
  nor (_07737_, _07736_, _06451_);
  and (_07738_, _07737_, _07735_);
  and (_07739_, _07738_, _06947_);
  and (_07740_, _06777_, _06468_);
  and (_07741_, _07740_, _07739_);
  not (_07742_, _07741_);
  and (_07743_, _07742_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_07744_, _06112_, _05616_);
  and (_07745_, _06680_, _06110_);
  nor (_07746_, _06745_, _07745_);
  and (_07747_, _07746_, _07744_);
  nor (_07748_, _06863_, _06748_);
  and (_07749_, _07748_, _07747_);
  nor (_07750_, _07749_, _05834_);
  not (_07751_, _07750_);
  and (_07752_, _07751_, _07269_);
  and (_07753_, _07752_, _07266_);
  and (_07754_, _07753_, _07259_);
  nor (_07755_, _07754_, _07742_);
  nor (_07756_, _07755_, _07743_);
  and (_07757_, _07742_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_07758_, _07749_, _05813_);
  not (_07759_, _07758_);
  and (_07760_, _07759_, _07198_);
  and (_07761_, _07760_, _07188_);
  nor (_07762_, _07761_, _07742_);
  nor (_07763_, _07762_, _07757_);
  and (_07764_, _07742_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_07765_, _07749_, _05667_);
  not (_07766_, _07765_);
  and (_07767_, _07766_, _07120_);
  and (_07768_, _07767_, _07107_);
  nor (_07769_, _07768_, _07742_);
  nor (_07770_, _07769_, _07764_);
  and (_07771_, _07742_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_07772_, _07749_, _05795_);
  not (_07773_, _07772_);
  and (_07774_, _07773_, _07034_);
  and (_07775_, _07774_, _07054_);
  and (_07776_, _07775_, _07051_);
  nor (_07777_, _07776_, _07742_);
  nor (_07778_, _07777_, _07771_);
  and (_07779_, _07742_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_07780_, _07749_, _06958_);
  not (_07781_, _07780_);
  and (_07782_, _07781_, _06978_);
  and (_07783_, _07782_, _06967_);
  nor (_07784_, _07783_, _07742_);
  nor (_07785_, _07784_, _07779_);
  and (_07786_, _07742_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_07787_, _07749_, _06687_);
  not (_07788_, _07787_);
  and (_07789_, _07788_, _06917_);
  and (_07790_, _07789_, _06935_);
  nor (_07791_, _07790_, _07742_);
  nor (_07792_, _07791_, _07786_);
  nor (_07793_, _07741_, _06493_);
  nor (_07794_, _07749_, _05943_);
  not (_07795_, _07794_);
  and (_07796_, _07795_, _06862_);
  and (_07797_, _07796_, _06853_);
  not (_07798_, _07797_);
  and (_07799_, _07798_, _07741_);
  nor (_07800_, _07799_, _07793_);
  and (_07801_, _07800_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_07802_, _07801_, _07792_);
  and (_07803_, _07802_, _07785_);
  and (_07804_, _07803_, _07778_);
  and (_07805_, _07804_, _07770_);
  and (_07806_, _07805_, _07763_);
  and (_07807_, _07806_, _07756_);
  nor (_07808_, _07741_, _06437_);
  nand (_07809_, _07808_, _07807_);
  or (_07810_, _07808_, _07807_);
  and (_07811_, _07810_, _06403_);
  and (_07812_, _07811_, _07809_);
  or (_07813_, _07812_, _06441_);
  and (_07814_, _07813_, _07742_);
  or (_07815_, _07749_, _05865_);
  and (_07816_, _07815_, _06740_);
  and (_07817_, _07816_, _06759_);
  and (_07818_, _07817_, _06716_);
  nor (_07819_, _07818_, _07742_);
  or (_07820_, _07819_, _07814_);
  and (_05586_, _07820_, _12493_);
  not (_07821_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_07822_, _07800_, _07821_);
  nor (_07823_, _07800_, _07821_);
  nor (_07824_, _07823_, _07822_);
  and (_07825_, _07824_, _06403_);
  nor (_07826_, _07825_, _06494_);
  nor (_07827_, _07826_, _07741_);
  nor (_07828_, _07827_, _07799_);
  nand (_05587_, _07828_, _12493_);
  nor (_07829_, _07801_, _07792_);
  nor (_07830_, _07829_, _07802_);
  nor (_07831_, _07830_, _06402_);
  nor (_07832_, _07831_, _06501_);
  nor (_07833_, _07832_, _07741_);
  nor (_07834_, _07833_, _07791_);
  nand (_05588_, _07834_, _12493_);
  nor (_07835_, _07802_, _07785_);
  nor (_07836_, _07835_, _07803_);
  nor (_07837_, _07836_, _06402_);
  nor (_07838_, _07837_, _06512_);
  nor (_07839_, _07838_, _07741_);
  nor (_07840_, _07839_, _07784_);
  nand (_05589_, _07840_, _12493_);
  nor (_07841_, _07803_, _07778_);
  nor (_07842_, _07841_, _07804_);
  nor (_07843_, _07842_, _06402_);
  nor (_07844_, _07843_, _06459_);
  nor (_07845_, _07844_, _07741_);
  nor (_07846_, _07845_, _07777_);
  nor (_05590_, _07846_, rst);
  nor (_07847_, _07804_, _07770_);
  nor (_07848_, _07847_, _07805_);
  nor (_07849_, _07848_, _06402_);
  nor (_07850_, _07849_, _06478_);
  nor (_07851_, _07850_, _07741_);
  nor (_07852_, _07851_, _07769_);
  nor (_05591_, _07852_, rst);
  nor (_07853_, _07805_, _07763_);
  nor (_07854_, _07853_, _07806_);
  nor (_07855_, _07854_, _06402_);
  nor (_07856_, _07855_, _06427_);
  nor (_07857_, _07856_, _07741_);
  nor (_07858_, _07857_, _07762_);
  nor (_05592_, _07858_, rst);
  nor (_07859_, _07806_, _07756_);
  nor (_07860_, _07859_, _07807_);
  nor (_07861_, _07860_, _06402_);
  nor (_07862_, _07861_, _06406_);
  nor (_07863_, _07862_, _07741_);
  nor (_07864_, _07863_, _07755_);
  nor (_05593_, _07864_, rst);
  and (_07865_, _07740_, _07073_);
  nand (_07866_, _07865_, _07738_);
  nor (_07867_, _07866_, _06770_);
  and (_07868_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05610_);
  and (_07869_, _07868_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_07870_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_07871_, _07870_, _07869_);
  or (_07872_, _07871_, _07867_);
  not (_07873_, _07869_);
  nor (_07874_, _06746_, _05684_);
  nor (_07875_, _06806_, _05795_);
  and (_07876_, _06625_, _05698_);
  not (_07877_, _07876_);
  nor (_07878_, _05865_, _06587_);
  and (_07879_, _07878_, _06693_);
  and (_07880_, _07879_, _05726_);
  and (_07881_, _07880_, _06563_);
  and (_07882_, _07881_, _06630_);
  nor (_07883_, _07882_, _06695_);
  and (_07884_, _06625_, _05750_);
  nor (_07885_, _07884_, _07883_);
  and (_07886_, _07885_, _07877_);
  and (_07887_, _06701_, _05865_);
  and (_07888_, _05712_, _05763_);
  nor (_07889_, _05726_, _05777_);
  and (_07890_, _07889_, _07888_);
  and (_07891_, _07890_, _07887_);
  and (_07892_, _05698_, _05750_);
  and (_07893_, _07892_, _07891_);
  nor (_07894_, _07893_, _06625_);
  not (_07895_, _07894_);
  and (_07896_, _07895_, _07886_);
  and (_07897_, _06625_, _05743_);
  nor (_07898_, _07897_, _07247_);
  and (_07899_, _07898_, _07896_);
  nor (_07900_, _07899_, _06708_);
  and (_07901_, _07899_, _06708_);
  nor (_07902_, _07901_, _07900_);
  and (_07903_, _07902_, _06686_);
  and (_07904_, _06625_, _06708_);
  nor (_07905_, _07904_, _06792_);
  nor (_07906_, _07905_, _06713_);
  or (_07907_, _07906_, _07903_);
  or (_07908_, _07907_, _07875_);
  and (_07909_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_07910_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_07911_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_07912_, _07911_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07913_, _07912_, _07910_);
  nor (_07914_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_07915_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_07916_, _07915_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07917_, _07916_, _07914_);
  nor (_07918_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_07919_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_07920_, _07919_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07921_, _07920_, _07918_);
  not (_07922_, _07921_);
  nor (_07923_, _07922_, _06783_);
  nor (_07924_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_07925_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_07926_, _07925_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07927_, _07926_, _07924_);
  and (_07928_, _07927_, _07923_);
  nor (_07929_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_07930_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_07931_, _07930_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07932_, _07931_, _07929_);
  and (_07933_, _07932_, _07928_);
  and (_07934_, _07933_, _07917_);
  nor (_07935_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_07936_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_07937_, _07936_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07938_, _07937_, _07935_);
  and (_07939_, _07938_, _07934_);
  and (_07940_, _07939_, _07913_);
  nor (_07941_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_07942_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_07943_, _07942_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07944_, _07943_, _07941_);
  and (_07945_, _07944_, _07940_);
  nor (_07946_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_07947_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_07948_, _07947_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07949_, _07948_, _07946_);
  nor (_07950_, _07949_, _07945_);
  and (_07951_, _07949_, _07945_);
  or (_07952_, _07951_, _07950_);
  nor (_07953_, _07952_, _06682_);
  and (_07954_, _06082_, _05616_);
  or (_07955_, _07954_, _07953_);
  or (_07956_, _07955_, _07909_);
  or (_07957_, _07956_, _07908_);
  or (_07958_, _07957_, _07874_);
  or (_07959_, _07958_, _07873_);
  and (_07960_, _07959_, _12493_);
  and (_05594_, _07960_, _07872_);
  and (_07961_, _07740_, _07014_);
  and (_07962_, _07961_, _07738_);
  nor (_07963_, _07962_, _07869_);
  not (_07964_, _07963_);
  nand (_07965_, _07964_, _06770_);
  not (_07966_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_07967_, _07963_, _07966_);
  and (_07968_, _07967_, _12493_);
  and (_05595_, _07968_, _07965_);
  nor (_07969_, _07866_, _06877_);
  and (_07970_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_07971_, _07970_, _07869_);
  or (_07972_, _07971_, _07969_);
  and (_07973_, _07922_, _06783_);
  nor (_07974_, _07973_, _07923_);
  and (_07975_, _07974_, _06681_);
  nand (_07976_, _06336_, _06112_);
  nor (_07977_, _06792_, _06711_);
  not (_07978_, _07977_);
  nor (_07979_, _07978_, _06703_);
  nor (_07980_, _07979_, _05777_);
  and (_07981_, _07979_, _05777_);
  nor (_07982_, _07981_, _07980_);
  and (_07983_, _07982_, _06686_);
  and (_07984_, _06745_, _05777_);
  and (_07985_, _06057_, _05616_);
  nor (_07986_, _06806_, _05667_);
  nor (_07987_, _06713_, _05943_);
  or (_07988_, _07987_, _07986_);
  or (_07989_, _07988_, _07985_);
  nor (_07990_, _07989_, _07984_);
  not (_07991_, _07990_);
  nor (_07992_, _07991_, _07983_);
  nand (_07993_, _07992_, _07976_);
  or (_07994_, _07993_, _07975_);
  or (_07995_, _07994_, _07873_);
  and (_07996_, _07995_, _12493_);
  and (_05596_, _07996_, _07972_);
  nor (_07997_, _07866_, _06939_);
  and (_07998_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_07999_, _07998_, _07869_);
  or (_08000_, _07999_, _07997_);
  nor (_08001_, _07927_, _07923_);
  nor (_08002_, _08001_, _07928_);
  and (_08003_, _08002_, _06681_);
  not (_08004_, _08003_);
  and (_08005_, _06236_, _06112_);
  not (_08006_, _08005_);
  and (_08007_, _06745_, _05726_);
  and (_08008_, _07879_, _06625_);
  and (_08009_, _07887_, _06587_);
  and (_08010_, _08009_, _06695_);
  nor (_08011_, _08010_, _08008_);
  nor (_08012_, _08011_, _06139_);
  and (_08013_, _08011_, _06139_);
  or (_08014_, _08013_, _06963_);
  nor (_08015_, _08014_, _08012_);
  and (_08016_, _06059_, _05616_);
  nor (_08017_, _06806_, _05813_);
  and (_08018_, _06712_, _05892_);
  or (_08019_, _08018_, _08017_);
  or (_08020_, _08019_, _08016_);
  or (_08021_, _08020_, _08015_);
  nor (_08022_, _08021_, _08007_);
  and (_08023_, _08022_, _08006_);
  and (_08024_, _08023_, _08004_);
  nand (_08025_, _08024_, _07869_);
  and (_08026_, _08025_, _12493_);
  and (_05597_, _08026_, _08000_);
  nor (_08027_, _07866_, _07000_);
  and (_08028_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_08029_, _08028_, _07869_);
  or (_08030_, _08029_, _08027_);
  nor (_08031_, _07932_, _07928_);
  nor (_08032_, _08031_, _07933_);
  and (_08033_, _08032_, _06681_);
  not (_08034_, _08033_);
  and (_08035_, _08009_, _06139_);
  and (_08036_, _08035_, _06695_);
  and (_08037_, _07880_, _06625_);
  nor (_08038_, _08037_, _08036_);
  and (_08039_, _08038_, _05763_);
  nor (_08040_, _08038_, _05763_);
  nor (_08041_, _08040_, _08039_);
  and (_08042_, _08041_, _06686_);
  and (_08043_, _06061_, _05616_);
  and (_08044_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_08045_, _06806_, _05834_);
  and (_08046_, _06712_, _05907_);
  nor (_08047_, _06746_, _05763_);
  or (_08048_, _08047_, _08046_);
  or (_08049_, _08048_, _08045_);
  nor (_08050_, _08049_, _08044_);
  not (_08051_, _08050_);
  nor (_08052_, _08051_, _08043_);
  not (_08053_, _08052_);
  nor (_08054_, _08053_, _08042_);
  and (_08055_, _08054_, _08034_);
  nand (_08056_, _08055_, _07869_);
  and (_08057_, _08056_, _12493_);
  and (_05598_, _08057_, _08030_);
  not (_08058_, _07065_);
  nor (_08059_, _07866_, _08058_);
  and (_08060_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_08061_, _08060_, _07869_);
  or (_08062_, _08061_, _08059_);
  nor (_08063_, _07933_, _07917_);
  nor (_08064_, _08063_, _07934_);
  and (_08065_, _08064_, _06681_);
  not (_08066_, _08065_);
  nor (_08067_, _07881_, _06630_);
  not (_08068_, _08067_);
  and (_08069_, _08068_, _07883_);
  and (_08070_, _08035_, _05763_);
  nor (_08071_, _08070_, _05712_);
  nor (_08072_, _08071_, _07891_);
  nor (_08073_, _08072_, _06625_);
  nor (_08074_, _08073_, _08069_);
  nor (_08075_, _08074_, _06963_);
  nor (_08076_, _06746_, _05712_);
  or (_08077_, _08076_, _06807_);
  nor (_08078_, _08077_, _08075_);
  and (_08079_, _06064_, _05616_);
  nor (_08080_, _06713_, _05795_);
  and (_08081_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_08082_, _08081_, _08080_);
  nor (_08083_, _08082_, _08079_);
  and (_08084_, _08083_, _08078_);
  and (_08085_, _08084_, _08066_);
  nand (_08086_, _08085_, _07869_);
  and (_08087_, _08086_, _12493_);
  and (_05599_, _08087_, _08062_);
  nor (_08088_, _07866_, _07134_);
  and (_08089_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_08090_, _08089_, _07869_);
  or (_08091_, _08090_, _08088_);
  nor (_08092_, _07938_, _07934_);
  not (_08093_, _08092_);
  nor (_08094_, _07939_, _06682_);
  and (_08095_, _08094_, _08093_);
  not (_08096_, _08095_);
  and (_08097_, _06068_, _05616_);
  nor (_08098_, _07891_, _06625_);
  nor (_08099_, _08098_, _07883_);
  nor (_08100_, _08099_, _06544_);
  and (_08101_, _08099_, _06544_);
  nor (_08102_, _08101_, _08100_);
  and (_08103_, _08102_, _06686_);
  and (_08104_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_08105_, _06625_, _05668_);
  or (_08106_, _08105_, _06713_);
  nor (_08107_, _08106_, _07884_);
  nor (_08108_, _06806_, _05943_);
  nor (_08109_, _06746_, _05750_);
  or (_08110_, _08109_, _08108_);
  or (_08111_, _08110_, _08107_);
  nor (_08112_, _08111_, _08104_);
  not (_08113_, _08112_);
  nor (_08114_, _08113_, _08103_);
  not (_08115_, _08114_);
  nor (_08116_, _08115_, _08097_);
  and (_08117_, _08116_, _08096_);
  nand (_08118_, _08117_, _07869_);
  and (_08119_, _08118_, _12493_);
  and (_05600_, _08119_, _08091_);
  not (_08120_, _07213_);
  nor (_08121_, _07866_, _08120_);
  and (_08122_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_08123_, _08122_, _07869_);
  or (_08124_, _08123_, _08121_);
  nor (_08125_, _07939_, _07913_);
  nor (_08126_, _08125_, _07940_);
  and (_08127_, _08126_, _06681_);
  not (_08128_, _08127_);
  and (_08129_, _06075_, _05616_);
  and (_08130_, _07891_, _05750_);
  nor (_08131_, _08130_, _06625_);
  not (_08132_, _08131_);
  and (_08133_, _08132_, _07885_);
  and (_08134_, _08133_, _05698_);
  nor (_08135_, _08133_, _05698_);
  or (_08136_, _08135_, _08134_);
  and (_08137_, _08136_, _06686_);
  and (_08138_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_08139_, _07250_, _06713_);
  and (_08140_, _08139_, _07877_);
  and (_08141_, _06805_, _05892_);
  nor (_08142_, _06746_, _05698_);
  or (_08143_, _08142_, _08141_);
  or (_08144_, _08143_, _08140_);
  nor (_08145_, _08144_, _08138_);
  not (_08146_, _08145_);
  nor (_08147_, _08146_, _08137_);
  not (_08148_, _08147_);
  nor (_08149_, _08148_, _08129_);
  and (_08150_, _08149_, _08128_);
  nand (_08151_, _08150_, _07869_);
  and (_08152_, _08151_, _12493_);
  and (_05601_, _08152_, _08124_);
  nor (_08153_, _07866_, _07285_);
  and (_08154_, _07866_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_08155_, _08154_, _07869_);
  or (_08156_, _08155_, _08153_);
  nor (_08157_, _07944_, _07940_);
  not (_08158_, _08157_);
  nor (_08159_, _07945_, _06682_);
  and (_08160_, _08159_, _08158_);
  not (_08161_, _08160_);
  and (_08162_, _06079_, _05616_);
  and (_08163_, _07896_, _05743_);
  nor (_08164_, _07896_, _05743_);
  nor (_08165_, _08164_, _08163_);
  nor (_08166_, _08165_, _06963_);
  and (_08167_, _06112_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_08168_, _06625_, _05836_);
  or (_08169_, _08168_, _06713_);
  nor (_08170_, _08169_, _07897_);
  and (_08171_, _06805_, _05907_);
  nor (_08172_, _06746_, _05743_);
  or (_08173_, _08172_, _08171_);
  or (_08174_, _08173_, _08170_);
  nor (_08175_, _08174_, _08167_);
  not (_08176_, _08175_);
  nor (_08177_, _08176_, _08166_);
  not (_08178_, _08177_);
  nor (_08179_, _08178_, _08162_);
  and (_08180_, _08179_, _08161_);
  nand (_08181_, _08180_, _07869_);
  and (_08182_, _08181_, _12493_);
  and (_05602_, _08182_, _08156_);
  nand (_08183_, _07964_, _06877_);
  or (_08184_, _07964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_08185_, _08184_, _12493_);
  and (_05603_, _08185_, _08183_);
  nand (_08186_, _07964_, _06939_);
  or (_08187_, _07964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_08188_, _08187_, _12493_);
  and (_05604_, _08188_, _08186_);
  nand (_08189_, _07964_, _07000_);
  not (_08190_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_08191_, _07963_, _08190_);
  and (_08192_, _08191_, _12493_);
  and (_05605_, _08192_, _08189_);
  or (_08193_, _07963_, _07065_);
  or (_08194_, _07964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_08195_, _08194_, _12493_);
  and (_05606_, _08195_, _08193_);
  nand (_08196_, _07964_, _07134_);
  or (_08197_, _07964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_08198_, _08197_, _12493_);
  and (_05607_, _08198_, _08196_);
  or (_08199_, _07963_, _07213_);
  or (_08200_, _07964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_08201_, _08200_, _12493_);
  and (_05608_, _08201_, _08199_);
  nand (_08202_, _07964_, _07285_);
  or (_08203_, _07964_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_08204_, _08203_, _12493_);
  and (_05609_, _08204_, _08202_);
  nor (_08205_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_08206_, _08205_, _06829_);
  nor (_08207_, _06451_, _06423_);
  and (_08208_, _06485_, _06435_);
  and (_08209_, _08208_, _08207_);
  and (_08210_, _08209_, _06835_);
  and (_08211_, _08205_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_08212_, _08211_, _08210_);
  or (_08213_, _08212_, _08206_);
  and (_08214_, _06777_, _06522_);
  and (_08215_, _08214_, _08209_);
  not (_08216_, _08215_);
  nor (_08217_, _07293_, _06829_);
  not (_08218_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_08219_, _06832_, _08218_);
  nand (_08220_, _08219_, _08210_);
  or (_08221_, _08220_, _08217_);
  and (_08222_, _08221_, _08216_);
  and (_08223_, _08222_, _08213_);
  nor (_08224_, _08216_, _07818_);
  or (_08225_, _08224_, _08223_);
  and (_05620_, _08225_, _12493_);
  nand (_08226_, _08215_, _07790_);
  not (_08227_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_08228_, _08210_, _06947_);
  nor (_08229_, _08228_, _08227_);
  or (_08230_, _08229_, _08215_);
  and (_08231_, _08228_, _06885_);
  or (_08232_, _08231_, _08230_);
  and (_08233_, _08232_, _08226_);
  and (_06067_, _08233_, _12493_);
  or (_08234_, _06090_, _06085_);
  or (_08235_, _08234_, _06096_);
  or (_08236_, _08235_, _06099_);
  or (_08237_, _08236_, _06102_);
  or (_08238_, _08237_, _06105_);
  or (_08239_, _08238_, _06107_);
  and (_08240_, _08239_, _05616_);
  and (_08241_, _06786_, _06639_);
  not (_08242_, _06639_);
  and (_08243_, _06787_, _08242_);
  or (_08244_, _08243_, _08241_);
  and (_08245_, _08244_, _06528_);
  not (_08246_, _06530_);
  nand (_08247_, _06676_, _08246_);
  or (_08248_, _06676_, _06531_);
  and (_08249_, _06681_, _08248_);
  and (_08250_, _08249_, _08247_);
  and (_08251_, _07892_, _06221_);
  and (_08252_, _07890_, _06112_);
  nand (_08253_, _08252_, _08251_);
  nand (_08254_, _08253_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_08255_, _08254_, _08250_);
  nor (_08256_, _08255_, _08245_);
  nand (_08257_, _08256_, _06525_);
  or (_08258_, _08257_, _08240_);
  nor (_08259_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_08260_, _08259_, _08210_);
  and (_08261_, _08260_, _08258_);
  not (_08262_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_08263_, _07014_, _08262_);
  or (_08264_, _08263_, _07015_);
  and (_08265_, _08264_, _08210_);
  or (_08266_, _08265_, _08215_);
  or (_08267_, _08266_, _08261_);
  nand (_08268_, _08215_, _07783_);
  and (_08269_, _08268_, _08267_);
  and (_06069_, _08269_, _12493_);
  and (_08270_, _08210_, _07073_);
  nand (_08271_, _08270_, _06829_);
  or (_08272_, _08270_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_08273_, _08272_, _08216_);
  and (_08274_, _08273_, _08271_);
  nor (_08275_, _08216_, _07776_);
  or (_08276_, _08275_, _08274_);
  and (_06070_, _08276_, _12493_);
  and (_08277_, _07145_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_08278_, _08277_, _07150_);
  and (_08279_, _08278_, _08210_);
  nor (_08280_, _08216_, _07768_);
  not (_08281_, _08210_);
  or (_08282_, _08281_, _07146_);
  not (_08283_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_08284_, _08215_, _08283_);
  and (_08285_, _08284_, _08282_);
  or (_08286_, _08285_, _08280_);
  or (_08287_, _08286_, _08279_);
  and (_06072_, _08287_, _12493_);
  nand (_08288_, _08215_, _07761_);
  and (_08289_, _07228_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_08290_, _08289_, _07227_);
  and (_08291_, _08290_, _08210_);
  or (_08292_, _08281_, _07221_);
  and (_08293_, _08292_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_08294_, _08293_, _08215_);
  or (_08295_, _08294_, _08291_);
  and (_08296_, _08295_, _08288_);
  and (_06074_, _08296_, _12493_);
  or (_08297_, _07296_, _07055_);
  nand (_08298_, _08297_, _08210_);
  or (_08299_, _08298_, _07298_);
  and (_08300_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_08301_, _06681_, _06664_);
  and (_08302_, _06635_, _06528_);
  or (_08303_, _08302_, _08301_);
  and (_08304_, _08303_, _08300_);
  nand (_08305_, _08300_, _06746_);
  and (_08306_, _08305_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_08307_, _08306_, _08210_);
  or (_08308_, _08307_, _08304_);
  and (_08309_, _08308_, _08216_);
  and (_08310_, _08309_, _08299_);
  nor (_08311_, _08216_, _07754_);
  or (_08312_, _08311_, _08310_);
  and (_06076_, _08312_, _12493_);
  not (_08313_, _07868_);
  and (_08314_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05610_);
  and (_08315_, _08314_, _08313_);
  not (_08316_, _06435_);
  and (_08317_, _06522_, _08316_);
  and (_08318_, _06484_, _06468_);
  and (_08319_, _08318_, _06777_);
  and (_08320_, _08319_, _08317_);
  and (_08321_, _08320_, _08207_);
  nor (_08322_, _08321_, _08315_);
  or (_08323_, _08322_, _06770_);
  not (_08324_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_08325_, _07868_, _08324_);
  nand (_08326_, _08318_, _06436_);
  and (_08327_, _06835_, _06452_);
  not (_08328_, _08327_);
  nor (_08329_, _08328_, _08326_);
  and (_08330_, _08329_, _06832_);
  and (_08331_, _08330_, _06829_);
  nor (_08332_, _08330_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_08333_, _08325_);
  and (_08334_, _08333_, _08322_);
  not (_08335_, _08334_);
  nor (_08336_, _08335_, _08332_);
  not (_08337_, _08336_);
  nor (_08338_, _08337_, _08331_);
  nor (_08339_, _08338_, _08325_);
  nand (_08340_, _08339_, _08323_);
  or (_08341_, _08333_, _07958_);
  and (_08342_, _08341_, _08340_);
  and (_06136_, _08342_, _12493_);
  or (_08343_, _08322_, _06877_);
  and (_08344_, _08329_, _06522_);
  and (_08345_, _08344_, _06829_);
  nor (_08346_, _08344_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_08347_, _08346_, _08335_);
  not (_08348_, _08347_);
  nor (_08349_, _08348_, _08345_);
  nor (_08350_, _08349_, _08325_);
  nand (_08351_, _08350_, _08343_);
  or (_08352_, _08333_, _07994_);
  and (_08353_, _08352_, _08351_);
  and (_06308_, _08353_, _12493_);
  or (_08354_, _08322_, _06939_);
  and (_08355_, _08329_, _06947_);
  and (_08356_, _08355_, _06829_);
  nor (_08357_, _08355_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_08358_, _08357_, _08335_);
  not (_08359_, _08358_);
  nor (_08360_, _08359_, _08356_);
  nor (_08361_, _08360_, _08325_);
  nand (_08362_, _08361_, _08354_);
  and (_08363_, _08325_, _08024_);
  not (_08364_, _08363_);
  and (_08365_, _08364_, _08362_);
  and (_06310_, _08365_, _12493_);
  or (_08366_, _08322_, _07000_);
  and (_08367_, _08329_, _07014_);
  and (_08368_, _08367_, _06829_);
  nor (_08369_, _08367_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_08370_, _08369_, _08335_);
  not (_08371_, _08370_);
  nor (_08372_, _08371_, _08368_);
  nor (_08373_, _08372_, _08325_);
  nand (_08374_, _08373_, _08366_);
  and (_08375_, _08325_, _08055_);
  not (_08376_, _08375_);
  and (_08377_, _08376_, _08374_);
  and (_06312_, _08377_, _12493_);
  nor (_08378_, _08333_, _08085_);
  not (_08379_, _08378_);
  or (_08380_, _08322_, _07065_);
  not (_08381_, _08322_);
  and (_08382_, _08318_, _06452_);
  and (_08383_, _06835_, _06436_);
  and (_08384_, _08383_, _08382_);
  nor (_08385_, _08384_, _05709_);
  nor (_08386_, _08385_, _08381_);
  not (_08387_, _08384_);
  nor (_08388_, _07073_, _05709_);
  nor (_08389_, _08388_, _07075_);
  or (_08390_, _08389_, _08387_);
  and (_08391_, _08390_, _08386_);
  nor (_08392_, _08391_, _08325_);
  nand (_08393_, _08392_, _08380_);
  nand (_08394_, _08393_, _08379_);
  and (_06314_, _08394_, _12493_);
  or (_08395_, _08322_, _07134_);
  and (_08396_, _08329_, _07144_);
  and (_08397_, _08396_, _06829_);
  nor (_08398_, _08396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_08399_, _08398_, _08335_);
  not (_08400_, _08399_);
  nor (_08401_, _08400_, _08397_);
  nor (_08402_, _08401_, _08325_);
  nand (_08403_, _08402_, _08395_);
  and (_08404_, _08325_, _08117_);
  not (_08405_, _08404_);
  and (_08406_, _08405_, _08403_);
  and (_06316_, _08406_, _12493_);
  nor (_08407_, _08333_, _08150_);
  not (_08408_, _08407_);
  or (_08409_, _08322_, _07213_);
  nor (_08410_, _07225_, _05695_);
  nor (_08411_, _08410_, _07227_);
  nor (_08412_, _08411_, _08387_);
  nor (_08413_, _08384_, _05695_);
  nor (_08414_, _08413_, _08381_);
  not (_08415_, _08414_);
  nor (_08416_, _08415_, _08412_);
  nor (_08417_, _08416_, _08325_);
  nand (_08418_, _08417_, _08409_);
  nand (_08419_, _08418_, _08408_);
  and (_06318_, _08419_, _12493_);
  or (_08420_, _08322_, _07285_);
  and (_08421_, _08329_, _07296_);
  and (_08422_, _08421_, _06829_);
  nor (_08423_, _08421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_08424_, _08423_, _08335_);
  not (_08425_, _08424_);
  nor (_08426_, _08425_, _08422_);
  nor (_08427_, _08426_, _08325_);
  nand (_08428_, _08427_, _08420_);
  and (_08429_, _08325_, _08180_);
  not (_08430_, _08429_);
  and (_08431_, _08430_, _08428_);
  and (_06320_, _08431_, _12493_);
  and (_08432_, _07738_, _06468_);
  and (_08433_, _08432_, _06832_);
  nand (_08434_, _08433_, _06829_);
  or (_08435_, _08433_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_08436_, _08435_, _06835_);
  and (_08437_, _08436_, _08434_);
  and (_08438_, _08432_, _06522_);
  nand (_08439_, _08438_, _07818_);
  or (_08440_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_08441_, _08440_, _06777_);
  and (_08442_, _08441_, _08439_);
  not (_08443_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_08444_, _06776_, _08443_);
  or (_08445_, _08444_, rst);
  or (_08446_, _08445_, _08442_);
  or (_07330_, _08446_, _08437_);
  and (_08447_, _07735_, _06486_);
  and (_08448_, _08447_, _06832_);
  nand (_08449_, _08448_, _06829_);
  or (_08450_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_08451_, _08450_, _06835_);
  and (_08452_, _08451_, _08449_);
  not (_08453_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_08454_, _08447_, _06522_);
  nor (_08455_, _08454_, _08453_);
  not (_08456_, _08454_);
  nor (_08457_, _08456_, _07818_);
  or (_08458_, _08457_, _08455_);
  and (_08459_, _08458_, _06777_);
  nor (_08460_, _06776_, _08453_);
  or (_08461_, _08460_, rst);
  or (_08462_, _08461_, _08459_);
  or (_07333_, _08462_, _08452_);
  and (_08463_, _08316_, _06423_);
  and (_08464_, _08463_, _08382_);
  and (_08465_, _08464_, _06832_);
  nand (_08466_, _08465_, _06829_);
  or (_08467_, _08465_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_08468_, _08467_, _06835_);
  and (_08469_, _08468_, _08466_);
  and (_08470_, _08464_, _06522_);
  not (_08471_, _08470_);
  nor (_08472_, _08471_, _07818_);
  not (_08473_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_08474_, _08470_, _08473_);
  or (_08475_, _08474_, _08472_);
  and (_08476_, _08475_, _06777_);
  nor (_08477_, _06776_, _08473_);
  or (_08478_, _08477_, rst);
  or (_08479_, _08478_, _08476_);
  or (_07336_, _08479_, _08469_);
  and (_08480_, _08463_, _06486_);
  not (_08481_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_08482_, _06832_, _08481_);
  or (_08483_, _08482_, _08217_);
  and (_08484_, _08483_, _08480_);
  nor (_08485_, _08480_, _08481_);
  or (_08486_, _08485_, _08484_);
  and (_08487_, _08486_, _06835_);
  and (_08488_, _06522_, _06485_);
  and (_08489_, _08488_, _06452_);
  and (_08490_, _08463_, _08489_);
  nor (_08491_, _08490_, _08481_);
  not (_08492_, _08490_);
  nor (_08493_, _08492_, _07818_);
  or (_08494_, _08493_, _08491_);
  and (_08495_, _08494_, _06777_);
  nor (_08496_, _06776_, _08481_);
  or (_08497_, _08496_, rst);
  or (_08498_, _08497_, _08495_);
  or (_07339_, _08498_, _08487_);
  or (_08499_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_08500_, _08438_, _06829_);
  and (_08501_, _08500_, _06835_);
  nand (_08502_, _08438_, _07797_);
  and (_08503_, _08502_, _06777_);
  or (_08504_, _08503_, _08501_);
  and (_08505_, _08504_, _08499_);
  not (_08506_, _06776_);
  and (_08507_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_08508_, _08507_, rst);
  or (_09974_, _08508_, _08505_);
  and (_08509_, _08432_, _06947_);
  nand (_08510_, _08509_, _06829_);
  or (_08511_, _08509_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_08512_, _08511_, _06835_);
  and (_08513_, _08512_, _08510_);
  nand (_08514_, _08438_, _07790_);
  or (_08515_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_08516_, _08515_, _06777_);
  and (_08517_, _08516_, _08514_);
  and (_08518_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_08519_, _08518_, rst);
  or (_08520_, _08519_, _08517_);
  or (_09976_, _08520_, _08513_);
  not (_08521_, _07077_);
  nand (_08522_, _08432_, _08521_);
  and (_08523_, _08522_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_08524_, _06521_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_08525_, _08524_, _07015_);
  and (_08526_, _08525_, _08432_);
  or (_08527_, _08526_, _08523_);
  and (_08528_, _08527_, _06835_);
  nand (_08529_, _08438_, _07783_);
  or (_08530_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_08531_, _08530_, _06777_);
  and (_08532_, _08531_, _08529_);
  not (_08533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_08534_, _06776_, _08533_);
  or (_08535_, _08534_, rst);
  or (_08536_, _08535_, _08532_);
  or (_09978_, _08536_, _08528_);
  nand (_08537_, _08432_, _06520_);
  and (_08538_, _08537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_08539_, _08521_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_08540_, _08539_, _07075_);
  and (_08541_, _08540_, _08432_);
  or (_08542_, _08541_, _08538_);
  and (_08543_, _08542_, _06835_);
  nand (_08544_, _08438_, _07776_);
  or (_08545_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_08546_, _08545_, _06777_);
  and (_08547_, _08546_, _08544_);
  and (_08548_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_08549_, _08548_, rst);
  or (_08550_, _08549_, _08547_);
  or (_09980_, _08550_, _08543_);
  and (_08551_, _08432_, _07144_);
  nand (_08552_, _08551_, _06829_);
  or (_08553_, _08551_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_08554_, _08553_, _06835_);
  and (_08555_, _08554_, _08552_);
  nand (_08556_, _08438_, _07768_);
  or (_08557_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_08558_, _08557_, _06777_);
  and (_08559_, _08558_, _08556_);
  and (_08560_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_08561_, _08560_, rst);
  or (_08562_, _08561_, _08559_);
  or (_09982_, _08562_, _08555_);
  and (_08563_, _08432_, _07225_);
  nand (_08564_, _08563_, _06829_);
  or (_08565_, _08563_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_08566_, _08565_, _06835_);
  and (_08567_, _08566_, _08564_);
  nand (_08568_, _08438_, _07761_);
  or (_08569_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_08570_, _08569_, _06777_);
  and (_08571_, _08570_, _08568_);
  and (_08572_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_08573_, _08572_, rst);
  or (_08574_, _08573_, _08571_);
  or (_09984_, _08574_, _08567_);
  nand (_08575_, _08432_, _07293_);
  and (_08576_, _08575_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_08577_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_08578_, _06831_, _08577_);
  or (_08579_, _08578_, _07298_);
  and (_08580_, _08579_, _08432_);
  or (_08581_, _08580_, _08576_);
  and (_08582_, _08581_, _06835_);
  nand (_08583_, _08438_, _07754_);
  or (_08584_, _08438_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_08585_, _08584_, _06777_);
  and (_08586_, _08585_, _08583_);
  nor (_08587_, _06776_, _08577_);
  or (_08588_, _08587_, rst);
  or (_08589_, _08588_, _08586_);
  or (_09986_, _08589_, _08582_);
  nand (_08590_, _08454_, _06829_);
  or (_08591_, _08454_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_08592_, _08591_, _06835_);
  and (_08593_, _08592_, _08590_);
  and (_08594_, _08456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_08595_, _08454_, _07798_);
  or (_08596_, _08595_, _08594_);
  and (_08597_, _08596_, _06777_);
  and (_08598_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_08599_, _08598_, rst);
  or (_08600_, _08599_, _08597_);
  or (_09988_, _08600_, _08593_);
  and (_08601_, _08447_, _06947_);
  nand (_08602_, _08601_, _06829_);
  or (_08603_, _08601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_08604_, _08603_, _06835_);
  and (_08605_, _08604_, _08602_);
  and (_08606_, _08456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_08607_, _08456_, _07790_);
  or (_08608_, _08607_, _08606_);
  and (_08609_, _08608_, _06777_);
  and (_08610_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_08611_, _08610_, rst);
  or (_08612_, _08611_, _08609_);
  or (_09990_, _08612_, _08605_);
  and (_08613_, _08447_, _07014_);
  nand (_08614_, _08613_, _06829_);
  or (_08615_, _08613_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_08616_, _08615_, _06835_);
  and (_08617_, _08616_, _08614_);
  not (_08618_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_08619_, _08454_, _08618_);
  nor (_08620_, _08456_, _07783_);
  or (_08621_, _08620_, _08619_);
  and (_08622_, _08621_, _06777_);
  nor (_08623_, _06776_, _08618_);
  or (_08624_, _08623_, rst);
  or (_08625_, _08624_, _08622_);
  or (_09992_, _08625_, _08617_);
  and (_08626_, _08447_, _07073_);
  nand (_08627_, _08626_, _06829_);
  or (_08628_, _08626_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_08629_, _08628_, _06835_);
  and (_08630_, _08629_, _08627_);
  and (_08631_, _08456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_08632_, _08456_, _07776_);
  or (_08633_, _08632_, _08631_);
  and (_08634_, _08633_, _06777_);
  and (_08635_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_08636_, _08635_, rst);
  or (_08637_, _08636_, _08634_);
  or (_09994_, _08637_, _08630_);
  and (_08638_, _08447_, _07144_);
  nand (_08639_, _08638_, _06829_);
  or (_08640_, _08638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_08641_, _08640_, _06835_);
  and (_08642_, _08641_, _08639_);
  and (_08643_, _08456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_08644_, _08456_, _07768_);
  or (_08645_, _08644_, _08643_);
  and (_08646_, _08645_, _06777_);
  and (_08647_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_08648_, _08647_, rst);
  or (_08649_, _08648_, _08646_);
  or (_09995_, _08649_, _08642_);
  and (_08650_, _08447_, _07225_);
  nand (_08651_, _08650_, _06829_);
  or (_08652_, _08650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_08653_, _08652_, _06835_);
  and (_08654_, _08653_, _08651_);
  and (_08655_, _08456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_08656_, _08456_, _07761_);
  or (_08657_, _08656_, _08655_);
  and (_08658_, _08657_, _06777_);
  and (_08659_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_08660_, _08659_, rst);
  or (_08661_, _08660_, _08658_);
  or (_09997_, _08661_, _08654_);
  and (_08662_, _08447_, _07296_);
  nand (_08663_, _08662_, _06829_);
  or (_08664_, _08662_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_08665_, _08664_, _06835_);
  and (_08666_, _08665_, _08663_);
  and (_08667_, _08456_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_08668_, _08456_, _07754_);
  or (_08669_, _08668_, _08667_);
  and (_08670_, _08669_, _06777_);
  and (_08671_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_08672_, _08671_, rst);
  or (_08673_, _08672_, _08670_);
  or (_09999_, _08673_, _08666_);
  nand (_08674_, _08470_, _06829_);
  or (_08675_, _08470_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_08676_, _08675_, _06835_);
  and (_08677_, _08676_, _08674_);
  and (_08678_, _08470_, _07798_);
  and (_08679_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_08680_, _08679_, _08678_);
  and (_08681_, _08680_, _06777_);
  and (_08682_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_08683_, _08682_, rst);
  or (_08684_, _08683_, _08681_);
  or (_10001_, _08684_, _08677_);
  and (_08685_, _08464_, _06947_);
  nand (_08686_, _08685_, _06829_);
  or (_08687_, _08685_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_08688_, _08687_, _06835_);
  and (_08689_, _08688_, _08686_);
  nor (_08690_, _08471_, _07790_);
  and (_08691_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_08692_, _08691_, _08690_);
  and (_08693_, _08692_, _06777_);
  and (_08694_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_08695_, _08694_, rst);
  or (_08696_, _08695_, _08693_);
  or (_10003_, _08696_, _08689_);
  and (_08697_, _08464_, _07014_);
  nand (_08698_, _08697_, _06829_);
  or (_08699_, _08697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_08700_, _08699_, _06835_);
  and (_08701_, _08700_, _08698_);
  nor (_08702_, _08471_, _07783_);
  not (_08703_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_08704_, _08470_, _08703_);
  or (_08705_, _08704_, _08702_);
  and (_08706_, _08705_, _06777_);
  nor (_08707_, _06776_, _08703_);
  or (_08708_, _08707_, rst);
  or (_08709_, _08708_, _08706_);
  or (_10005_, _08709_, _08701_);
  and (_08710_, _08464_, _07073_);
  nand (_08711_, _08710_, _06829_);
  or (_08712_, _08710_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_08713_, _08712_, _06835_);
  and (_08714_, _08713_, _08711_);
  nor (_08715_, _08471_, _07776_);
  and (_08716_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_08717_, _08716_, _08715_);
  and (_08718_, _08717_, _06777_);
  and (_08719_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_08720_, _08719_, rst);
  or (_08721_, _08720_, _08718_);
  or (_10007_, _08721_, _08714_);
  and (_08722_, _08464_, _07144_);
  nand (_08723_, _08722_, _06829_);
  or (_08724_, _08722_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_08725_, _08724_, _06835_);
  and (_08726_, _08725_, _08723_);
  nor (_08727_, _08471_, _07768_);
  and (_08728_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_08729_, _08728_, _08727_);
  and (_08730_, _08729_, _06777_);
  and (_08731_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_08732_, _08731_, rst);
  or (_08733_, _08732_, _08730_);
  or (_10009_, _08733_, _08726_);
  and (_08734_, _08464_, _07225_);
  nand (_08735_, _08734_, _06829_);
  or (_08736_, _08734_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_08737_, _08736_, _06835_);
  and (_08738_, _08737_, _08735_);
  nor (_08739_, _08471_, _07761_);
  and (_08740_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_08741_, _08740_, _08739_);
  and (_08742_, _08741_, _06777_);
  and (_08743_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_08744_, _08743_, rst);
  or (_08745_, _08744_, _08742_);
  or (_10011_, _08745_, _08738_);
  and (_08746_, _08464_, _07296_);
  nand (_08747_, _08746_, _06829_);
  or (_08748_, _08746_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_08749_, _08748_, _06835_);
  and (_08750_, _08749_, _08747_);
  nor (_08751_, _08471_, _07754_);
  and (_08752_, _08471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_08753_, _08752_, _08751_);
  and (_08754_, _08753_, _06777_);
  and (_08755_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_08756_, _08755_, rst);
  or (_08757_, _08756_, _08754_);
  or (_10013_, _08757_, _08750_);
  nand (_08758_, _06829_, _06522_);
  or (_08759_, _06522_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_08760_, _08759_, _08480_);
  and (_08761_, _08760_, _08758_);
  not (_08762_, _08480_);
  and (_08763_, _08762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_08764_, _08763_, _08761_);
  and (_08765_, _08764_, _06835_);
  and (_08766_, _08492_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_08767_, _08492_, _07797_);
  or (_08768_, _08767_, _08766_);
  and (_08769_, _08768_, _06777_);
  and (_08770_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_08771_, _08770_, rst);
  or (_08772_, _08771_, _08769_);
  or (_10015_, _08772_, _08765_);
  nand (_08773_, _06947_, _06829_);
  or (_08774_, _06947_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_08775_, _08774_, _08480_);
  and (_08776_, _08775_, _08773_);
  and (_08777_, _08762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_08778_, _08777_, _08776_);
  and (_08779_, _08778_, _06835_);
  and (_08780_, _08492_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_08781_, _08492_, _07790_);
  or (_08782_, _08781_, _08780_);
  and (_08783_, _08782_, _06777_);
  and (_08784_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_08785_, _08784_, rst);
  or (_08786_, _08785_, _08783_);
  or (_10017_, _08786_, _08779_);
  not (_08787_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_08788_, _07014_, _08787_);
  or (_08789_, _08788_, _07015_);
  and (_08790_, _08789_, _08480_);
  nor (_08791_, _08480_, _08787_);
  or (_08792_, _08791_, _08790_);
  and (_08793_, _08792_, _06835_);
  nor (_08794_, _08490_, _08787_);
  nor (_08795_, _08492_, _07783_);
  or (_08796_, _08795_, _08794_);
  and (_08797_, _08796_, _06777_);
  nor (_08798_, _06776_, _08787_);
  or (_08799_, _08798_, rst);
  or (_08800_, _08799_, _08797_);
  or (_10019_, _08800_, _08793_);
  and (_08801_, _07074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_08802_, _08801_, _07075_);
  and (_08803_, _08802_, _08480_);
  and (_08804_, _08762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_08805_, _08804_, _08803_);
  and (_08806_, _08805_, _06835_);
  and (_08807_, _08492_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_08808_, _08492_, _07776_);
  or (_08809_, _08808_, _08807_);
  and (_08810_, _08809_, _06777_);
  and (_08811_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_08812_, _08811_, rst);
  or (_08813_, _08812_, _08810_);
  or (_10021_, _08813_, _08806_);
  and (_08814_, _07149_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_08815_, _08814_, _07150_);
  and (_08816_, _08815_, _08480_);
  and (_08817_, _08762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_08818_, _08817_, _08816_);
  and (_08819_, _08818_, _06835_);
  and (_08820_, _08492_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_08821_, _08492_, _07768_);
  or (_08822_, _08821_, _08820_);
  and (_08823_, _08822_, _06777_);
  and (_08824_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_08825_, _08824_, rst);
  or (_08826_, _08825_, _08823_);
  or (_10023_, _08826_, _08819_);
  and (_08827_, _07226_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_08828_, _08827_, _07227_);
  and (_08829_, _08828_, _08480_);
  and (_08830_, _08762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_08831_, _08830_, _08829_);
  and (_08832_, _08831_, _06835_);
  and (_08833_, _08492_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_08834_, _08492_, _07761_);
  or (_08835_, _08834_, _08833_);
  and (_08836_, _08835_, _06777_);
  and (_08837_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_08838_, _08837_, rst);
  or (_08839_, _08838_, _08836_);
  or (_10025_, _08839_, _08832_);
  and (_08840_, _07297_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_08841_, _08840_, _07298_);
  and (_08842_, _08841_, _08480_);
  and (_08843_, _08762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_08844_, _08843_, _08842_);
  and (_08845_, _08844_, _06835_);
  and (_08846_, _08492_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_08847_, _08492_, _07754_);
  or (_08848_, _08847_, _08846_);
  and (_08849_, _08848_, _06777_);
  and (_08850_, _08506_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_08851_, _08850_, rst);
  or (_08852_, _08851_, _08849_);
  or (_10027_, _08852_, _08845_);
  and (_08853_, _06451_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_08854_, _08853_, _08316_);
  nor (_08855_, _06520_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_08856_, _08855_, _08854_);
  not (_08857_, _08856_);
  and (_08858_, _07657_, _07616_);
  not (_08859_, _07693_);
  and (_08860_, _08859_, _07658_);
  nor (_08861_, _07683_, _07667_);
  nor (_08862_, _07675_, _07670_);
  and (_08863_, _08862_, _08861_);
  and (_08864_, _07692_, _07680_);
  and (_08865_, _08864_, _08863_);
  and (_08866_, _08865_, _08860_);
  nor (_08867_, _08866_, _07308_);
  nor (_08868_, _08867_, _08858_);
  not (_08869_, _08868_);
  not (_08870_, _07624_);
  and (_08871_, _07718_, _08870_);
  and (_08872_, _08871_, _07733_);
  and (_08873_, _06774_, _06449_);
  not (_08874_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_08875_, _06521_, _08874_);
  and (_08876_, _08875_, _08873_);
  and (_08877_, _07360_, _06830_);
  nor (_08878_, _07360_, _06830_);
  nor (_08879_, _08878_, _08877_);
  and (_08880_, _08879_, _08876_);
  not (_08881_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_08882_, _08215_, _08881_);
  nor (_08883_, _08882_, _08275_);
  and (_08884_, _08883_, _06469_);
  nor (_08885_, _08883_, _06469_);
  nor (_08886_, _08885_, _08884_);
  and (_08887_, _08886_, _08880_);
  not (_08888_, _08887_);
  nor (_08889_, _08888_, _07783_);
  and (_08890_, _08853_, _06423_);
  nor (_08891_, _08853_, _06469_);
  nor (_08892_, _08891_, _08890_);
  nor (_08893_, _08892_, _08883_);
  not (_08894_, _08893_);
  and (_08895_, _08892_, _08883_);
  and (_08896_, _08853_, _06469_);
  nor (_08897_, _06498_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_08898_, _08897_, _08896_);
  and (_08899_, _08898_, _07601_);
  nor (_08900_, _08898_, _07601_);
  nor (_08901_, _08900_, _08899_);
  and (_08902_, _08853_, _07736_);
  nor (_08903_, _06509_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_08904_, _08903_, _08902_);
  and (_08905_, _08904_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_08906_, _08905_, _08856_);
  and (_08907_, _08906_, _08901_);
  not (_08908_, _08907_);
  nor (_08909_, _08908_, _08895_);
  and (_08910_, _08909_, _08894_);
  not (_08911_, _08910_);
  and (_08912_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _06592_);
  nand (_08913_, _08912_, _06600_);
  nor (_08914_, _08913_, _06829_);
  nor (_08915_, _07783_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_08916_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_08917_, _08912_, _06593_);
  nor (_08918_, _08917_, _08916_);
  nand (_08919_, _08912_, _06602_);
  nand (_08920_, _08919_, _08918_);
  and (_08921_, _08920_, _05754_);
  or (_08922_, _08921_, _08915_);
  or (_08923_, _08922_, _08914_);
  or (_08924_, _08923_, _08911_);
  and (_08925_, _08883_, _07360_);
  and (_08926_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_08927_, _08883_, _07601_);
  and (_08928_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_08929_, _08928_, _08926_);
  nor (_08930_, _08883_, _07360_);
  and (_08931_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_08932_, _08883_, _07601_);
  and (_08933_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_08934_, _08933_, _08931_);
  or (_08935_, _08934_, _08929_);
  or (_08936_, _08935_, _08910_);
  and (_08937_, _08936_, _08888_);
  and (_08938_, _08937_, _08924_);
  or (_08939_, _08938_, _08889_);
  and (_08940_, _08939_, _08872_);
  not (_08941_, _08940_);
  and (_08942_, _07733_, _07719_);
  not (_08943_, _07840_);
  and (_08944_, _08943_, _08942_);
  not (_08945_, _08944_);
  and (_08946_, _07733_, _07624_);
  and (_08947_, _08946_, _07718_);
  and (_08948_, _08947_, _07552_);
  nor (_08949_, _07718_, _08870_);
  and (_08950_, _08949_, _07733_);
  not (_08951_, _07312_);
  and (_08952_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_08953_, _07319_, _07312_);
  not (_08954_, _08953_);
  and (_08955_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_08956_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_08957_, _08956_, _08955_);
  and (_08958_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not (_08959_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_08960_, _07324_, _08959_);
  nor (_08961_, _08960_, _08958_);
  and (_08962_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_08963_, _07329_, _07365_);
  nor (_08964_, _08963_, _08962_);
  and (_08965_, _08964_, _08961_);
  and (_08966_, _08965_, _08957_);
  nor (_08967_, _08966_, _08954_);
  nor (_08968_, _08967_, _08952_);
  not (_08969_, _08968_);
  and (_08970_, _08969_, _08950_);
  nor (_08971_, _08970_, _08948_);
  and (_08972_, _08971_, _08945_);
  and (_08973_, _08972_, _08941_);
  nor (_08974_, _08973_, _08869_);
  and (_08975_, _06603_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_08976_, _08975_);
  and (_08977_, _05689_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_08978_, _08977_, _08976_);
  and (_08979_, _08916_, _06603_);
  and (_08980_, _08979_, _06885_);
  nor (_08981_, _07761_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_08982_, _08981_, _08980_);
  or (_08983_, _08982_, _08978_);
  nor (_08984_, _08983_, _08911_);
  and (_08985_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_08986_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_08987_, _08986_, _08985_);
  and (_08988_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_08989_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_08990_, _08989_, _08988_);
  and (_08991_, _08990_, _08987_);
  and (_08992_, _08991_, _08911_);
  or (_08993_, _08992_, _08984_);
  and (_08994_, _08993_, _08888_);
  and (_08995_, _08887_, _07761_);
  nor (_08996_, _08995_, _08994_);
  nand (_08997_, _08996_, _08872_);
  not (_08998_, _08942_);
  nor (_08999_, _07858_, _08998_);
  and (_09000_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_09001_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_09002_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_09003_, _09002_, _09001_);
  and (_09004_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_09005_, _07329_, _07498_);
  nor (_09006_, _09005_, _09004_);
  and (_09007_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not (_09008_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_09009_, _07324_, _09008_);
  nor (_09010_, _09009_, _09007_);
  and (_09011_, _09010_, _09006_);
  and (_09012_, _09011_, _09003_);
  nor (_09013_, _09012_, _08954_);
  nor (_09014_, _09013_, _09000_);
  not (_09015_, _09014_);
  and (_09016_, _09015_, _08950_);
  not (_09017_, _08949_);
  nor (_09018_, _08871_, _07733_);
  and (_09019_, _09018_, _09017_);
  nor (_09020_, _09019_, _09016_);
  not (_09021_, _09020_);
  nor (_09022_, _09021_, _08999_);
  and (_09023_, _09022_, _08997_);
  not (_09024_, _09023_);
  nand (_09025_, _07559_, _07654_);
  and (_09026_, _07710_, _09025_);
  nor (_09027_, _09026_, _07706_);
  not (_09028_, _07690_);
  and (_09029_, _07566_, _07707_);
  and (_09030_, _09029_, _07559_);
  nor (_09031_, _09030_, _07670_);
  and (_09032_, _09031_, _09028_);
  and (_09033_, _09032_, _08859_);
  and (_09034_, _09029_, _07441_);
  not (_09035_, _09034_);
  and (_09036_, _09035_, _09026_);
  and (_09037_, _07524_, _07561_);
  and (_09038_, _07588_, _09037_);
  and (_09039_, _09038_, _07441_);
  nor (_09040_, _09039_, _07677_);
  and (_09041_, _09040_, _07709_);
  and (_09042_, _09041_, _09036_);
  and (_09043_, _09042_, _09033_);
  and (_09044_, _09043_, _08861_);
  nor (_09045_, _09044_, _07308_);
  nor (_09046_, _09045_, _09027_);
  not (_09047_, _06593_);
  and (_09048_, _08916_, _09047_);
  nor (_09049_, _09048_, _08912_);
  not (_09050_, _09049_);
  and (_09051_, _09050_, _05672_);
  and (_09052_, _08916_, _06593_);
  and (_09053_, _09052_, _06885_);
  nor (_09054_, _07818_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_09055_, _09054_, _09053_);
  or (_09056_, _09055_, _09051_);
  nor (_09057_, _09056_, _08911_);
  and (_09058_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_09059_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_09060_, _09059_, _09058_);
  and (_09061_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_09062_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_09063_, _09062_, _09061_);
  and (_09064_, _09063_, _09060_);
  and (_09065_, _09064_, _08911_);
  or (_09066_, _09065_, _09057_);
  and (_09067_, _09066_, _08888_);
  and (_09068_, _08887_, _07818_);
  nor (_09069_, _09068_, _09067_);
  nand (_09070_, _09069_, _08872_);
  not (_09071_, _07733_);
  and (_09072_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_09073_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_09074_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_09075_, _09074_, _09073_);
  and (_09076_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_09077_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_09078_, _07324_, _09077_);
  nor (_09079_, _09078_, _09076_);
  and (_09080_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_09081_, _07329_, _07449_);
  nor (_09082_, _09081_, _09080_);
  and (_09083_, _09082_, _09079_);
  and (_09084_, _09083_, _09075_);
  nor (_09085_, _09084_, _08954_);
  nor (_09086_, _09085_, _09072_);
  not (_09087_, _09086_);
  and (_09088_, _09087_, _08949_);
  nor (_09089_, _09088_, _09071_);
  nand (_09090_, _07820_, _07719_);
  and (_09091_, _09090_, _09089_);
  and (_09092_, _09091_, _09070_);
  not (_09093_, _09092_);
  nor (_09094_, _09093_, _09046_);
  and (_09095_, _09094_, _09024_);
  nor (_09096_, _09095_, _08974_);
  and (_09097_, _09096_, _08857_);
  not (_09098_, _08898_);
  and (_09099_, _08912_, _06596_);
  and (_09100_, _09099_, _06829_);
  not (_09101_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_09102_, _07797_, _09101_);
  nor (_09103_, _05768_, _09101_);
  nor (_09104_, _09103_, _09102_);
  nor (_09105_, _09104_, _09099_);
  nor (_09106_, _09105_, _09100_);
  nor (_09107_, _09106_, _08911_);
  and (_09108_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_09109_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_09110_, _09109_, _09108_);
  and (_09111_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_09112_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_09113_, _09112_, _09111_);
  and (_09114_, _09113_, _09110_);
  and (_09115_, _09114_, _08911_);
  nor (_09116_, _09115_, _09107_);
  nor (_09117_, _09116_, _08887_);
  and (_09118_, _08887_, _07797_);
  nor (_09119_, _09118_, _09117_);
  and (_09120_, _09119_, _08872_);
  not (_09121_, _09120_);
  not (_09122_, _07828_);
  and (_09123_, _09122_, _08942_);
  not (_09124_, _09123_);
  and (_09125_, _08947_, _07601_);
  and (_09126_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_09127_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_09128_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_09129_, _09128_, _09127_);
  not (_09130_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_09131_, _07324_, _09130_);
  nor (_09132_, _07329_, _07320_);
  nor (_09133_, _09132_, _09131_);
  and (_09134_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_09135_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_09136_, _09135_, _09134_);
  and (_09137_, _09136_, _09133_);
  and (_09138_, _09137_, _09129_);
  nor (_09139_, _09138_, _08954_);
  nor (_09140_, _09139_, _09126_);
  not (_09141_, _09140_);
  and (_09142_, _09141_, _08950_);
  nor (_09143_, _09142_, _09125_);
  and (_09144_, _09143_, _09124_);
  and (_09145_, _09144_, _09121_);
  nor (_09146_, _09145_, _08869_);
  not (_09147_, _07776_);
  and (_09148_, _08887_, _09147_);
  and (_09149_, _08917_, _06885_);
  nor (_09150_, _07776_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_09151_, _08912_, _09047_);
  or (_09152_, _09151_, _08916_);
  and (_09153_, _09152_, _05703_);
  or (_09154_, _09153_, _09150_);
  or (_09155_, _09154_, _09149_);
  or (_09156_, _09155_, _08911_);
  and (_09157_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_09158_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_09159_, _09158_, _09157_);
  and (_09160_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_09161_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_09162_, _09161_, _09160_);
  or (_09163_, _09162_, _09159_);
  or (_09164_, _09163_, _08910_);
  and (_09165_, _09164_, _08888_);
  and (_09166_, _09165_, _09156_);
  or (_09167_, _09166_, _09148_);
  and (_09168_, _09167_, _08872_);
  not (_09169_, _09168_);
  not (_09170_, _07846_);
  and (_09171_, _09170_, _08942_);
  not (_09172_, _09171_);
  not (_09173_, _08883_);
  and (_09174_, _08947_, _09173_);
  and (_09175_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_09176_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  not (_09177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_09178_, _07324_, _09177_);
  nor (_09179_, _09178_, _09176_);
  and (_09180_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_09181_, _07329_, _07389_);
  nor (_09182_, _09181_, _09180_);
  and (_09183_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_09184_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_09185_, _09184_, _09183_);
  and (_09186_, _09185_, _09182_);
  and (_09187_, _09186_, _09179_);
  nor (_09188_, _09187_, _08954_);
  nor (_09189_, _09188_, _09175_);
  not (_09190_, _09189_);
  and (_09191_, _09190_, _08950_);
  nor (_09192_, _09191_, _09174_);
  and (_09193_, _09192_, _09172_);
  and (_09194_, _09193_, _09169_);
  not (_09195_, _09194_);
  and (_09196_, _09195_, _09094_);
  nor (_09197_, _09196_, _09146_);
  nor (_09198_, _09197_, _09098_);
  nor (_09199_, _09198_, _09097_);
  nor (_09200_, _09096_, _08857_);
  not (_09201_, _09200_);
  not (_09202_, _08892_);
  and (_09203_, _09092_, _08869_);
  nor (_09204_, _09195_, _09203_);
  not (_09205_, _07754_);
  and (_09206_, _08887_, _09205_);
  nand (_09207_, _08916_, _06600_);
  nor (_09208_, _09207_, _06829_);
  nor (_09209_, _07754_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_09210_, _06600_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_09211_, _05734_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_09212_, _09211_, _09210_);
  or (_09213_, _09212_, _09209_);
  or (_09214_, _09213_, _09208_);
  or (_09215_, _09214_, _08911_);
  and (_09216_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_09217_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_09218_, _09217_, _09216_);
  and (_09219_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_09220_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_09221_, _09220_, _09219_);
  or (_09222_, _09221_, _09218_);
  or (_09223_, _09222_, _08910_);
  and (_09224_, _09223_, _08888_);
  and (_09225_, _09224_, _09215_);
  or (_09226_, _09225_, _09206_);
  and (_09227_, _09226_, _08872_);
  not (_09228_, _09227_);
  nor (_09229_, _07864_, _08998_);
  and (_09230_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_09231_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_09232_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_09233_, _09232_, _09231_);
  and (_09234_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_09235_, _07329_, _07475_);
  nor (_09236_, _09235_, _09234_);
  and (_09237_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not (_09238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_09239_, _07324_, _09238_);
  nor (_09240_, _09239_, _09237_);
  and (_09241_, _09240_, _09236_);
  and (_09242_, _09241_, _09233_);
  nor (_09243_, _09242_, _08954_);
  nor (_09244_, _09243_, _09230_);
  not (_09245_, _09244_);
  and (_09246_, _09245_, _08949_);
  nor (_09247_, _09246_, _09018_);
  not (_09248_, _09247_);
  nor (_09249_, _09248_, _09229_);
  and (_09250_, _09249_, _09228_);
  and (_09251_, _09250_, _09203_);
  nor (_09252_, _09251_, _09204_);
  nor (_09253_, _09252_, _09202_);
  and (_09254_, _09252_, _09202_);
  nor (_09255_, _09254_, _09253_);
  and (_09256_, _09255_, _09201_);
  nor (_09257_, _07790_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_09258_, _08912_, _06603_);
  and (_09259_, _09258_, _06885_);
  and (_09260_, _08912_, _06599_);
  not (_09261_, _09260_);
  and (_09262_, _08918_, _09261_);
  not (_09263_, _09262_);
  and (_09264_, _09263_, _05717_);
  or (_09265_, _09264_, _09259_);
  or (_09266_, _09265_, _09257_);
  nor (_09267_, _09266_, _08911_);
  and (_09268_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_09269_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_09270_, _09269_, _09268_);
  and (_09271_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_09272_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_09273_, _09272_, _09271_);
  and (_09274_, _09273_, _09270_);
  and (_09275_, _09274_, _08911_);
  or (_09276_, _09275_, _09267_);
  and (_09277_, _09276_, _08888_);
  and (_09278_, _08887_, _07790_);
  nor (_09279_, _09278_, _09277_);
  nand (_09280_, _09279_, _08872_);
  and (_09281_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_09282_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_09283_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_09284_, _09283_, _09282_);
  and (_09285_, _07420_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_09286_, _07417_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_09287_, _09286_, _09285_);
  and (_09288_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_09289_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_09290_, _09289_, _09288_);
  and (_09291_, _09290_, _09287_);
  and (_09292_, _09291_, _09284_);
  nor (_09293_, _09292_, _08954_);
  nor (_09294_, _09293_, _09281_);
  not (_09295_, _09294_);
  and (_09296_, _09295_, _08950_);
  and (_09297_, _08871_, _09071_);
  not (_09298_, _07834_);
  and (_09299_, _09298_, _08942_);
  and (_09300_, _08947_, _07439_);
  or (_09301_, _09300_, _09299_);
  or (_09302_, _09301_, _09297_);
  nor (_09303_, _09302_, _09296_);
  and (_09304_, _09303_, _09280_);
  nor (_09305_, _09304_, _08869_);
  and (_09306_, _06596_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_09307_, _09306_);
  and (_09308_, _05653_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_09309_, _09308_, _09307_);
  and (_09310_, _08916_, _06596_);
  and (_09311_, _09310_, _06885_);
  nor (_09312_, _07768_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_09313_, _09312_, _09311_);
  or (_09314_, _09313_, _09309_);
  nor (_09315_, _09314_, _08911_);
  and (_09316_, _08932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_09317_, _08927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_09318_, _09317_, _09316_);
  and (_09319_, _08925_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_09320_, _08930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_09321_, _09320_, _09319_);
  and (_09322_, _09321_, _09318_);
  and (_09323_, _09322_, _08911_);
  or (_09324_, _09323_, _09315_);
  and (_09325_, _09324_, _08888_);
  and (_09326_, _08887_, _07768_);
  nor (_09327_, _09326_, _09325_);
  nand (_09328_, _09327_, _08872_);
  nor (_09329_, _07852_, _08998_);
  and (_09330_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_09331_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_09332_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_09333_, _09332_, _09331_);
  and (_09334_, _07417_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_09335_, _07329_, _07530_);
  nor (_09336_, _09335_, _09334_);
  and (_09337_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_09338_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_09339_, _09338_, _09337_);
  and (_09340_, _09339_, _09336_);
  and (_09341_, _09340_, _09333_);
  nor (_09342_, _09341_, _08954_);
  nor (_09343_, _09342_, _09330_);
  not (_09344_, _09343_);
  and (_09345_, _09344_, _08950_);
  nor (_09346_, _09345_, _09329_);
  and (_09347_, _09071_, _07624_);
  nor (_09348_, _08284_, _08280_);
  not (_09349_, _09348_);
  and (_09350_, _09349_, _08947_);
  or (_09351_, _09350_, _09347_);
  not (_09352_, _09351_);
  and (_09353_, _09352_, _09346_);
  and (_09354_, _09353_, _09328_);
  not (_09355_, _09354_);
  and (_09356_, _09355_, _09094_);
  nor (_09357_, _09356_, _09305_);
  nand (_09358_, _09357_, _08904_);
  or (_09359_, _09357_, _08904_);
  and (_09360_, _09359_, _09358_);
  not (_09361_, _09360_);
  not (_09362_, _08873_);
  and (_09363_, _09197_, _09098_);
  nor (_09364_, _09363_, _09362_);
  and (_09365_, _09364_, _09361_);
  and (_09366_, _09365_, _09256_);
  and (_09367_, _09366_, _09199_);
  not (_09368_, _09096_);
  and (_09369_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_09370_, _09197_);
  and (_09371_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_09372_, _09371_, _09369_);
  and (_09373_, _09372_, _09357_);
  not (_09374_, _09357_);
  not (_09375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_09376_, _09197_, _09375_);
  and (_09377_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_09378_, _09377_, _09376_);
  and (_09379_, _09378_, _09374_);
  or (_09380_, _09379_, _09373_);
  or (_09381_, _09380_, _09368_);
  not (_09382_, _09252_);
  and (_09383_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_09384_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_09385_, _09384_, _09383_);
  and (_09386_, _09385_, _09357_);
  not (_09387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_09388_, _09197_, _09387_);
  and (_09389_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_09390_, _09389_, _09388_);
  and (_09391_, _09390_, _09374_);
  or (_09392_, _09391_, _09386_);
  or (_09393_, _09392_, _09096_);
  and (_09394_, _09393_, _09382_);
  and (_09395_, _09394_, _09381_);
  or (_09396_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_09397_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_09398_, _09397_, _09396_);
  and (_09399_, _09398_, _09357_);
  or (_09400_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_09401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_09402_, _09197_, _09401_);
  and (_09403_, _09402_, _09400_);
  and (_09404_, _09403_, _09374_);
  or (_09405_, _09404_, _09399_);
  or (_09406_, _09405_, _09368_);
  or (_09407_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_09408_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_09409_, _09408_, _09407_);
  and (_09410_, _09409_, _09357_);
  or (_09411_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_09412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_09413_, _09197_, _09412_);
  and (_09414_, _09413_, _09411_);
  and (_09415_, _09414_, _09374_);
  or (_09416_, _09415_, _09410_);
  or (_09417_, _09416_, _09096_);
  and (_09418_, _09417_, _09252_);
  and (_09419_, _09418_, _09406_);
  or (_09420_, _09419_, _09395_);
  or (_09421_, _09420_, _09367_);
  not (_09422_, _09367_);
  or (_09423_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_09424_, _09423_, _12493_);
  and (_10115_, _09424_, _09421_);
  nor (_09425_, _08898_, _09362_);
  nor (_09426_, _08904_, _09362_);
  and (_09427_, _09426_, _09425_);
  nor (_09428_, _08856_, _09362_);
  and (_09429_, _08892_, _08873_);
  and (_09430_, _09429_, _09428_);
  and (_09431_, _09430_, _09427_);
  and (_09432_, _09056_, _08873_);
  and (_09433_, _09432_, _09431_);
  not (_09434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_09435_, _09431_, _09434_);
  or (_10127_, _09435_, _09433_);
  nor (_09436_, _09426_, _09425_);
  nor (_09437_, _09429_, _09428_);
  and (_09438_, _09437_, _08873_);
  and (_09439_, _09438_, _09436_);
  and (_09440_, _09106_, _08873_);
  and (_09441_, _09440_, _09439_);
  not (_09442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_09443_, _09439_, _09442_);
  or (_10374_, _09443_, _09441_);
  and (_09444_, _09266_, _08873_);
  and (_09445_, _09444_, _09439_);
  not (_09446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_09447_, _09439_, _09446_);
  or (_10380_, _09447_, _09445_);
  and (_09448_, _08923_, _08873_);
  and (_09449_, _09448_, _09439_);
  not (_09450_, _09439_);
  and (_09451_, _09450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_10385_, _09451_, _09449_);
  and (_09452_, _09155_, _08873_);
  and (_09453_, _09452_, _09439_);
  and (_09454_, _09450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_10390_, _09454_, _09453_);
  and (_09455_, _09314_, _08873_);
  and (_09456_, _09455_, _09439_);
  and (_09457_, _09450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_10395_, _09457_, _09456_);
  and (_09458_, _08983_, _08873_);
  and (_09459_, _09458_, _09439_);
  and (_09460_, _09450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_10400_, _09460_, _09459_);
  and (_09461_, _09214_, _08873_);
  and (_09462_, _09461_, _09439_);
  and (_09463_, _09450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_10405_, _09463_, _09462_);
  and (_09464_, _09439_, _09432_);
  and (_09465_, _09450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_10408_, _09465_, _09464_);
  and (_09466_, _09425_, _08904_);
  and (_09467_, _09466_, _09437_);
  and (_09468_, _09467_, _09440_);
  not (_09469_, _09467_);
  and (_09470_, _09469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_10415_, _09470_, _09468_);
  and (_09471_, _09467_, _09444_);
  and (_09472_, _09469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_10419_, _09472_, _09471_);
  and (_09473_, _09467_, _09448_);
  and (_09474_, _09469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_10422_, _09474_, _09473_);
  and (_09475_, _09467_, _09452_);
  and (_09476_, _09469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_10426_, _09476_, _09475_);
  and (_09477_, _09467_, _09455_);
  not (_09478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_09479_, _09467_, _09478_);
  or (_10429_, _09479_, _09477_);
  and (_09480_, _09467_, _09458_);
  not (_09481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_09482_, _09467_, _09481_);
  or (_10433_, _09482_, _09480_);
  and (_09483_, _09467_, _09461_);
  and (_09484_, _09469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_10436_, _09484_, _09483_);
  and (_09485_, _09467_, _09432_);
  and (_09486_, _09469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_10439_, _09486_, _09485_);
  and (_09487_, _09426_, _08898_);
  and (_09488_, _09487_, _09437_);
  and (_09489_, _09488_, _09440_);
  not (_09490_, _09488_);
  and (_09491_, _09490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_10446_, _09491_, _09489_);
  and (_09492_, _09488_, _09444_);
  and (_09493_, _09490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_10449_, _09493_, _09492_);
  and (_09494_, _09488_, _09448_);
  not (_09495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_09496_, _09488_, _09495_);
  or (_10453_, _09496_, _09494_);
  and (_09497_, _09488_, _09452_);
  and (_09498_, _09490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_10456_, _09498_, _09497_);
  and (_09499_, _09488_, _09455_);
  not (_09500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_09501_, _09488_, _09500_);
  or (_10460_, _09501_, _09499_);
  and (_09502_, _09488_, _09458_);
  not (_09503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_09504_, _09488_, _09503_);
  or (_10463_, _09504_, _09502_);
  and (_09505_, _09488_, _09461_);
  and (_09506_, _09490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_10467_, _09506_, _09505_);
  and (_09507_, _09488_, _09432_);
  not (_09508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_09509_, _09488_, _09508_);
  or (_10469_, _09509_, _09507_);
  and (_09510_, _09437_, _09427_);
  and (_09511_, _09510_, _09440_);
  not (_09512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_09513_, _09510_, _09512_);
  or (_10475_, _09513_, _09511_);
  and (_09514_, _09510_, _09444_);
  not (_09515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_09516_, _09510_, _09515_);
  or (_10478_, _09516_, _09514_);
  and (_09517_, _09510_, _09448_);
  not (_09518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_09519_, _09510_, _09518_);
  or (_10482_, _09519_, _09517_);
  and (_09520_, _09510_, _09452_);
  not (_09521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_09522_, _09510_, _09521_);
  or (_10485_, _09522_, _09520_);
  and (_09523_, _09510_, _09455_);
  not (_09524_, _09510_);
  and (_09525_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_10489_, _09525_, _09523_);
  and (_09526_, _09510_, _09458_);
  and (_09527_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_10492_, _09527_, _09526_);
  and (_09528_, _09510_, _09461_);
  and (_09529_, _09524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_10496_, _09529_, _09528_);
  and (_09530_, _09510_, _09432_);
  nor (_09531_, _09510_, _09375_);
  or (_10498_, _09531_, _09530_);
  and (_09532_, _09428_, _09202_);
  and (_09533_, _09532_, _09436_);
  and (_09534_, _09533_, _09440_);
  not (_09535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_09536_, _09533_, _09535_);
  or (_10505_, _09536_, _09534_);
  and (_09537_, _09533_, _09444_);
  not (_09538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_09539_, _09533_, _09538_);
  or (_10509_, _09539_, _09537_);
  and (_09540_, _09533_, _09448_);
  not (_09541_, _09533_);
  and (_09542_, _09541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_10512_, _09542_, _09540_);
  and (_09543_, _09533_, _09452_);
  not (_09544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_09545_, _09533_, _09544_);
  or (_10516_, _09545_, _09543_);
  and (_09546_, _09533_, _09455_);
  and (_09547_, _09541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_10519_, _09547_, _09546_);
  and (_09548_, _09533_, _09458_);
  and (_09549_, _09541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_10523_, _09549_, _09548_);
  and (_09550_, _09533_, _09461_);
  not (_09551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_09552_, _09533_, _09551_);
  or (_10526_, _09552_, _09550_);
  and (_09553_, _09533_, _09432_);
  and (_09554_, _09541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_10529_, _09554_, _09553_);
  and (_09555_, _09532_, _09466_);
  and (_09556_, _09555_, _09440_);
  not (_09557_, _09555_);
  and (_09558_, _09557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_10533_, _09558_, _09556_);
  and (_09559_, _09555_, _09444_);
  and (_09560_, _09557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_10537_, _09560_, _09559_);
  and (_09561_, _09555_, _09448_);
  and (_09562_, _09557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_10540_, _09562_, _09561_);
  and (_09563_, _09555_, _09452_);
  not (_09564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_09565_, _09555_, _09564_);
  or (_10544_, _09565_, _09563_);
  and (_09566_, _09555_, _09455_);
  not (_09567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_09568_, _09555_, _09567_);
  or (_10547_, _09568_, _09566_);
  and (_09569_, _09555_, _09458_);
  not (_09570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_09571_, _09555_, _09570_);
  or (_10551_, _09571_, _09569_);
  and (_09572_, _09555_, _09461_);
  and (_09573_, _09557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_10554_, _09573_, _09572_);
  and (_09574_, _09555_, _09432_);
  and (_09575_, _09557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_10557_, _09575_, _09574_);
  and (_09576_, _09532_, _09487_);
  and (_09577_, _09576_, _09440_);
  not (_09578_, _09576_);
  and (_09579_, _09578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_10561_, _09579_, _09577_);
  and (_09580_, _09576_, _09444_);
  and (_09581_, _09578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_10565_, _09581_, _09580_);
  and (_09582_, _09576_, _09448_);
  not (_09583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_09584_, _09576_, _09583_);
  or (_10568_, _09584_, _09582_);
  and (_09585_, _09576_, _09452_);
  and (_09586_, _09578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_10572_, _09586_, _09585_);
  and (_09587_, _09576_, _09455_);
  not (_09588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_09589_, _09576_, _09588_);
  or (_10575_, _09589_, _09587_);
  and (_09590_, _09576_, _09458_);
  not (_09591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_09592_, _09576_, _09591_);
  or (_10579_, _09592_, _09590_);
  and (_09593_, _09576_, _09461_);
  not (_09594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_09595_, _09576_, _09594_);
  or (_10582_, _09595_, _09593_);
  and (_09596_, _09576_, _09432_);
  not (_09597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_09598_, _09576_, _09597_);
  or (_10585_, _09598_, _09596_);
  and (_09599_, _09532_, _09427_);
  and (_09600_, _09599_, _09440_);
  not (_09601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_09602_, _09599_, _09601_);
  or (_10589_, _09602_, _09600_);
  and (_09603_, _09599_, _09444_);
  not (_09604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_09605_, _09599_, _09604_);
  or (_10593_, _09605_, _09603_);
  and (_09606_, _09599_, _09448_);
  not (_09607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_09608_, _09599_, _09607_);
  or (_10596_, _09608_, _09606_);
  and (_09609_, _09599_, _09452_);
  not (_09610_, _09599_);
  and (_09611_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_10600_, _09611_, _09609_);
  and (_09612_, _09599_, _09455_);
  and (_09613_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_10603_, _09613_, _09612_);
  and (_09614_, _09599_, _09458_);
  and (_09615_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_10607_, _09615_, _09614_);
  and (_09616_, _09599_, _09461_);
  and (_09617_, _09610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_10610_, _09617_, _09616_);
  and (_09618_, _09599_, _09432_);
  nor (_09619_, _09599_, _09387_);
  or (_10613_, _09619_, _09618_);
  and (_09620_, _09429_, _08856_);
  and (_09621_, _09620_, _09436_);
  and (_09622_, _09621_, _09440_);
  not (_09623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_09624_, _09621_, _09623_);
  or (_10620_, _09624_, _09622_);
  and (_09625_, _09621_, _09444_);
  not (_09626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_09627_, _09621_, _09626_);
  or (_10623_, _09627_, _09625_);
  and (_09628_, _09621_, _09448_);
  not (_09629_, _09621_);
  and (_09630_, _09629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_10627_, _09630_, _09628_);
  and (_09631_, _09621_, _09452_);
  and (_09632_, _09629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_10630_, _09632_, _09631_);
  and (_09633_, _09621_, _09455_);
  and (_09634_, _09629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_10634_, _09634_, _09633_);
  and (_09635_, _09621_, _09458_);
  and (_09636_, _09629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_10637_, _09636_, _09635_);
  and (_09637_, _09621_, _09461_);
  and (_09638_, _09629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_10641_, _09638_, _09637_);
  and (_09639_, _09621_, _09432_);
  and (_09640_, _09629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_10644_, _09640_, _09639_);
  and (_09641_, _09620_, _09466_);
  and (_09642_, _09641_, _09440_);
  not (_09643_, _09641_);
  and (_09644_, _09643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_10648_, _09644_, _09642_);
  and (_09645_, _09641_, _09444_);
  and (_09646_, _09643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_10652_, _09646_, _09645_);
  and (_09647_, _09641_, _09448_);
  and (_09648_, _09643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_10655_, _09648_, _09647_);
  and (_09649_, _09641_, _09452_);
  and (_09650_, _09643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_10659_, _09650_, _09649_);
  and (_09651_, _09641_, _09455_);
  not (_09652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_09653_, _09641_, _09652_);
  or (_10662_, _09653_, _09651_);
  and (_09654_, _09641_, _09458_);
  not (_09655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_09656_, _09641_, _09655_);
  or (_10666_, _09656_, _09654_);
  and (_09657_, _09641_, _09461_);
  and (_09658_, _09643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_10669_, _09658_, _09657_);
  and (_09659_, _09641_, _09432_);
  and (_09660_, _09643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_10672_, _09660_, _09659_);
  and (_09661_, _09620_, _09487_);
  and (_09662_, _09661_, _09440_);
  not (_09663_, _09661_);
  and (_09664_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_10676_, _09664_, _09662_);
  and (_09665_, _09661_, _09444_);
  and (_09666_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_10680_, _09666_, _09665_);
  and (_09667_, _09661_, _09448_);
  not (_09668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_09669_, _09661_, _09668_);
  or (_10683_, _09669_, _09667_);
  and (_09670_, _09661_, _09452_);
  not (_09671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_09672_, _09661_, _09671_);
  or (_10687_, _09672_, _09670_);
  and (_09673_, _09661_, _09455_);
  not (_09674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_09675_, _09661_, _09674_);
  or (_10690_, _09675_, _09673_);
  and (_09676_, _09661_, _09458_);
  not (_09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_09678_, _09661_, _09677_);
  or (_10694_, _09678_, _09676_);
  and (_09679_, _09661_, _09461_);
  and (_09680_, _09663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_10697_, _09680_, _09679_);
  and (_09681_, _09661_, _09432_);
  nor (_09682_, _09661_, _09401_);
  or (_10700_, _09682_, _09681_);
  and (_09683_, _09620_, _09427_);
  and (_09684_, _09683_, _09440_);
  not (_09685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_09686_, _09683_, _09685_);
  or (_10704_, _09686_, _09684_);
  and (_09687_, _09683_, _09444_);
  not (_09688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_09689_, _09683_, _09688_);
  or (_10708_, _09689_, _09687_);
  and (_09690_, _09683_, _09448_);
  not (_09691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_09692_, _09683_, _09691_);
  or (_10711_, _09692_, _09690_);
  and (_09693_, _09683_, _09452_);
  not (_09694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_09695_, _09683_, _09694_);
  or (_10715_, _09695_, _09693_);
  and (_09696_, _09683_, _09455_);
  not (_09697_, _09683_);
  and (_09698_, _09697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_10718_, _09698_, _09696_);
  and (_09699_, _09683_, _09458_);
  and (_09700_, _09697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_10722_, _09700_, _09699_);
  and (_09701_, _09683_, _09461_);
  and (_09702_, _09697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_10725_, _09702_, _09701_);
  and (_09703_, _09683_, _09432_);
  not (_09704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_09705_, _09683_, _09704_);
  or (_10728_, _09705_, _09703_);
  and (_09706_, _09436_, _09430_);
  and (_09707_, _09706_, _09440_);
  not (_09708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_09709_, _09706_, _09708_);
  or (_10733_, _09709_, _09707_);
  and (_09710_, _09706_, _09444_);
  not (_09711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_09712_, _09706_, _09711_);
  or (_10737_, _09712_, _09710_);
  and (_09713_, _09706_, _09448_);
  not (_09714_, _09706_);
  and (_09715_, _09714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_10740_, _09715_, _09713_);
  and (_09716_, _09706_, _09452_);
  not (_09717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_09718_, _09706_, _09717_);
  or (_10744_, _09718_, _09716_);
  and (_09719_, _09706_, _09455_);
  and (_09720_, _09714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_10747_, _09720_, _09719_);
  and (_09721_, _09706_, _09458_);
  and (_09722_, _09714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_10751_, _09722_, _09721_);
  and (_09723_, _09706_, _09461_);
  not (_09724_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_09725_, _09706_, _09724_);
  or (_10754_, _09725_, _09723_);
  and (_09726_, _09706_, _09432_);
  and (_09727_, _09714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_10757_, _09727_, _09726_);
  and (_09728_, _09466_, _09430_);
  and (_09729_, _09728_, _09440_);
  not (_09730_, _09728_);
  and (_09731_, _09730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_10761_, _09731_, _09729_);
  and (_09732_, _09728_, _09444_);
  and (_09733_, _09730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_10765_, _09733_, _09732_);
  and (_09734_, _09728_, _09448_);
  and (_09735_, _09730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_10768_, _09735_, _09734_);
  and (_09736_, _09728_, _09452_);
  not (_09737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_09738_, _09728_, _09737_);
  or (_10772_, _09738_, _09736_);
  and (_09739_, _09728_, _09455_);
  not (_09740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_09741_, _09728_, _09740_);
  or (_10775_, _09741_, _09739_);
  and (_09742_, _09728_, _09458_);
  not (_09743_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_09744_, _09728_, _09743_);
  or (_10779_, _09744_, _09742_);
  and (_09745_, _09728_, _09461_);
  not (_09746_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_09747_, _09728_, _09746_);
  or (_10782_, _09747_, _09745_);
  and (_09748_, _09728_, _09432_);
  and (_09749_, _09730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_10785_, _09749_, _09748_);
  and (_09750_, _09487_, _09430_);
  and (_09751_, _09750_, _09440_);
  not (_09752_, _09750_);
  and (_09753_, _09752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_10789_, _09753_, _09751_);
  and (_09754_, _09750_, _09444_);
  and (_09755_, _09752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_10793_, _09755_, _09754_);
  and (_09756_, _09750_, _09448_);
  not (_09757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_09758_, _09750_, _09757_);
  or (_10796_, _09758_, _09756_);
  and (_09759_, _09750_, _09452_);
  not (_09760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_09761_, _09750_, _09760_);
  or (_10800_, _09761_, _09759_);
  and (_09762_, _09750_, _09455_);
  not (_09763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_09764_, _09750_, _09763_);
  or (_10803_, _09764_, _09762_);
  and (_09765_, _09750_, _09458_);
  not (_09766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_09767_, _09750_, _09766_);
  or (_10807_, _09767_, _09765_);
  and (_09768_, _09750_, _09461_);
  not (_09769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_09770_, _09750_, _09769_);
  or (_10810_, _09770_, _09768_);
  and (_09771_, _09750_, _09432_);
  nor (_09772_, _09750_, _09412_);
  or (_10813_, _09772_, _09771_);
  and (_09773_, _09440_, _09431_);
  not (_09774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_09775_, _09431_, _09774_);
  or (_10817_, _09775_, _09773_);
  and (_09776_, _09444_, _09431_);
  not (_09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_09778_, _09431_, _09777_);
  or (_10821_, _09778_, _09776_);
  and (_09779_, _09448_, _09431_);
  not (_09780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_09781_, _09431_, _09780_);
  or (_10824_, _09781_, _09779_);
  and (_09782_, _09452_, _09431_);
  not (_09783_, _09431_);
  and (_09784_, _09783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_10828_, _09784_, _09782_);
  and (_09785_, _09455_, _09431_);
  and (_09786_, _09783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_10831_, _09786_, _09785_);
  and (_09787_, _09458_, _09431_);
  and (_09788_, _09783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_10835_, _09788_, _09787_);
  and (_09789_, _09461_, _09431_);
  not (_09790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_09791_, _09431_, _09790_);
  or (_10838_, _09791_, _09789_);
  or (_09792_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_09793_, _09197_, _09442_);
  and (_09794_, _09793_, _09357_);
  and (_09795_, _09794_, _09792_);
  nor (_09796_, _09197_, _09512_);
  and (_09797_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_09798_, _09797_, _09796_);
  and (_09799_, _09798_, _09374_);
  or (_09800_, _09799_, _09795_);
  or (_09801_, _09800_, _09368_);
  or (_09802_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_09803_, _09197_, _09535_);
  and (_09804_, _09803_, _09357_);
  and (_09805_, _09804_, _09802_);
  nor (_09806_, _09197_, _09601_);
  and (_09807_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_09808_, _09807_, _09806_);
  and (_09809_, _09808_, _09374_);
  or (_09810_, _09809_, _09805_);
  or (_09811_, _09810_, _09096_);
  and (_09812_, _09811_, _09382_);
  and (_09813_, _09812_, _09801_);
  nand (_09814_, _09197_, _09623_);
  or (_09815_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_09816_, _09815_, _09814_);
  and (_09817_, _09816_, _09357_);
  and (_09818_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_09819_, _09197_, _09685_);
  or (_09820_, _09819_, _09818_);
  and (_09821_, _09820_, _09374_);
  or (_09822_, _09821_, _09817_);
  or (_09823_, _09822_, _09368_);
  nand (_09824_, _09197_, _09708_);
  or (_09825_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_09826_, _09825_, _09824_);
  and (_09827_, _09826_, _09357_);
  and (_09828_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_09829_, _09197_, _09774_);
  or (_09830_, _09829_, _09828_);
  and (_09831_, _09830_, _09374_);
  or (_09832_, _09831_, _09827_);
  or (_09833_, _09832_, _09096_);
  and (_09834_, _09833_, _09252_);
  and (_09835_, _09834_, _09823_);
  or (_09836_, _09835_, _09813_);
  or (_09837_, _09836_, _09367_);
  or (_09838_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_09839_, _09838_, _12493_);
  and (_12471_, _09839_, _09837_);
  or (_09840_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_09841_, _09197_, _09446_);
  and (_09842_, _09841_, _09357_);
  and (_09843_, _09842_, _09840_);
  nor (_09844_, _09197_, _09515_);
  and (_09845_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_09846_, _09845_, _09844_);
  and (_09847_, _09846_, _09374_);
  or (_09848_, _09847_, _09843_);
  or (_09849_, _09848_, _09368_);
  or (_09850_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_09851_, _09197_, _09538_);
  and (_09852_, _09851_, _09357_);
  and (_09853_, _09852_, _09850_);
  nor (_09854_, _09197_, _09604_);
  and (_09855_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_09856_, _09855_, _09854_);
  and (_09857_, _09856_, _09374_);
  or (_09858_, _09857_, _09853_);
  or (_09859_, _09858_, _09096_);
  and (_09860_, _09859_, _09382_);
  and (_09861_, _09860_, _09849_);
  nand (_09862_, _09197_, _09626_);
  or (_09863_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_09864_, _09863_, _09862_);
  and (_09865_, _09864_, _09357_);
  and (_09866_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_09867_, _09197_, _09688_);
  or (_09868_, _09867_, _09866_);
  and (_09869_, _09868_, _09374_);
  or (_09870_, _09869_, _09865_);
  or (_09871_, _09870_, _09368_);
  nand (_09872_, _09197_, _09711_);
  or (_09873_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_09874_, _09873_, _09872_);
  and (_09875_, _09874_, _09357_);
  and (_09876_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_09877_, _09197_, _09777_);
  or (_09878_, _09877_, _09876_);
  and (_09879_, _09878_, _09374_);
  or (_09880_, _09879_, _09875_);
  or (_09881_, _09880_, _09096_);
  and (_09882_, _09881_, _09252_);
  and (_09883_, _09882_, _09871_);
  or (_09884_, _09883_, _09861_);
  or (_09885_, _09884_, _09367_);
  or (_09886_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_09887_, _09886_, _12493_);
  and (_12473_, _09887_, _09885_);
  and (_09888_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_09889_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_09890_, _09889_, _09888_);
  and (_09891_, _09890_, _09357_);
  nor (_09892_, _09197_, _09518_);
  and (_09893_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_09894_, _09893_, _09892_);
  and (_09895_, _09894_, _09374_);
  or (_09896_, _09895_, _09891_);
  or (_09897_, _09896_, _09368_);
  and (_09898_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_09899_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_09900_, _09899_, _09898_);
  and (_09901_, _09900_, _09357_);
  nor (_09902_, _09197_, _09607_);
  and (_09903_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_09904_, _09903_, _09902_);
  and (_09905_, _09904_, _09374_);
  or (_09906_, _09905_, _09901_);
  or (_09907_, _09906_, _09096_);
  and (_09908_, _09907_, _09382_);
  and (_09909_, _09908_, _09897_);
  or (_09910_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_09911_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_09912_, _09911_, _09910_);
  and (_09913_, _09912_, _09357_);
  or (_09914_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_09915_, _09197_, _09668_);
  and (_09916_, _09915_, _09914_);
  and (_09917_, _09916_, _09374_);
  or (_09918_, _09917_, _09913_);
  or (_09919_, _09918_, _09368_);
  or (_09920_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_09921_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_09922_, _09921_, _09920_);
  and (_09923_, _09922_, _09357_);
  or (_09924_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_09925_, _09197_, _09757_);
  and (_09926_, _09925_, _09924_);
  and (_09927_, _09926_, _09374_);
  or (_09928_, _09927_, _09923_);
  or (_09929_, _09928_, _09096_);
  and (_09930_, _09929_, _09252_);
  and (_09931_, _09930_, _09919_);
  or (_09932_, _09931_, _09909_);
  or (_09933_, _09932_, _09367_);
  or (_09934_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_09935_, _09934_, _12493_);
  and (_12475_, _09935_, _09933_);
  and (_09936_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_09937_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_09938_, _09937_, _09936_);
  and (_09939_, _09938_, _09357_);
  nor (_09940_, _09197_, _09521_);
  and (_09941_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_09942_, _09941_, _09940_);
  and (_09943_, _09942_, _09374_);
  or (_09944_, _09943_, _09939_);
  or (_09945_, _09944_, _09368_);
  and (_09946_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_09947_, _09197_, _09564_);
  or (_09948_, _09947_, _09946_);
  and (_09949_, _09948_, _09357_);
  and (_09950_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_09951_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_09952_, _09951_, _09950_);
  and (_09953_, _09952_, _09374_);
  or (_09954_, _09953_, _09949_);
  or (_09955_, _09954_, _09096_);
  and (_09956_, _09955_, _09382_);
  and (_09957_, _09956_, _09945_);
  or (_09958_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_09959_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_09960_, _09959_, _09958_);
  and (_09961_, _09960_, _09357_);
  or (_09962_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_09963_, _09197_, _09671_);
  and (_09964_, _09963_, _09962_);
  and (_09965_, _09964_, _09374_);
  or (_09966_, _09965_, _09961_);
  or (_09967_, _09966_, _09368_);
  nand (_09968_, _09197_, _09717_);
  or (_09969_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_09970_, _09969_, _09968_);
  and (_09971_, _09970_, _09357_);
  or (_09972_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_09973_, _09197_, _09760_);
  and (_09975_, _09973_, _09972_);
  and (_09977_, _09975_, _09374_);
  or (_09979_, _09977_, _09971_);
  or (_09981_, _09979_, _09096_);
  and (_09983_, _09981_, _09252_);
  and (_09985_, _09983_, _09967_);
  or (_09987_, _09985_, _09957_);
  or (_09989_, _09987_, _09367_);
  or (_09991_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_09993_, _09991_, _12493_);
  and (_12477_, _09993_, _09989_);
  and (_09996_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_09998_, _09197_, _09478_);
  or (_10000_, _09998_, _09996_);
  and (_10002_, _10000_, _09357_);
  or (_10004_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_10006_, _09197_, _09500_);
  and (_10008_, _10006_, _10004_);
  and (_10010_, _10008_, _09374_);
  or (_10012_, _10010_, _10002_);
  or (_10014_, _10012_, _09368_);
  and (_10016_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_10018_, _09197_, _09567_);
  or (_10020_, _10018_, _10016_);
  and (_10022_, _10020_, _09357_);
  or (_10024_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_10026_, _09197_, _09588_);
  and (_10028_, _10026_, _10024_);
  and (_10029_, _10028_, _09374_);
  or (_10030_, _10029_, _10022_);
  or (_10031_, _10030_, _09096_);
  and (_10032_, _10031_, _09382_);
  and (_10033_, _10032_, _10014_);
  and (_10034_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_10035_, _09197_, _09652_);
  or (_10036_, _10035_, _10034_);
  and (_10037_, _10036_, _09357_);
  or (_10038_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_10039_, _09197_, _09674_);
  and (_10040_, _10039_, _10038_);
  and (_10041_, _10040_, _09374_);
  or (_10042_, _10041_, _10037_);
  or (_10043_, _10042_, _09368_);
  and (_10044_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_10045_, _09197_, _09740_);
  or (_10046_, _10045_, _10044_);
  and (_10047_, _10046_, _09357_);
  or (_10048_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_10049_, _09197_, _09763_);
  and (_10050_, _10049_, _10048_);
  and (_10051_, _10050_, _09374_);
  or (_10052_, _10051_, _10047_);
  or (_10053_, _10052_, _09096_);
  and (_10054_, _10053_, _09252_);
  and (_10055_, _10054_, _10043_);
  or (_10056_, _10055_, _10033_);
  or (_10057_, _10056_, _09367_);
  or (_10058_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_10059_, _10058_, _12493_);
  and (_12478_, _10059_, _10057_);
  and (_10060_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_10061_, _09197_, _09481_);
  or (_10062_, _10061_, _10060_);
  and (_10063_, _10062_, _09357_);
  or (_10064_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_10065_, _09197_, _09503_);
  and (_10066_, _10065_, _10064_);
  and (_10067_, _10066_, _09374_);
  or (_10068_, _10067_, _10063_);
  or (_10069_, _10068_, _09368_);
  and (_10070_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_10071_, _09197_, _09570_);
  or (_10072_, _10071_, _10070_);
  and (_10073_, _10072_, _09357_);
  or (_10074_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_10075_, _09197_, _09591_);
  and (_10076_, _10075_, _10074_);
  and (_10077_, _10076_, _09374_);
  or (_10078_, _10077_, _10073_);
  or (_10079_, _10078_, _09096_);
  and (_10080_, _10079_, _09382_);
  and (_10081_, _10080_, _10069_);
  and (_10082_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_10083_, _09197_, _09655_);
  or (_10084_, _10083_, _10082_);
  and (_10085_, _10084_, _09357_);
  or (_10086_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_10087_, _09197_, _09677_);
  and (_10088_, _10087_, _10086_);
  and (_10089_, _10088_, _09374_);
  or (_10090_, _10089_, _10085_);
  or (_10091_, _10090_, _09368_);
  and (_10092_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_10093_, _09197_, _09743_);
  or (_10094_, _10093_, _10092_);
  and (_10095_, _10094_, _09357_);
  or (_10096_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_10097_, _09197_, _09766_);
  and (_10098_, _10097_, _10096_);
  and (_10099_, _10098_, _09374_);
  or (_10100_, _10099_, _10095_);
  or (_10101_, _10100_, _09096_);
  and (_10102_, _10101_, _09252_);
  and (_10103_, _10102_, _10091_);
  or (_10104_, _10103_, _10081_);
  or (_10105_, _10104_, _09367_);
  or (_10106_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_10107_, _10106_, _12493_);
  and (_12480_, _10107_, _10105_);
  and (_10108_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_10109_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_10110_, _10109_, _10108_);
  and (_10111_, _10110_, _09357_);
  and (_10112_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_10113_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_10114_, _10113_, _10112_);
  and (_10116_, _10114_, _09374_);
  or (_10117_, _10116_, _10111_);
  or (_10118_, _10117_, _09368_);
  or (_10119_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand (_10120_, _09197_, _09551_);
  and (_10121_, _10120_, _09357_);
  and (_10122_, _10121_, _10119_);
  or (_10123_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nand (_10124_, _09197_, _09594_);
  and (_10125_, _10124_, _10123_);
  and (_10126_, _10125_, _09374_);
  or (_10128_, _10126_, _10122_);
  or (_10129_, _10128_, _09096_);
  and (_10130_, _10129_, _09382_);
  and (_10131_, _10130_, _10118_);
  or (_10132_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_10133_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_10134_, _10133_, _10132_);
  and (_10135_, _10134_, _09357_);
  or (_10136_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_10137_, _09370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_10138_, _10137_, _10136_);
  and (_10139_, _10138_, _09374_);
  or (_10140_, _10139_, _10135_);
  or (_10141_, _10140_, _09368_);
  nand (_10142_, _09197_, _09724_);
  or (_10143_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_10144_, _10143_, _10142_);
  and (_10145_, _10144_, _09357_);
  or (_10146_, _09197_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_10147_, _09197_, _09769_);
  and (_10148_, _10147_, _10146_);
  and (_10149_, _10148_, _09374_);
  or (_10150_, _10149_, _10145_);
  or (_10151_, _10150_, _09096_);
  and (_10152_, _10151_, _09252_);
  and (_10153_, _10152_, _10141_);
  or (_10154_, _10153_, _10131_);
  or (_10155_, _10154_, _09367_);
  or (_10156_, _09422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_10157_, _10156_, _12493_);
  and (_12482_, _10157_, _10155_);
  nor (_10158_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_10159_, \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10160_, _10159_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nor (_10161_, _10160_, _10158_);
  or (_10162_, _10161_, rst);
  or (_10163_, \oc8051_gm_cxrom_1.cell0.data [7], _12493_);
  and (_12490_, _10163_, _10162_);
  nor (_10164_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10165_, \oc8051_gm_cxrom_1.cell0.data [0], _10159_);
  nor (_10166_, _10165_, _10164_);
  or (_10167_, _10166_, rst);
  or (_10168_, \oc8051_gm_cxrom_1.cell0.data [0], _12493_);
  and (_12497_, _10168_, _10167_);
  nor (_10169_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10170_, \oc8051_gm_cxrom_1.cell0.data [1], _10159_);
  nor (_10171_, _10170_, _10169_);
  or (_10172_, _10171_, rst);
  or (_10173_, \oc8051_gm_cxrom_1.cell0.data [1], _12493_);
  and (_12501_, _10173_, _10172_);
  nor (_10174_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10175_, \oc8051_gm_cxrom_1.cell0.data [2], _10159_);
  nor (_10176_, _10175_, _10174_);
  or (_10177_, _10176_, rst);
  or (_10178_, \oc8051_gm_cxrom_1.cell0.data [2], _12493_);
  and (_12504_, _10178_, _10177_);
  nor (_10179_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10180_, \oc8051_gm_cxrom_1.cell0.data [3], _10159_);
  nor (_10181_, _10180_, _10179_);
  or (_10182_, _10181_, rst);
  or (_10183_, \oc8051_gm_cxrom_1.cell0.data [3], _12493_);
  and (_12508_, _10183_, _10182_);
  nor (_10184_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10185_, \oc8051_gm_cxrom_1.cell0.data [4], _10159_);
  nor (_10186_, _10185_, _10184_);
  or (_10187_, _10186_, rst);
  or (_10188_, \oc8051_gm_cxrom_1.cell0.data [4], _12493_);
  and (_12512_, _10188_, _10187_);
  nor (_10189_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10190_, \oc8051_gm_cxrom_1.cell0.data [5], _10159_);
  nor (_10191_, _10190_, _10189_);
  or (_10192_, _10191_, rst);
  or (_10193_, \oc8051_gm_cxrom_1.cell0.data [5], _12493_);
  and (_12516_, _10193_, _10192_);
  nor (_10194_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  nor (_10195_, \oc8051_gm_cxrom_1.cell0.data [6], _10159_);
  nor (_10196_, _10195_, _10194_);
  or (_10197_, _10196_, rst);
  or (_10198_, \oc8051_gm_cxrom_1.cell0.data [6], _12493_);
  and (_12520_, _10198_, _10197_);
  nor (_10199_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_10200_, \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10201_, _10200_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nor (_10202_, _10201_, _10199_);
  or (_10203_, _10202_, rst);
  or (_10204_, \oc8051_gm_cxrom_1.cell1.data [7], _12493_);
  and (_12541_, _10204_, _10203_);
  nor (_10205_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10206_, \oc8051_gm_cxrom_1.cell1.data [0], _10200_);
  nor (_10207_, _10206_, _10205_);
  or (_10208_, _10207_, rst);
  or (_10209_, \oc8051_gm_cxrom_1.cell1.data [0], _12493_);
  and (_12548_, _10209_, _10208_);
  nor (_10210_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10211_, \oc8051_gm_cxrom_1.cell1.data [1], _10200_);
  nor (_10212_, _10211_, _10210_);
  or (_10213_, _10212_, rst);
  or (_10214_, \oc8051_gm_cxrom_1.cell1.data [1], _12493_);
  and (_12551_, _10214_, _10213_);
  nor (_10215_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10216_, \oc8051_gm_cxrom_1.cell1.data [2], _10200_);
  nor (_10217_, _10216_, _10215_);
  or (_10218_, _10217_, rst);
  or (_10219_, \oc8051_gm_cxrom_1.cell1.data [2], _12493_);
  and (_12555_, _10219_, _10218_);
  nor (_10220_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10221_, \oc8051_gm_cxrom_1.cell1.data [3], _10200_);
  nor (_10222_, _10221_, _10220_);
  or (_10223_, _10222_, rst);
  or (_10224_, \oc8051_gm_cxrom_1.cell1.data [3], _12493_);
  and (_12559_, _10224_, _10223_);
  nor (_10225_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10226_, \oc8051_gm_cxrom_1.cell1.data [4], _10200_);
  nor (_10227_, _10226_, _10225_);
  or (_10228_, _10227_, rst);
  or (_10229_, \oc8051_gm_cxrom_1.cell1.data [4], _12493_);
  and (_12563_, _10229_, _10228_);
  nor (_10230_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10231_, \oc8051_gm_cxrom_1.cell1.data [5], _10200_);
  nor (_10232_, _10231_, _10230_);
  or (_10233_, _10232_, rst);
  or (_10234_, \oc8051_gm_cxrom_1.cell1.data [5], _12493_);
  and (_12567_, _10234_, _10233_);
  nor (_10235_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  nor (_10236_, \oc8051_gm_cxrom_1.cell1.data [6], _10200_);
  nor (_10237_, _10236_, _10235_);
  or (_10238_, _10237_, rst);
  or (_10239_, \oc8051_gm_cxrom_1.cell1.data [6], _12493_);
  and (_12571_, _10239_, _10238_);
  nor (_10240_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_10241_, \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10242_, _10241_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nor (_10243_, _10242_, _10240_);
  or (_10244_, _10243_, rst);
  or (_10245_, \oc8051_gm_cxrom_1.cell2.data [7], _12493_);
  and (_12592_, _10245_, _10244_);
  nor (_10246_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10247_, \oc8051_gm_cxrom_1.cell2.data [0], _10241_);
  nor (_10248_, _10247_, _10246_);
  or (_10249_, _10248_, rst);
  or (_10250_, \oc8051_gm_cxrom_1.cell2.data [0], _12493_);
  and (_12599_, _10250_, _10249_);
  nor (_10251_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10252_, \oc8051_gm_cxrom_1.cell2.data [1], _10241_);
  nor (_10253_, _10252_, _10251_);
  or (_10254_, _10253_, rst);
  or (_10255_, \oc8051_gm_cxrom_1.cell2.data [1], _12493_);
  and (_12602_, _10255_, _10254_);
  nor (_10256_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10257_, \oc8051_gm_cxrom_1.cell2.data [2], _10241_);
  nor (_10258_, _10257_, _10256_);
  or (_10259_, _10258_, rst);
  or (_10260_, \oc8051_gm_cxrom_1.cell2.data [2], _12493_);
  and (_12606_, _10260_, _10259_);
  nor (_10261_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10262_, \oc8051_gm_cxrom_1.cell2.data [3], _10241_);
  nor (_10263_, _10262_, _10261_);
  or (_10264_, _10263_, rst);
  or (_10265_, \oc8051_gm_cxrom_1.cell2.data [3], _12493_);
  and (_00012_, _10265_, _10264_);
  nor (_10266_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10267_, \oc8051_gm_cxrom_1.cell2.data [4], _10241_);
  nor (_10268_, _10267_, _10266_);
  or (_10269_, _10268_, rst);
  or (_10270_, \oc8051_gm_cxrom_1.cell2.data [4], _12493_);
  and (_00016_, _10270_, _10269_);
  nor (_10271_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10272_, \oc8051_gm_cxrom_1.cell2.data [5], _10241_);
  nor (_10273_, _10272_, _10271_);
  or (_10274_, _10273_, rst);
  or (_10275_, \oc8051_gm_cxrom_1.cell2.data [5], _12493_);
  and (_00020_, _10275_, _10274_);
  nor (_10276_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  nor (_10277_, \oc8051_gm_cxrom_1.cell2.data [6], _10241_);
  nor (_10278_, _10277_, _10276_);
  or (_10279_, _10278_, rst);
  or (_10280_, \oc8051_gm_cxrom_1.cell2.data [6], _12493_);
  and (_00024_, _10280_, _10279_);
  nor (_10281_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_10282_, \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10283_, _10282_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nor (_10284_, _10283_, _10281_);
  or (_10285_, _10284_, rst);
  or (_10286_, \oc8051_gm_cxrom_1.cell3.data [7], _12493_);
  and (_00045_, _10286_, _10285_);
  nor (_10287_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10288_, \oc8051_gm_cxrom_1.cell3.data [0], _10282_);
  nor (_10289_, _10288_, _10287_);
  or (_10290_, _10289_, rst);
  or (_10291_, \oc8051_gm_cxrom_1.cell3.data [0], _12493_);
  and (_00052_, _10291_, _10290_);
  nor (_10292_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10293_, \oc8051_gm_cxrom_1.cell3.data [1], _10282_);
  nor (_10294_, _10293_, _10292_);
  or (_10295_, _10294_, rst);
  or (_10296_, \oc8051_gm_cxrom_1.cell3.data [1], _12493_);
  and (_00056_, _10296_, _10295_);
  nor (_10297_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10298_, \oc8051_gm_cxrom_1.cell3.data [2], _10282_);
  nor (_10299_, _10298_, _10297_);
  or (_10300_, _10299_, rst);
  or (_10301_, \oc8051_gm_cxrom_1.cell3.data [2], _12493_);
  and (_00060_, _10301_, _10300_);
  nor (_10302_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10303_, \oc8051_gm_cxrom_1.cell3.data [3], _10282_);
  nor (_10304_, _10303_, _10302_);
  or (_10305_, _10304_, rst);
  or (_10306_, \oc8051_gm_cxrom_1.cell3.data [3], _12493_);
  and (_00064_, _10306_, _10305_);
  nor (_10307_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10308_, \oc8051_gm_cxrom_1.cell3.data [4], _10282_);
  nor (_10309_, _10308_, _10307_);
  or (_10310_, _10309_, rst);
  or (_10311_, \oc8051_gm_cxrom_1.cell3.data [4], _12493_);
  and (_00067_, _10311_, _10310_);
  nor (_10312_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10313_, \oc8051_gm_cxrom_1.cell3.data [5], _10282_);
  nor (_10314_, _10313_, _10312_);
  or (_10315_, _10314_, rst);
  or (_10316_, \oc8051_gm_cxrom_1.cell3.data [5], _12493_);
  and (_00071_, _10316_, _10315_);
  nor (_10317_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  nor (_10318_, \oc8051_gm_cxrom_1.cell3.data [6], _10282_);
  nor (_10319_, _10318_, _10317_);
  or (_10320_, _10319_, rst);
  or (_10321_, \oc8051_gm_cxrom_1.cell3.data [6], _12493_);
  and (_00075_, _10321_, _10320_);
  nor (_10322_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_10323_, \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10324_, _10323_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nor (_10325_, _10324_, _10322_);
  or (_10326_, _10325_, rst);
  or (_10327_, \oc8051_gm_cxrom_1.cell4.data [7], _12493_);
  and (_00096_, _10327_, _10326_);
  nor (_10328_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10329_, \oc8051_gm_cxrom_1.cell4.data [0], _10323_);
  nor (_10330_, _10329_, _10328_);
  or (_10331_, _10330_, rst);
  or (_10332_, \oc8051_gm_cxrom_1.cell4.data [0], _12493_);
  and (_00103_, _10332_, _10331_);
  nor (_10333_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10334_, \oc8051_gm_cxrom_1.cell4.data [1], _10323_);
  nor (_10335_, _10334_, _10333_);
  or (_10336_, _10335_, rst);
  or (_10337_, \oc8051_gm_cxrom_1.cell4.data [1], _12493_);
  and (_00107_, _10337_, _10336_);
  nor (_10338_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10339_, \oc8051_gm_cxrom_1.cell4.data [2], _10323_);
  nor (_10340_, _10339_, _10338_);
  or (_10341_, _10340_, rst);
  or (_10342_, \oc8051_gm_cxrom_1.cell4.data [2], _12493_);
  and (_00111_, _10342_, _10341_);
  nor (_10343_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10344_, \oc8051_gm_cxrom_1.cell4.data [3], _10323_);
  nor (_10345_, _10344_, _10343_);
  or (_10346_, _10345_, rst);
  or (_10347_, \oc8051_gm_cxrom_1.cell4.data [3], _12493_);
  and (_00115_, _10347_, _10346_);
  nor (_10348_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10349_, \oc8051_gm_cxrom_1.cell4.data [4], _10323_);
  nor (_10350_, _10349_, _10348_);
  or (_10351_, _10350_, rst);
  or (_10352_, \oc8051_gm_cxrom_1.cell4.data [4], _12493_);
  and (_00119_, _10352_, _10351_);
  nor (_10353_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10354_, \oc8051_gm_cxrom_1.cell4.data [5], _10323_);
  nor (_10355_, _10354_, _10353_);
  or (_10356_, _10355_, rst);
  or (_10357_, \oc8051_gm_cxrom_1.cell4.data [5], _12493_);
  and (_00123_, _10357_, _10356_);
  nor (_10358_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  nor (_10359_, \oc8051_gm_cxrom_1.cell4.data [6], _10323_);
  nor (_10360_, _10359_, _10358_);
  or (_10361_, _10360_, rst);
  or (_10362_, \oc8051_gm_cxrom_1.cell4.data [6], _12493_);
  and (_00127_, _10362_, _10361_);
  nor (_10363_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_10364_, \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10365_, _10364_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nor (_10366_, _10365_, _10363_);
  or (_10367_, _10366_, rst);
  or (_10368_, \oc8051_gm_cxrom_1.cell5.data [7], _12493_);
  and (_00148_, _10368_, _10367_);
  nor (_10369_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10370_, \oc8051_gm_cxrom_1.cell5.data [0], _10364_);
  nor (_10371_, _10370_, _10369_);
  or (_10372_, _10371_, rst);
  or (_10373_, \oc8051_gm_cxrom_1.cell5.data [0], _12493_);
  and (_00155_, _10373_, _10372_);
  nor (_10375_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10376_, \oc8051_gm_cxrom_1.cell5.data [1], _10364_);
  nor (_10377_, _10376_, _10375_);
  or (_10378_, _10377_, rst);
  or (_10379_, \oc8051_gm_cxrom_1.cell5.data [1], _12493_);
  and (_00158_, _10379_, _10378_);
  nor (_10381_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10382_, \oc8051_gm_cxrom_1.cell5.data [2], _10364_);
  nor (_10383_, _10382_, _10381_);
  or (_10384_, _10383_, rst);
  or (_10386_, \oc8051_gm_cxrom_1.cell5.data [2], _12493_);
  and (_00162_, _10386_, _10384_);
  nor (_10387_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10388_, \oc8051_gm_cxrom_1.cell5.data [3], _10364_);
  nor (_10389_, _10388_, _10387_);
  or (_10391_, _10389_, rst);
  or (_10392_, \oc8051_gm_cxrom_1.cell5.data [3], _12493_);
  and (_00166_, _10392_, _10391_);
  nor (_10393_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10394_, \oc8051_gm_cxrom_1.cell5.data [4], _10364_);
  nor (_10396_, _10394_, _10393_);
  or (_10397_, _10396_, rst);
  or (_10398_, \oc8051_gm_cxrom_1.cell5.data [4], _12493_);
  and (_00170_, _10398_, _10397_);
  nor (_10399_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10401_, \oc8051_gm_cxrom_1.cell5.data [5], _10364_);
  nor (_10402_, _10401_, _10399_);
  or (_10403_, _10402_, rst);
  or (_10404_, \oc8051_gm_cxrom_1.cell5.data [5], _12493_);
  and (_00174_, _10404_, _10403_);
  nor (_10406_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  nor (_10407_, \oc8051_gm_cxrom_1.cell5.data [6], _10364_);
  nor (_10409_, _10407_, _10406_);
  or (_10410_, _10409_, rst);
  or (_10411_, \oc8051_gm_cxrom_1.cell5.data [6], _12493_);
  and (_00178_, _10411_, _10410_);
  nor (_10412_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_10413_, \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10414_, _10413_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nor (_10416_, _10414_, _10412_);
  or (_10417_, _10416_, rst);
  or (_10418_, \oc8051_gm_cxrom_1.cell6.data [7], _12493_);
  and (_00198_, _10418_, _10417_);
  nor (_10420_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10421_, \oc8051_gm_cxrom_1.cell6.data [0], _10413_);
  nor (_10423_, _10421_, _10420_);
  or (_10424_, _10423_, rst);
  or (_10425_, \oc8051_gm_cxrom_1.cell6.data [0], _12493_);
  and (_00204_, _10425_, _10424_);
  nor (_10427_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10428_, \oc8051_gm_cxrom_1.cell6.data [1], _10413_);
  nor (_10430_, _10428_, _10427_);
  or (_10431_, _10430_, rst);
  or (_10432_, \oc8051_gm_cxrom_1.cell6.data [1], _12493_);
  and (_00208_, _10432_, _10431_);
  nor (_10434_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10435_, \oc8051_gm_cxrom_1.cell6.data [2], _10413_);
  nor (_10437_, _10435_, _10434_);
  or (_10438_, _10437_, rst);
  or (_10440_, \oc8051_gm_cxrom_1.cell6.data [2], _12493_);
  and (_00212_, _10440_, _10438_);
  nor (_10441_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10442_, \oc8051_gm_cxrom_1.cell6.data [3], _10413_);
  nor (_10443_, _10442_, _10441_);
  or (_10444_, _10443_, rst);
  or (_10445_, \oc8051_gm_cxrom_1.cell6.data [3], _12493_);
  and (_00215_, _10445_, _10444_);
  nor (_10447_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10448_, \oc8051_gm_cxrom_1.cell6.data [4], _10413_);
  nor (_10450_, _10448_, _10447_);
  or (_10451_, _10450_, rst);
  or (_10452_, \oc8051_gm_cxrom_1.cell6.data [4], _12493_);
  and (_00219_, _10452_, _10451_);
  nor (_10454_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10455_, \oc8051_gm_cxrom_1.cell6.data [5], _10413_);
  nor (_10457_, _10455_, _10454_);
  or (_10458_, _10457_, rst);
  or (_10459_, \oc8051_gm_cxrom_1.cell6.data [5], _12493_);
  and (_00222_, _10459_, _10458_);
  nor (_10461_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  nor (_10462_, \oc8051_gm_cxrom_1.cell6.data [6], _10413_);
  nor (_10464_, _10462_, _10461_);
  or (_10465_, _10464_, rst);
  or (_10466_, \oc8051_gm_cxrom_1.cell6.data [6], _12493_);
  and (_00226_, _10466_, _10465_);
  nor (_10468_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_10470_, \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10471_, _10470_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nor (_10472_, _10471_, _10468_);
  or (_10473_, _10472_, rst);
  or (_10474_, \oc8051_gm_cxrom_1.cell7.data [7], _12493_);
  and (_00245_, _10474_, _10473_);
  nor (_10476_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10477_, \oc8051_gm_cxrom_1.cell7.data [0], _10470_);
  nor (_10479_, _10477_, _10476_);
  or (_10480_, _10479_, rst);
  or (_10481_, \oc8051_gm_cxrom_1.cell7.data [0], _12493_);
  and (_00252_, _10481_, _10480_);
  nor (_10483_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10484_, \oc8051_gm_cxrom_1.cell7.data [1], _10470_);
  nor (_10486_, _10484_, _10483_);
  or (_10487_, _10486_, rst);
  or (_10488_, \oc8051_gm_cxrom_1.cell7.data [1], _12493_);
  and (_00256_, _10488_, _10487_);
  nor (_10490_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10491_, \oc8051_gm_cxrom_1.cell7.data [2], _10470_);
  nor (_10493_, _10491_, _10490_);
  or (_10494_, _10493_, rst);
  or (_10495_, \oc8051_gm_cxrom_1.cell7.data [2], _12493_);
  and (_00259_, _10495_, _10494_);
  nor (_10497_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10499_, \oc8051_gm_cxrom_1.cell7.data [3], _10470_);
  nor (_10500_, _10499_, _10497_);
  or (_10501_, _10500_, rst);
  or (_10502_, \oc8051_gm_cxrom_1.cell7.data [3], _12493_);
  and (_00263_, _10502_, _10501_);
  nor (_10503_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10504_, \oc8051_gm_cxrom_1.cell7.data [4], _10470_);
  nor (_10506_, _10504_, _10503_);
  or (_10507_, _10506_, rst);
  or (_10508_, \oc8051_gm_cxrom_1.cell7.data [4], _12493_);
  and (_00266_, _10508_, _10507_);
  nor (_10510_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10511_, \oc8051_gm_cxrom_1.cell7.data [5], _10470_);
  nor (_10513_, _10511_, _10510_);
  or (_10514_, _10513_, rst);
  or (_10515_, \oc8051_gm_cxrom_1.cell7.data [5], _12493_);
  and (_00270_, _10515_, _10514_);
  nor (_10517_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  nor (_10518_, \oc8051_gm_cxrom_1.cell7.data [6], _10470_);
  nor (_10520_, _10518_, _10517_);
  or (_10521_, _10520_, rst);
  or (_10522_, \oc8051_gm_cxrom_1.cell7.data [6], _12493_);
  and (_00274_, _10522_, _10521_);
  nor (_10524_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_10525_, \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10527_, _10525_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nor (_10528_, _10527_, _10524_);
  or (_10530_, _10528_, rst);
  or (_10531_, \oc8051_gm_cxrom_1.cell8.data [7], _12493_);
  and (_00293_, _10531_, _10530_);
  nor (_10532_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10534_, \oc8051_gm_cxrom_1.cell8.data [0], _10525_);
  nor (_10535_, _10534_, _10532_);
  or (_10536_, _10535_, rst);
  or (_10538_, \oc8051_gm_cxrom_1.cell8.data [0], _12493_);
  and (_00299_, _10538_, _10536_);
  nor (_10539_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10541_, \oc8051_gm_cxrom_1.cell8.data [1], _10525_);
  nor (_10542_, _10541_, _10539_);
  or (_10543_, _10542_, rst);
  or (_10545_, \oc8051_gm_cxrom_1.cell8.data [1], _12493_);
  and (_00303_, _10545_, _10543_);
  nor (_10546_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10548_, \oc8051_gm_cxrom_1.cell8.data [2], _10525_);
  nor (_10549_, _10548_, _10546_);
  or (_10550_, _10549_, rst);
  or (_10552_, \oc8051_gm_cxrom_1.cell8.data [2], _12493_);
  and (_00307_, _10552_, _10550_);
  nor (_10553_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10555_, \oc8051_gm_cxrom_1.cell8.data [3], _10525_);
  nor (_10556_, _10555_, _10553_);
  or (_10558_, _10556_, rst);
  or (_10559_, \oc8051_gm_cxrom_1.cell8.data [3], _12493_);
  and (_00310_, _10559_, _10558_);
  nor (_10560_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10562_, \oc8051_gm_cxrom_1.cell8.data [4], _10525_);
  nor (_10563_, _10562_, _10560_);
  or (_10564_, _10563_, rst);
  or (_10566_, \oc8051_gm_cxrom_1.cell8.data [4], _12493_);
  and (_00314_, _10566_, _10564_);
  nor (_10567_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10569_, \oc8051_gm_cxrom_1.cell8.data [5], _10525_);
  nor (_10570_, _10569_, _10567_);
  or (_10571_, _10570_, rst);
  or (_10573_, \oc8051_gm_cxrom_1.cell8.data [5], _12493_);
  and (_00318_, _10573_, _10571_);
  nor (_10574_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  nor (_10576_, \oc8051_gm_cxrom_1.cell8.data [6], _10525_);
  nor (_10577_, _10576_, _10574_);
  or (_10578_, _10577_, rst);
  or (_10580_, \oc8051_gm_cxrom_1.cell8.data [6], _12493_);
  and (_00319_, _10580_, _10578_);
  nor (_10581_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_10583_, \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10584_, _10583_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nor (_10586_, _10584_, _10581_);
  or (_10587_, _10586_, rst);
  or (_10588_, \oc8051_gm_cxrom_1.cell9.data [7], _12493_);
  and (_00333_, _10588_, _10587_);
  nor (_10590_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10591_, \oc8051_gm_cxrom_1.cell9.data [0], _10583_);
  nor (_10592_, _10591_, _10590_);
  or (_10594_, _10592_, rst);
  or (_10595_, \oc8051_gm_cxrom_1.cell9.data [0], _12493_);
  and (_00339_, _10595_, _10594_);
  nor (_10597_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10598_, \oc8051_gm_cxrom_1.cell9.data [1], _10583_);
  nor (_10599_, _10598_, _10597_);
  or (_10601_, _10599_, rst);
  or (_10602_, \oc8051_gm_cxrom_1.cell9.data [1], _12493_);
  and (_00342_, _10602_, _10601_);
  nor (_10604_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10605_, \oc8051_gm_cxrom_1.cell9.data [2], _10583_);
  nor (_10606_, _10605_, _10604_);
  or (_10608_, _10606_, rst);
  or (_10609_, \oc8051_gm_cxrom_1.cell9.data [2], _12493_);
  and (_00346_, _10609_, _10608_);
  nor (_10611_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10612_, \oc8051_gm_cxrom_1.cell9.data [3], _10583_);
  nor (_10614_, _10612_, _10611_);
  or (_10615_, _10614_, rst);
  or (_10616_, \oc8051_gm_cxrom_1.cell9.data [3], _12493_);
  and (_00349_, _10616_, _10615_);
  nor (_10617_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10618_, \oc8051_gm_cxrom_1.cell9.data [4], _10583_);
  nor (_10619_, _10618_, _10617_);
  or (_10621_, _10619_, rst);
  or (_10622_, \oc8051_gm_cxrom_1.cell9.data [4], _12493_);
  and (_00352_, _10622_, _10621_);
  nor (_10624_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10625_, \oc8051_gm_cxrom_1.cell9.data [5], _10583_);
  nor (_10626_, _10625_, _10624_);
  or (_10628_, _10626_, rst);
  or (_10629_, \oc8051_gm_cxrom_1.cell9.data [5], _12493_);
  and (_00356_, _10629_, _10628_);
  nor (_10631_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  nor (_10632_, \oc8051_gm_cxrom_1.cell9.data [6], _10583_);
  nor (_10633_, _10632_, _10631_);
  or (_10635_, _10633_, rst);
  or (_10636_, \oc8051_gm_cxrom_1.cell9.data [6], _12493_);
  and (_00359_, _10636_, _10635_);
  nor (_10638_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_10639_, \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10640_, _10639_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nor (_10642_, _10640_, _10638_);
  or (_10643_, _10642_, rst);
  or (_10645_, \oc8051_gm_cxrom_1.cell10.data [7], _12493_);
  and (_00374_, _10645_, _10643_);
  nor (_10646_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10647_, \oc8051_gm_cxrom_1.cell10.data [0], _10639_);
  nor (_10649_, _10647_, _10646_);
  or (_10650_, _10649_, rst);
  or (_10651_, \oc8051_gm_cxrom_1.cell10.data [0], _12493_);
  and (_00379_, _10651_, _10650_);
  nor (_10653_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10654_, \oc8051_gm_cxrom_1.cell10.data [1], _10639_);
  nor (_10656_, _10654_, _10653_);
  or (_10657_, _10656_, rst);
  or (_10658_, \oc8051_gm_cxrom_1.cell10.data [1], _12493_);
  and (_00383_, _10658_, _10657_);
  nor (_10660_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10661_, \oc8051_gm_cxrom_1.cell10.data [2], _10639_);
  nor (_10663_, _10661_, _10660_);
  or (_10664_, _10663_, rst);
  or (_10665_, \oc8051_gm_cxrom_1.cell10.data [2], _12493_);
  and (_00386_, _10665_, _10664_);
  nor (_10667_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10668_, \oc8051_gm_cxrom_1.cell10.data [3], _10639_);
  nor (_10670_, _10668_, _10667_);
  or (_10671_, _10670_, rst);
  or (_10673_, \oc8051_gm_cxrom_1.cell10.data [3], _12493_);
  and (_00389_, _10673_, _10671_);
  nor (_10674_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10675_, \oc8051_gm_cxrom_1.cell10.data [4], _10639_);
  nor (_10677_, _10675_, _10674_);
  or (_10678_, _10677_, rst);
  or (_10679_, \oc8051_gm_cxrom_1.cell10.data [4], _12493_);
  and (_00392_, _10679_, _10678_);
  nor (_10681_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10682_, \oc8051_gm_cxrom_1.cell10.data [5], _10639_);
  nor (_10684_, _10682_, _10681_);
  or (_10685_, _10684_, rst);
  or (_10686_, \oc8051_gm_cxrom_1.cell10.data [5], _12493_);
  and (_00396_, _10686_, _10685_);
  nor (_10688_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  nor (_10689_, \oc8051_gm_cxrom_1.cell10.data [6], _10639_);
  nor (_10691_, _10689_, _10688_);
  or (_10692_, _10691_, rst);
  or (_10693_, \oc8051_gm_cxrom_1.cell10.data [6], _12493_);
  and (_00399_, _10693_, _10692_);
  nor (_10695_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_10696_, \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10698_, _10696_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nor (_10699_, _10698_, _10695_);
  or (_10701_, _10699_, rst);
  or (_10702_, \oc8051_gm_cxrom_1.cell11.data [7], _12493_);
  and (_00416_, _10702_, _10701_);
  nor (_10703_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10705_, \oc8051_gm_cxrom_1.cell11.data [0], _10696_);
  nor (_10706_, _10705_, _10703_);
  or (_10707_, _10706_, rst);
  or (_10709_, \oc8051_gm_cxrom_1.cell11.data [0], _12493_);
  and (_00421_, _10709_, _10707_);
  nor (_10710_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10712_, \oc8051_gm_cxrom_1.cell11.data [1], _10696_);
  nor (_10713_, _10712_, _10710_);
  or (_10714_, _10713_, rst);
  or (_10716_, \oc8051_gm_cxrom_1.cell11.data [1], _12493_);
  and (_00425_, _10716_, _10714_);
  nor (_10717_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10719_, \oc8051_gm_cxrom_1.cell11.data [2], _10696_);
  nor (_10720_, _10719_, _10717_);
  or (_10721_, _10720_, rst);
  or (_10723_, \oc8051_gm_cxrom_1.cell11.data [2], _12493_);
  and (_00428_, _10723_, _10721_);
  nor (_10724_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10726_, \oc8051_gm_cxrom_1.cell11.data [3], _10696_);
  nor (_10727_, _10726_, _10724_);
  or (_10729_, _10727_, rst);
  or (_10730_, \oc8051_gm_cxrom_1.cell11.data [3], _12493_);
  and (_00431_, _10730_, _10729_);
  nor (_10731_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10732_, \oc8051_gm_cxrom_1.cell11.data [4], _10696_);
  nor (_10734_, _10732_, _10731_);
  or (_10735_, _10734_, rst);
  or (_10736_, \oc8051_gm_cxrom_1.cell11.data [4], _12493_);
  and (_00434_, _10736_, _10735_);
  nor (_10738_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10739_, \oc8051_gm_cxrom_1.cell11.data [5], _10696_);
  nor (_10741_, _10739_, _10738_);
  or (_10742_, _10741_, rst);
  or (_10743_, \oc8051_gm_cxrom_1.cell11.data [5], _12493_);
  and (_00438_, _10743_, _10742_);
  nor (_10745_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  nor (_10746_, \oc8051_gm_cxrom_1.cell11.data [6], _10696_);
  nor (_10748_, _10746_, _10745_);
  or (_10749_, _10748_, rst);
  or (_10750_, \oc8051_gm_cxrom_1.cell11.data [6], _12493_);
  and (_00441_, _10750_, _10749_);
  nor (_10752_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_10753_, \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10755_, _10753_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nor (_10756_, _10755_, _10752_);
  or (_10758_, _10756_, rst);
  or (_10759_, \oc8051_gm_cxrom_1.cell12.data [7], _12493_);
  and (_00458_, _10759_, _10758_);
  nor (_10760_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10762_, \oc8051_gm_cxrom_1.cell12.data [0], _10753_);
  nor (_10763_, _10762_, _10760_);
  or (_10764_, _10763_, rst);
  or (_10766_, \oc8051_gm_cxrom_1.cell12.data [0], _12493_);
  and (_00463_, _10766_, _10764_);
  nor (_10767_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10769_, \oc8051_gm_cxrom_1.cell12.data [1], _10753_);
  nor (_10770_, _10769_, _10767_);
  or (_10771_, _10770_, rst);
  or (_10773_, \oc8051_gm_cxrom_1.cell12.data [1], _12493_);
  and (_00467_, _10773_, _10771_);
  nor (_10774_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10776_, \oc8051_gm_cxrom_1.cell12.data [2], _10753_);
  nor (_10777_, _10776_, _10774_);
  or (_10778_, _10777_, rst);
  or (_10780_, \oc8051_gm_cxrom_1.cell12.data [2], _12493_);
  and (_00470_, _10780_, _10778_);
  nor (_10781_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10783_, \oc8051_gm_cxrom_1.cell12.data [3], _10753_);
  nor (_10784_, _10783_, _10781_);
  or (_10786_, _10784_, rst);
  or (_10787_, \oc8051_gm_cxrom_1.cell12.data [3], _12493_);
  and (_00473_, _10787_, _10786_);
  nor (_10788_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10790_, \oc8051_gm_cxrom_1.cell12.data [4], _10753_);
  nor (_10791_, _10790_, _10788_);
  or (_10792_, _10791_, rst);
  or (_10794_, \oc8051_gm_cxrom_1.cell12.data [4], _12493_);
  and (_00476_, _10794_, _10792_);
  nor (_10795_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10797_, \oc8051_gm_cxrom_1.cell12.data [5], _10753_);
  nor (_10798_, _10797_, _10795_);
  or (_10799_, _10798_, rst);
  or (_10801_, \oc8051_gm_cxrom_1.cell12.data [5], _12493_);
  and (_00480_, _10801_, _10799_);
  nor (_10802_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  nor (_10804_, \oc8051_gm_cxrom_1.cell12.data [6], _10753_);
  nor (_10805_, _10804_, _10802_);
  or (_10806_, _10805_, rst);
  or (_10808_, \oc8051_gm_cxrom_1.cell12.data [6], _12493_);
  and (_00483_, _10808_, _10806_);
  nor (_10809_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_10811_, \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10812_, _10811_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nor (_10814_, _10812_, _10809_);
  or (_10815_, _10814_, rst);
  or (_10816_, \oc8051_gm_cxrom_1.cell13.data [7], _12493_);
  and (_00502_, _10816_, _10815_);
  nor (_10818_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10819_, \oc8051_gm_cxrom_1.cell13.data [0], _10811_);
  nor (_10820_, _10819_, _10818_);
  or (_10822_, _10820_, rst);
  or (_10823_, \oc8051_gm_cxrom_1.cell13.data [0], _12493_);
  and (_00508_, _10823_, _10822_);
  nor (_10825_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10826_, \oc8051_gm_cxrom_1.cell13.data [1], _10811_);
  nor (_10827_, _10826_, _10825_);
  or (_10829_, _10827_, rst);
  or (_10830_, \oc8051_gm_cxrom_1.cell13.data [1], _12493_);
  and (_00511_, _10830_, _10829_);
  nor (_10832_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10833_, \oc8051_gm_cxrom_1.cell13.data [2], _10811_);
  nor (_10834_, _10833_, _10832_);
  or (_10836_, _10834_, rst);
  or (_10837_, \oc8051_gm_cxrom_1.cell13.data [2], _12493_);
  and (_00515_, _10837_, _10836_);
  nor (_10839_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10840_, \oc8051_gm_cxrom_1.cell13.data [3], _10811_);
  nor (_10841_, _10840_, _10839_);
  or (_10842_, _10841_, rst);
  or (_10843_, \oc8051_gm_cxrom_1.cell13.data [3], _12493_);
  and (_00518_, _10843_, _10842_);
  nor (_10844_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10845_, \oc8051_gm_cxrom_1.cell13.data [4], _10811_);
  nor (_10846_, _10845_, _10844_);
  or (_10847_, _10846_, rst);
  or (_10848_, \oc8051_gm_cxrom_1.cell13.data [4], _12493_);
  and (_00522_, _10848_, _10847_);
  nor (_10849_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10850_, \oc8051_gm_cxrom_1.cell13.data [5], _10811_);
  nor (_10851_, _10850_, _10849_);
  or (_10852_, _10851_, rst);
  or (_10853_, \oc8051_gm_cxrom_1.cell13.data [5], _12493_);
  and (_00525_, _10853_, _10852_);
  nor (_10854_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  nor (_10855_, \oc8051_gm_cxrom_1.cell13.data [6], _10811_);
  nor (_10856_, _10855_, _10854_);
  or (_10857_, _10856_, rst);
  or (_10858_, \oc8051_gm_cxrom_1.cell13.data [6], _12493_);
  and (_00529_, _10858_, _10857_);
  nor (_10859_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_10860_, \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10861_, _10860_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nor (_10862_, _10861_, _10859_);
  or (_10863_, _10862_, rst);
  or (_10864_, \oc8051_gm_cxrom_1.cell14.data [7], _12493_);
  and (_12609_[7], _10864_, _10863_);
  nor (_10865_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10866_, \oc8051_gm_cxrom_1.cell14.data [0], _10860_);
  nor (_10867_, _10866_, _10865_);
  or (_10868_, _10867_, rst);
  or (_10869_, \oc8051_gm_cxrom_1.cell14.data [0], _12493_);
  and (_12609_[0], _10869_, _10868_);
  nor (_10870_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10871_, \oc8051_gm_cxrom_1.cell14.data [1], _10860_);
  nor (_10872_, _10871_, _10870_);
  or (_10873_, _10872_, rst);
  or (_10874_, \oc8051_gm_cxrom_1.cell14.data [1], _12493_);
  and (_12609_[1], _10874_, _10873_);
  nor (_10875_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10876_, \oc8051_gm_cxrom_1.cell14.data [2], _10860_);
  nor (_10877_, _10876_, _10875_);
  or (_10878_, _10877_, rst);
  or (_10879_, \oc8051_gm_cxrom_1.cell14.data [2], _12493_);
  and (_12609_[2], _10879_, _10878_);
  nor (_10880_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10881_, \oc8051_gm_cxrom_1.cell14.data [3], _10860_);
  nor (_10882_, _10881_, _10880_);
  or (_10883_, _10882_, rst);
  or (_10884_, \oc8051_gm_cxrom_1.cell14.data [3], _12493_);
  and (_12609_[3], _10884_, _10883_);
  nor (_10885_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10886_, \oc8051_gm_cxrom_1.cell14.data [4], _10860_);
  nor (_10887_, _10886_, _10885_);
  or (_10888_, _10887_, rst);
  or (_10889_, \oc8051_gm_cxrom_1.cell14.data [4], _12493_);
  and (_12609_[4], _10889_, _10888_);
  nor (_10890_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10891_, \oc8051_gm_cxrom_1.cell14.data [5], _10860_);
  nor (_10892_, _10891_, _10890_);
  or (_10893_, _10892_, rst);
  or (_10894_, \oc8051_gm_cxrom_1.cell14.data [5], _12493_);
  and (_12609_[5], _10894_, _10893_);
  nor (_10895_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  nor (_10896_, \oc8051_gm_cxrom_1.cell14.data [6], _10860_);
  nor (_10897_, _10896_, _10895_);
  or (_10898_, _10897_, rst);
  or (_10899_, \oc8051_gm_cxrom_1.cell14.data [6], _12493_);
  and (_12609_[6], _10899_, _10898_);
  nor (_10900_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_10901_, \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10902_, _10901_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nor (_10903_, _10902_, _10900_);
  or (_10904_, _10903_, rst);
  or (_10905_, \oc8051_gm_cxrom_1.cell15.data [7], _12493_);
  and (_12610_[7], _10905_, _10904_);
  nor (_10906_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10907_, \oc8051_gm_cxrom_1.cell15.data [0], _10901_);
  nor (_10908_, _10907_, _10906_);
  or (_10909_, _10908_, rst);
  or (_10910_, \oc8051_gm_cxrom_1.cell15.data [0], _12493_);
  and (_12610_[0], _10910_, _10909_);
  nor (_10911_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10912_, \oc8051_gm_cxrom_1.cell15.data [1], _10901_);
  nor (_10913_, _10912_, _10911_);
  or (_10914_, _10913_, rst);
  or (_10915_, \oc8051_gm_cxrom_1.cell15.data [1], _12493_);
  and (_12610_[1], _10915_, _10914_);
  nor (_10916_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10917_, \oc8051_gm_cxrom_1.cell15.data [2], _10901_);
  nor (_10918_, _10917_, _10916_);
  or (_10919_, _10918_, rst);
  or (_10920_, \oc8051_gm_cxrom_1.cell15.data [2], _12493_);
  and (_12610_[2], _10920_, _10919_);
  nor (_10921_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10922_, \oc8051_gm_cxrom_1.cell15.data [3], _10901_);
  nor (_10923_, _10922_, _10921_);
  or (_10924_, _10923_, rst);
  or (_10925_, \oc8051_gm_cxrom_1.cell15.data [3], _12493_);
  and (_12610_[3], _10925_, _10924_);
  nor (_10926_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10927_, \oc8051_gm_cxrom_1.cell15.data [4], _10901_);
  nor (_10928_, _10927_, _10926_);
  or (_10929_, _10928_, rst);
  or (_10930_, \oc8051_gm_cxrom_1.cell15.data [4], _12493_);
  and (_12610_[4], _10930_, _10929_);
  nor (_10931_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10932_, \oc8051_gm_cxrom_1.cell15.data [5], _10901_);
  nor (_10933_, _10932_, _10931_);
  or (_10934_, _10933_, rst);
  or (_10935_, \oc8051_gm_cxrom_1.cell15.data [5], _12493_);
  and (_12610_[5], _10935_, _10934_);
  nor (_10936_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  nor (_10937_, \oc8051_gm_cxrom_1.cell15.data [6], _10901_);
  nor (_10938_, _10937_, _10936_);
  or (_10939_, _10938_, rst);
  or (_10940_, \oc8051_gm_cxrom_1.cell15.data [6], _12493_);
  and (_12610_[6], _10940_, _10939_);
  nor (_12678_[2], _07731_, rst);
  and (_10941_, _07312_, _12493_);
  nand (_10942_, _10941_, _07595_);
  nor (_10943_, _07559_, _07440_);
  or (_12679_[2], _10943_, _10942_);
  and (_10944_, _07407_, _07381_);
  and (_10945_, _10944_, _07433_);
  and (_10946_, _10945_, _07355_);
  and (_10947_, _07488_, _07462_);
  and (_10948_, _10947_, _07515_);
  and (_10949_, _10948_, _10946_);
  and (_10950_, _10949_, _07546_);
  not (_10951_, _07462_);
  and (_10952_, _07488_, _10951_);
  not (_10953_, _07546_);
  not (_10954_, _07381_);
  and (_10955_, _07407_, _10954_);
  not (_10956_, _07355_);
  nor (_10957_, _07433_, _10956_);
  and (_10958_, _10957_, _10955_);
  and (_10959_, _10958_, _10953_);
  and (_10960_, _10959_, _10952_);
  and (_10961_, _10949_, _10953_);
  or (_10962_, _10961_, _10960_);
  or (_10963_, _10962_, _10950_);
  and (_10964_, _10953_, _07515_);
  and (_10965_, _10964_, _10952_);
  and (_10966_, _10957_, _10944_);
  and (_10967_, _10966_, _10965_);
  not (_10968_, _07515_);
  and (_10969_, _10952_, _10968_);
  and (_10970_, _07546_, _07433_);
  and (_10971_, _10970_, _10955_);
  not (_10972_, _07407_);
  and (_10973_, _07546_, _10972_);
  or (_10974_, _10973_, _10971_);
  and (_10975_, _10974_, _10969_);
  nor (_10976_, _10975_, _10967_);
  nor (_10977_, _10953_, _07515_);
  nor (_10978_, _10977_, _10964_);
  and (_10979_, _10978_, _10947_);
  and (_10980_, _10979_, _10966_);
  and (_10981_, _07546_, _07515_);
  nor (_10982_, _07488_, _07462_);
  and (_10983_, _10982_, _10981_);
  not (_10984_, _07433_);
  and (_10985_, _10955_, _10984_);
  and (_10986_, _10985_, _10956_);
  and (_10987_, _10986_, _10983_);
  nor (_10988_, _10987_, _10980_);
  nand (_10989_, _10988_, _10976_);
  and (_10990_, _10947_, _10968_);
  and (_10991_, _10990_, _10946_);
  and (_10992_, _10952_, _07515_);
  and (_10993_, _10945_, _10956_);
  and (_10994_, _10993_, _10992_);
  or (_10995_, _10994_, _10991_);
  and (_10996_, _10977_, _10952_);
  and (_10997_, _10996_, _10985_);
  nor (_10998_, _07546_, _07515_);
  and (_10999_, _10982_, _10998_);
  and (_11000_, _10999_, _10945_);
  or (_11001_, _11000_, _10997_);
  and (_11002_, _10982_, _10977_);
  and (_11003_, _11002_, _10945_);
  and (_11004_, _10983_, _10972_);
  or (_11005_, _11004_, _11003_);
  or (_11006_, _11005_, _11001_);
  or (_11007_, _11006_, _10995_);
  or (_11008_, _11007_, _10989_);
  and (_11009_, _10944_, _10984_);
  not (_11010_, _11009_);
  not (_11011_, _07488_);
  and (_11012_, _11011_, _07462_);
  and (_11013_, _11012_, _10998_);
  nor (_11014_, _11013_, _10956_);
  nor (_11015_, _11014_, _11010_);
  not (_11016_, _11015_);
  and (_11017_, _10977_, _10947_);
  and (_11018_, _11017_, _10966_);
  and (_11019_, _11012_, _10964_);
  and (_11020_, _11019_, _10966_);
  nor (_11021_, _11020_, _11018_);
  and (_11022_, _11021_, _11016_);
  and (_11023_, _10982_, _10968_);
  and (_11024_, _11023_, _10966_);
  and (_11025_, _11012_, _10977_);
  and (_11026_, _11025_, _10993_);
  and (_11027_, _11012_, _07546_);
  and (_11028_, _11027_, _10966_);
  or (_11029_, _11028_, _11026_);
  nor (_11030_, _11029_, _11024_);
  nand (_11031_, _11030_, _11022_);
  or (_11032_, _11031_, _11008_);
  or (_11033_, _11032_, _10963_);
  and (_11034_, _11033_, _07313_);
  not (_11035_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_11036_, _07311_, _05610_);
  and (_11037_, _11036_, _07614_);
  nor (_11038_, _11037_, _11035_);
  or (_11039_, _11038_, rst);
  or (_12680_[1], _11039_, _11034_);
  nand (_11040_, _07462_, _07307_);
  or (_11041_, _07307_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_11042_, _11041_, _12493_);
  and (_12681_[7], _11042_, _11040_);
  and (_11043_, \oc8051_top_1.oc8051_sfr1.wait_data , _12493_);
  and (_11044_, _11043_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_11045_, _07721_, _07630_);
  and (_11046_, _07602_, _07584_);
  and (_11047_, _11046_, _07551_);
  or (_11048_, _11047_, _11045_);
  and (_11049_, _07589_, _07559_);
  or (_11050_, _11049_, _07704_);
  or (_11051_, _11050_, _07679_);
  and (_11052_, _07564_, _07440_);
  and (_11053_, _07678_, _07602_);
  or (_11054_, _11053_, _11052_);
  nor (_11055_, _11054_, _11051_);
  nand (_11056_, _11055_, _07658_);
  or (_11057_, _11056_, _11048_);
  and (_11058_, _11057_, _10941_);
  or (_12682_, _11058_, _11044_);
  and (_11059_, _07551_, _07643_);
  and (_11060_, _11059_, _07562_);
  and (_11061_, _11060_, _07561_);
  or (_11062_, _11061_, _07583_);
  and (_11063_, _07553_, _07438_);
  and (_11064_, _11063_, _07678_);
  or (_11065_, _11064_, _11062_);
  and (_11066_, _07607_, _07559_);
  or (_11067_, _11066_, _07603_);
  or (_11068_, _11067_, _11065_);
  and (_11069_, _11068_, _07312_);
  and (_11070_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11071_, \oc8051_top_1.oc8051_decoder1.state [0], _05610_);
  and (_11072_, _11071_, _11035_);
  not (_11073_, _07724_);
  and (_11074_, _11073_, _11072_);
  or (_11075_, _11074_, _11070_);
  or (_11076_, _11075_, _11069_);
  and (_12683_[1], _11076_, _12493_);
  and (_11077_, _11043_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_11078_, _07721_, _07641_);
  or (_11079_, _07641_, _07564_);
  and (_11080_, _11079_, _07629_);
  or (_11081_, _11080_, _11078_);
  and (_11082_, _11063_, _07655_);
  or (_11083_, _11082_, _11081_);
  nor (_11084_, _07551_, _07412_);
  and (_11085_, _11084_, _07572_);
  and (_11086_, _11079_, _07643_);
  or (_11087_, _11086_, _11085_);
  or (_11088_, _11087_, _07575_);
  and (_11089_, _11084_, _07567_);
  and (_11090_, _07721_, _07632_);
  or (_11091_, _11090_, _11089_);
  or (_11092_, _11091_, _11067_);
  or (_11093_, _11092_, _11088_);
  or (_11094_, _11093_, _11083_);
  and (_11095_, _11094_, _10941_);
  or (_12684_[1], _11095_, _11077_);
  and (_11096_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11097_, _07694_, _07312_);
  or (_11098_, _11097_, _11096_);
  or (_11099_, _11098_, _11074_);
  and (_12685_[2], _11099_, _12493_);
  not (_11100_, _10943_);
  and (_11101_, _11100_, _07630_);
  nor (_11102_, _11101_, _11046_);
  not (_11103_, _11102_);
  and (_11104_, _11103_, _11072_);
  or (_11105_, _11104_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11106_, _07628_, _07413_);
  and (_11107_, _07572_, _07441_);
  nor (_11108_, _11107_, _11106_);
  nor (_11109_, _11108_, _07551_);
  and (_11110_, _11047_, _07727_);
  or (_11111_, _11110_, _11109_);
  and (_11112_, _11111_, _07614_);
  or (_11113_, _11112_, _11105_);
  or (_11114_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05610_);
  and (_11115_, _11114_, _12493_);
  and (_12686_[2], _11115_, _11113_);
  and (_11116_, _11043_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_11117_, _11084_, _07563_);
  or (_11118_, _11117_, _11085_);
  nor (_11119_, _07438_, _07552_);
  and (_11120_, _07412_, _07601_);
  and (_11121_, _11120_, _11119_);
  and (_11122_, _11121_, _07600_);
  or (_11123_, _07671_, _11122_);
  or (_11124_, _11123_, _11118_);
  and (_11125_, _07567_, _07441_);
  or (_11126_, _11082_, _11052_);
  or (_11127_, _11126_, _11125_);
  or (_11128_, _07678_, _07655_);
  and (_11129_, _11128_, _07554_);
  or (_11130_, _11061_, _07687_);
  or (_11131_, _11130_, _11129_);
  or (_11132_, _11131_, _11127_);
  or (_11133_, _11132_, _11124_);
  and (_11134_, _11133_, _10941_);
  or (_12687_[1], _11134_, _11116_);
  and (_11135_, _11043_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_11136_, _11064_, _07667_);
  and (_11137_, _07602_, _07494_);
  and (_11138_, _11063_, _07637_);
  or (_11139_, _11138_, _11137_);
  or (_11140_, _11139_, _11136_);
  or (_11141_, _11140_, _11087_);
  and (_11142_, _07570_, _07563_);
  or (_11143_, _07597_, _07556_);
  or (_11144_, _11143_, _11142_);
  and (_11145_, _07721_, _07662_);
  or (_11146_, _07670_, _07663_);
  or (_11147_, _11146_, _11145_);
  or (_11148_, _11147_, _11144_);
  or (_11149_, _11148_, _11141_);
  nor (_11150_, _07638_, _07573_);
  not (_11151_, _11150_);
  not (_11152_, _07676_);
  and (_11153_, _11059_, _07526_);
  or (_11154_, _11153_, _11060_);
  or (_11155_, _11154_, _11152_);
  or (_11156_, _11155_, _11151_);
  or (_11157_, _11156_, _11083_);
  or (_11158_, _11157_, _11149_);
  and (_11159_, _11158_, _10941_);
  or (_12688_[3], _11159_, _11135_);
  and (_11160_, _07554_, _07522_);
  and (_11161_, _11084_, _07584_);
  and (_11162_, _11063_, _07522_);
  or (_11163_, _11162_, _11161_);
  or (_11164_, _11163_, _11160_);
  and (_11165_, _07522_, _07643_);
  or (_11166_, _11165_, _07585_);
  or (_11167_, _11166_, _11164_);
  and (_11168_, _11063_, _07607_);
  or (_11169_, _11168_, _11073_);
  or (_11170_, _11169_, _11167_);
  and (_11171_, _11170_, _10941_);
  and (_11172_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_11173_, _11172_, _07728_);
  and (_11174_, _11173_, _12493_);
  or (_12689_[1], _11174_, _11171_);
  or (_11175_, _07690_, _07687_);
  not (_11176_, _07695_);
  or (_11177_, _11080_, _11176_);
  or (_11178_, _11177_, _11175_);
  and (_11179_, _07655_, _07441_);
  and (_11180_, _07594_, _07560_);
  and (_11181_, _11180_, _07629_);
  or (_11182_, _11181_, _07665_);
  or (_11183_, _11182_, _07663_);
  or (_11184_, _11183_, _11179_);
  nand (_11185_, _07680_, _07639_);
  or (_11186_, _11185_, _11184_);
  or (_11187_, _11186_, _11178_);
  and (_11188_, _07589_, _07643_);
  and (_11189_, _11084_, _07594_);
  or (_11190_, _11189_, _07644_);
  or (_11191_, _11190_, _11188_);
  or (_11192_, _11191_, _11062_);
  and (_11193_, _07570_, _07594_);
  or (_11194_, _11193_, _07573_);
  or (_11195_, _11194_, _07626_);
  and (_11196_, _11106_, _07560_);
  or (_11197_, _11196_, _07590_);
  or (_11198_, _11197_, _07684_);
  or (_11199_, _11198_, _11195_);
  or (_11200_, _11199_, _11192_);
  or (_11201_, _11200_, _11087_);
  or (_11202_, _11201_, _11187_);
  and (_11203_, _11202_, _07312_);
  and (_11204_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11205_, _07710_, _07706_);
  or (_11206_, _11179_, _11196_);
  and (_11207_, _11206_, _07616_);
  or (_11208_, _11207_, _11074_);
  or (_11209_, _11208_, _11205_);
  or (_11210_, _11209_, _11204_);
  or (_11211_, _11210_, _11203_);
  and (_12690_, _11211_, _12493_);
  nor (_12678_[0], _07622_, rst);
  nor (_12678_[1], _07716_, rst);
  nand (_12679_[0], _11103_, _10941_);
  nand (_11212_, _11046_, _10941_);
  or (_11213_, _10942_, _07653_);
  and (_12679_[1], _11213_, _11212_);
  or (_11214_, _10995_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_11215_, _11214_, _10960_);
  and (_11216_, _11215_, _11037_);
  nor (_11217_, _11036_, _07614_);
  or (_11218_, _11217_, rst);
  or (_12680_[0], _11218_, _11216_);
  nand (_11219_, _07355_, _07307_);
  or (_11220_, _07307_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_11221_, _11220_, _12493_);
  and (_12681_[0], _11221_, _11219_);
  not (_11222_, _07307_);
  or (_11223_, _07433_, _11222_);
  or (_11224_, _07307_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_11225_, _11224_, _12493_);
  and (_12681_[1], _11225_, _11223_);
  nand (_11226_, _07381_, _07307_);
  or (_11227_, _07307_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_11228_, _11227_, _12493_);
  and (_12681_[2], _11228_, _11226_);
  nand (_11229_, _07407_, _07307_);
  or (_11230_, _07307_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_11231_, _11230_, _12493_);
  and (_12681_[3], _11231_, _11229_);
  or (_11232_, _07546_, _11222_);
  or (_11233_, _07307_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_11234_, _11233_, _12493_);
  and (_12681_[4], _11234_, _11232_);
  nand (_11235_, _07515_, _07307_);
  or (_11236_, _07307_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_11237_, _11236_, _12493_);
  and (_12681_[5], _11237_, _11235_);
  nand (_11238_, _07488_, _07307_);
  or (_11239_, _07307_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_11240_, _11239_, _12493_);
  and (_12681_[6], _11240_, _11238_);
  or (_11241_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05610_);
  and (_11242_, _11241_, _11105_);
  and (_11243_, _11154_, _07467_);
  and (_11244_, _07595_, _07560_);
  and (_11245_, _11244_, _07721_);
  and (_11246_, _07721_, _07605_);
  and (_11247_, _11063_, _07630_);
  or (_11248_, _11247_, _11246_);
  nor (_11249_, _11248_, _11245_);
  nand (_11250_, _11249_, _07599_);
  or (_11251_, _11250_, _11243_);
  and (_11252_, _11063_, _07662_);
  or (_11253_, _11252_, _11066_);
  or (_11254_, _11253_, _11164_);
  and (_11255_, _11084_, _07579_);
  or (_11256_, _11255_, _11165_);
  or (_11257_, _07572_, _07564_);
  and (_11258_, _11257_, _07721_);
  or (_11259_, _11258_, _11256_);
  or (_11260_, _11259_, _11254_);
  and (_11261_, _07580_, _07554_);
  or (_11262_, _11261_, _11138_);
  and (_11263_, _11063_, _07580_);
  and (_11264_, _07630_, _07643_);
  or (_11265_, _11264_, _11263_);
  or (_11266_, _11265_, _11262_);
  and (_11267_, _07607_, _07554_);
  or (_11268_, _11168_, _11267_);
  or (_11269_, _11268_, _07603_);
  and (_11270_, _07637_, _07554_);
  or (_11271_, _11137_, _11270_);
  or (_11272_, _11271_, _11269_);
  or (_11273_, _11272_, _11266_);
  or (_11274_, _11273_, _11260_);
  or (_11275_, _11274_, _11251_);
  and (_11276_, _11275_, _07312_);
  or (_11277_, _11276_, _11242_);
  and (_12683_[0], _11277_, _12493_);
  and (_11278_, _11043_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_11279_, _07662_, _07637_);
  and (_11280_, _11279_, _07441_);
  or (_11281_, _11253_, _11154_);
  or (_11282_, _11281_, _11280_);
  or (_11283_, _11089_, _07571_);
  nor (_11284_, _11283_, _11090_);
  nand (_11285_, _11284_, _07688_);
  or (_11286_, _11285_, _11048_);
  not (_11287_, _07637_);
  nand (_11288_, _07581_, _11287_);
  and (_11289_, _11288_, _07721_);
  or (_11290_, _11289_, _11144_);
  or (_11291_, _11290_, _11286_);
  or (_11292_, _11291_, _11282_);
  and (_11293_, _11292_, _10941_);
  or (_12684_[0], _11293_, _11278_);
  or (_11294_, _11198_, _11188_);
  or (_11295_, _11294_, _11187_);
  and (_11296_, _11295_, _07312_);
  and (_11297_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11298_, _11297_, _11209_);
  or (_11299_, _11298_, _11296_);
  and (_12685_[0], _11299_, _12493_);
  and (_11300_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11301_, _11300_, _11208_);
  and (_11302_, _07636_, _07551_);
  or (_11303_, _11302_, _07583_);
  or (_11304_, _11303_, _11195_);
  or (_11305_, _11304_, _11109_);
  and (_11306_, _11305_, _07312_);
  or (_11307_, _11306_, _11301_);
  and (_12685_[1], _11307_, _12493_);
  or (_11308_, _11279_, _07605_);
  and (_11309_, _11308_, _07721_);
  or (_11310_, _11309_, _11109_);
  or (_11311_, _11161_, _07582_);
  or (_11312_, _11046_, _07723_);
  and (_11313_, _11162_, _07560_);
  or (_11314_, _11313_, _11263_);
  or (_11315_, _11314_, _11312_);
  or (_11316_, _11315_, _11311_);
  or (_11317_, _11316_, _11310_);
  and (_11318_, _07721_, _07678_);
  or (_11319_, _11168_, _11137_);
  or (_11320_, _11319_, _11318_);
  or (_11321_, _11320_, _11256_);
  and (_11322_, _11063_, _07666_);
  or (_11323_, _11322_, _11045_);
  or (_11324_, _11245_, _07722_);
  or (_11325_, _11324_, _11258_);
  or (_11326_, _11325_, _11323_);
  and (_11327_, _11244_, _07629_);
  and (_11328_, _11162_, _07551_);
  or (_11329_, _11328_, _07606_);
  or (_11330_, _11329_, _11327_);
  and (_11331_, _07684_, _07360_);
  or (_11332_, _11189_, _11267_);
  or (_11333_, _11332_, _11193_);
  or (_11334_, _11333_, _11331_);
  or (_11335_, _11334_, _11330_);
  or (_11336_, _11335_, _11326_);
  or (_11337_, _11336_, _11321_);
  or (_11338_, _11337_, _11317_);
  and (_11339_, _11338_, _07312_);
  and (_11340_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11341_, _11104_, _07728_);
  or (_11342_, _11341_, _11340_);
  or (_11343_, _11342_, _11339_);
  and (_12686_[0], _11343_, _12493_);
  or (_11344_, _07663_, _07638_);
  and (_11345_, _11344_, _07601_);
  and (_11346_, _07595_, _07570_);
  or (_11347_, _07723_, _11267_);
  or (_11348_, _11347_, _07684_);
  or (_11349_, _11348_, _11346_);
  or (_11350_, _11349_, _11311_);
  or (_11351_, _11350_, _11345_);
  and (_11352_, _11084_, _07595_);
  or (_11353_, _11181_, _11066_);
  nor (_11354_, _11353_, _11352_);
  nand (_11355_, _11354_, _07609_);
  or (_11356_, _11355_, _07649_);
  or (_11357_, _11356_, _11326_);
  or (_11358_, _11357_, _11321_);
  or (_11359_, _11358_, _11351_);
  and (_11360_, _11359_, _07312_);
  and (_11361_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11362_, _11361_, _11341_);
  or (_11363_, _11362_, _11360_);
  and (_12686_[1], _11363_, _12493_);
  and (_11364_, _11043_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  not (_11365_, _08861_);
  or (_11366_, _11168_, _11365_);
  and (_11367_, _07602_, _07572_);
  and (_11368_, _11367_, _07560_);
  and (_11369_, _11052_, _07601_);
  or (_11370_, _11369_, _11368_);
  or (_11371_, _11370_, _11124_);
  or (_11372_, _11371_, _11366_);
  not (_11373_, _08862_);
  or (_11374_, _11129_, _11373_);
  and (_11375_, _07721_, _07564_);
  or (_11376_, _11375_, _11082_);
  or (_11377_, _11376_, _11175_);
  or (_11378_, _11377_, _11374_);
  and (_11379_, _07602_, _07654_);
  and (_11380_, _11160_, _07560_);
  and (_11381_, _07602_, _07666_);
  or (_11382_, _11381_, _11380_);
  or (_11383_, _11382_, _11379_);
  or (_11384_, _11161_, _11061_);
  or (_11385_, _11384_, _11313_);
  and (_11386_, _07654_, _07643_);
  or (_11387_, _11386_, _11267_);
  or (_11388_, _11387_, _07693_);
  or (_11389_, _11388_, _11385_);
  or (_11390_, _11389_, _11383_);
  or (_11391_, _11390_, _11378_);
  or (_11392_, _11391_, _11372_);
  and (_11393_, _11392_, _10941_);
  or (_12687_[0], _11393_, _11364_);
  or (_11394_, _11328_, _11142_);
  or (_11395_, _11064_, _07674_);
  or (_11396_, _11395_, _11394_);
  or (_11397_, _11396_, _11147_);
  or (_11398_, _11397_, _11315_);
  or (_11399_, _11379_, _11375_);
  or (_11400_, _11368_, _11256_);
  or (_11401_, _11400_, _11399_);
  or (_11402_, _11060_, _07597_);
  or (_11403_, _07606_, _07603_);
  or (_11404_, _11403_, _11402_);
  not (_11405_, _07685_);
  or (_11406_, _11405_, _07582_);
  or (_11407_, _11406_, _11404_);
  or (_11408_, _11407_, _11401_);
  or (_11409_, _11408_, _11398_);
  and (_11410_, _11409_, _10941_);
  and (_11411_, _07308_, _12493_);
  and (_11412_, _11411_, _07723_);
  and (_11413_, _11043_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_11414_, _11413_, _11412_);
  or (_12688_[0], _11414_, _11410_);
  and (_11415_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11416_, _07723_, _05610_);
  or (_11417_, _11416_, _11415_);
  and (_11418_, _11417_, _12493_);
  or (_11419_, _11089_, _07675_);
  or (_11420_, _11419_, _11168_);
  or (_11421_, _11420_, _11323_);
  or (_11422_, _11261_, _11255_);
  and (_11423_, _07666_, _07440_);
  or (_11424_, _11423_, _11245_);
  or (_11425_, _11424_, _11422_);
  or (_11426_, _11425_, _11421_);
  not (_11427_, _07683_);
  nor (_11428_, _11263_, _07684_);
  and (_11429_, _11428_, _11427_);
  or (_11430_, _11064_, _07587_);
  and (_11431_, _07602_, _07522_);
  or (_11432_, _11431_, _11384_);
  nor (_11433_, _11432_, _11430_);
  nand (_11434_, _11433_, _11429_);
  or (_11435_, _11434_, _11426_);
  or (_11436_, _11088_, _11083_);
  or (_11437_, _11436_, _11435_);
  and (_11438_, _11437_, _10941_);
  or (_12688_[1], _11438_, _11418_);
  not (_11439_, _11428_);
  or (_11440_, _11439_, _11422_);
  or (_11441_, _11440_, _11424_);
  or (_11442_, _07583_, _07573_);
  nor (_11443_, _11442_, _11367_);
  nand (_11444_, _11443_, _08861_);
  or (_11445_, _11376_, _11130_);
  or (_11446_, _11445_, _11444_);
  or (_11447_, _11087_, _11081_);
  or (_11448_, _11447_, _11446_);
  or (_11449_, _11448_, _11441_);
  and (_11450_, _11449_, _07312_);
  and (_11451_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11452_, _07722_, _05610_);
  or (_11453_, _11452_, _11451_);
  or (_11454_, _11453_, _11450_);
  and (_12688_[2], _11454_, _12493_);
  and (_11455_, _11043_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_11456_, _11053_, _07691_);
  nand (_11457_, _11456_, _08862_);
  not (_11458_, _07413_);
  or (_11459_, _07602_, _11458_);
  and (_11460_, _11459_, _07666_);
  or (_11461_, _11460_, _11399_);
  or (_11462_, _11461_, _11457_);
  or (_11463_, _11370_, _11167_);
  or (_11464_, _11463_, _11366_);
  or (_11465_, _11464_, _11462_);
  and (_11466_, _11465_, _10941_);
  or (_12689_[0], _11466_, _11455_);
  nor (_12675_[7], _07462_, rst);
  nor (_12676_[7], _09086_, rst);
  and (_11467_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_11468_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_11469_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_11470_, _07329_, _09077_);
  nor (_11471_, _11470_, _11469_);
  and (_11472_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_11473_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_11474_, _11473_, _11472_);
  and (_11475_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  not (_11476_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_11477_, _07324_, _11476_);
  nor (_11478_, _11477_, _11475_);
  and (_11479_, _11478_, _11474_);
  and (_11480_, _11479_, _11471_);
  nor (_11481_, _11480_, _07318_);
  nor (_11482_, _11481_, _11468_);
  nor (_11483_, _11482_, _08951_);
  nor (_11484_, _11483_, _11467_);
  nor (_12677_[7], _11484_, rst);
  nor (_12675_[0], _07355_, rst);
  and (_12675_[1], _07433_, _12493_);
  nor (_12675_[2], _07381_, rst);
  nor (_12675_[3], _07407_, rst);
  and (_12675_[4], _07546_, _12493_);
  nor (_12675_[5], _07515_, rst);
  nor (_12675_[6], _07488_, rst);
  nor (_12676_[0], _09140_, rst);
  nor (_12676_[1], _09294_, rst);
  nor (_12676_[2], _08968_, rst);
  nor (_12676_[3], _09189_, rst);
  nor (_12676_[4], _09343_, rst);
  nor (_12676_[5], _09014_, rst);
  nor (_12676_[6], _09244_, rst);
  and (_11485_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_11486_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_11487_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_11488_, _07329_, _09130_);
  nor (_11489_, _11488_, _11487_);
  and (_11490_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_11491_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_11492_, _11491_, _11490_);
  and (_11493_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not (_11494_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_11495_, _07324_, _11494_);
  nor (_11496_, _11495_, _11493_);
  and (_11497_, _11496_, _11492_);
  and (_11498_, _11497_, _11489_);
  nor (_11499_, _11498_, _07318_);
  nor (_11500_, _11499_, _11486_);
  nor (_11501_, _11500_, _08951_);
  nor (_11502_, _11501_, _11485_);
  nor (_12677_[0], _11502_, rst);
  and (_11503_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_11504_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_11505_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_11506_, _07420_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_11507_, _11506_, _11505_);
  and (_11508_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_11509_, _07417_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_11510_, _11509_, _11508_);
  and (_11511_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_11512_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_11513_, _11512_, _11511_);
  and (_11514_, _11513_, _11510_);
  and (_11515_, _11514_, _11507_);
  nor (_11516_, _11515_, _07318_);
  nor (_11517_, _11516_, _11504_);
  nor (_11518_, _11517_, _08951_);
  nor (_11519_, _11518_, _11503_);
  nor (_12677_[1], _11519_, rst);
  and (_11520_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_11521_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_11522_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor (_11523_, _07329_, _08959_);
  nor (_11524_, _11523_, _11522_);
  and (_11525_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_11526_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11527_, _11526_, _11525_);
  and (_11528_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not (_11529_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_11530_, _07324_, _11529_);
  nor (_11531_, _11530_, _11528_);
  and (_11532_, _11531_, _11527_);
  and (_11533_, _11532_, _11524_);
  nor (_11534_, _11533_, _07318_);
  nor (_11535_, _11534_, _11521_);
  nor (_11536_, _11535_, _08951_);
  nor (_11537_, _11536_, _11520_);
  nor (_12677_[2], _11537_, rst);
  and (_11538_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_11539_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_11540_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_11541_, _07329_, _09177_);
  nor (_11542_, _11541_, _11540_);
  and (_11543_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_11544_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_11545_, _11544_, _11543_);
  and (_11546_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not (_11547_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_11548_, _07324_, _11547_);
  nor (_11549_, _11548_, _11546_);
  and (_11550_, _11549_, _11545_);
  and (_11551_, _11550_, _11542_);
  nor (_11552_, _11551_, _07318_);
  nor (_11553_, _11552_, _11539_);
  nor (_11554_, _11553_, _08951_);
  nor (_11555_, _11554_, _11538_);
  nor (_12677_[3], _11555_, rst);
  and (_11556_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_11557_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_11558_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_11559_, _07420_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_11560_, _11559_, _11558_);
  and (_11561_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_11562_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_11563_, _11562_, _11561_);
  and (_11564_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_11565_, _07417_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_11566_, _11565_, _11564_);
  and (_11567_, _11566_, _11563_);
  and (_11568_, _11567_, _11560_);
  nor (_11569_, _11568_, _07318_);
  nor (_11570_, _11569_, _11557_);
  nor (_11571_, _11570_, _08951_);
  nor (_11572_, _11571_, _11556_);
  nor (_12677_[4], _11572_, rst);
  and (_11573_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_11574_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_11575_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_11576_, _07329_, _09008_);
  nor (_11577_, _11576_, _11575_);
  and (_11578_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_11579_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_11580_, _11579_, _11578_);
  and (_11581_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  not (_11582_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_11583_, _07324_, _11582_);
  nor (_11584_, _11583_, _11581_);
  and (_11585_, _11584_, _11580_);
  and (_11586_, _11585_, _11577_);
  nor (_11587_, _11586_, _07318_);
  nor (_11588_, _11587_, _11574_);
  nor (_11589_, _11588_, _08951_);
  nor (_11590_, _11589_, _11573_);
  nor (_12677_[5], _11590_, rst);
  and (_11591_, _08951_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_11592_, _07318_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_11593_, _07345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_11594_, _07329_, _09238_);
  nor (_11595_, _11594_, _11593_);
  and (_11596_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not (_11597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_11598_, _07324_, _11597_);
  nor (_11599_, _11598_, _11596_);
  and (_11600_, _11599_, _11595_);
  and (_11601_, _07335_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_11602_, _07342_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_11603_, _11602_, _11601_);
  and (_11604_, _11603_, _11600_);
  nor (_11605_, _11604_, _07318_);
  nor (_11606_, _11605_, _11592_);
  nor (_11607_, _11606_, _08951_);
  nor (_11608_, _11607_, _11591_);
  nor (_12677_[6], _11608_, rst);
  and (_11609_, _07313_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_11610_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_11611_, _11609_, _07947_);
  and (_11612_, _11611_, _12493_);
  and (_12692_[15], _11612_, _11610_);
  not (_11613_, _11609_);
  or (_11614_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00002_, _11609_, _12493_);
  and (_11615_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _12493_);
  or (_11616_, _11615_, _00002_);
  and (_12693_[15], _11616_, _11614_);
  nor (_12694_, _09092_, rst);
  and (_12695_, \oc8051_top_1.oc8051_memory_interface1.dstb_o , _12493_);
  nor (_12696_[4], _09348_, rst);
  and (_12697_[7], _09069_, _12493_);
  not (_11617_, _07620_);
  not (_11618_, _06423_);
  nor (_11619_, _09250_, _11618_);
  and (_11620_, _09250_, _11618_);
  nor (_11621_, _11620_, _11619_);
  or (_11622_, _09092_, _06452_);
  nand (_11623_, _09092_, _06452_);
  and (_11624_, _11623_, _11622_);
  and (_11625_, _11624_, _11621_);
  or (_11626_, _09023_, _08316_);
  nand (_11627_, _09023_, _08316_);
  and (_11628_, _11627_, _11626_);
  or (_11629_, _09354_, _07736_);
  nand (_11630_, _09354_, _07736_);
  and (_11631_, _11630_, _11629_);
  and (_11632_, _11631_, _11628_);
  and (_11633_, _11632_, _11625_);
  nor (_11634_, _09145_, _06498_);
  and (_11635_, _09145_, _06498_);
  nor (_11636_, _11635_, _11634_);
  and (_11637_, _09304_, _07012_);
  nor (_11638_, _09304_, _07012_);
  or (_11639_, _11638_, _11637_);
  nor (_11640_, _11639_, _11636_);
  nor (_11641_, _09194_, _06469_);
  and (_11642_, _09194_, _06469_);
  nor (_11643_, _11642_, _11641_);
  nor (_11644_, _08973_, _06520_);
  and (_11645_, _08973_, _06520_);
  nor (_11646_, _11645_, _11644_);
  not (_11647_, _11646_);
  and (_11648_, _11647_, _11643_);
  and (_11649_, _11648_, _11640_);
  and (_11650_, _11649_, _11633_);
  and (_11651_, _11650_, _06776_);
  nor (_11652_, _06451_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_11653_, _11652_, _11651_);
  not (_11654_, _11653_);
  and (_11655_, _11633_, _11643_);
  nor (_11656_, _07658_, _11071_);
  and (_11657_, _07293_, _06777_);
  and (_11658_, _11657_, _11656_);
  and (_11659_, _11658_, _11655_);
  and (_11660_, _06969_, _06586_);
  nand (_11661_, _11660_, _07030_);
  nor (_11662_, _11661_, _07089_);
  and (_11663_, _11662_, _07161_);
  and (_11664_, _11663_, _07239_);
  and (_11665_, _09026_, _07709_);
  nor (_11666_, _11665_, _11071_);
  nor (_11667_, _11666_, _07705_);
  and (_11668_, _11667_, _06845_);
  and (_11669_, _11668_, _11664_);
  and (_11670_, _11669_, _06642_);
  and (_11671_, _11656_, _06619_);
  nor (_11672_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_11673_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_11674_, _11673_, _11672_);
  nor (_11675_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_11676_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_11677_, _11676_, _11675_);
  and (_11678_, _11677_, _11674_);
  and (_11679_, _11678_, _07618_);
  not (_11680_, _07705_);
  nor (_11681_, _11656_, _07520_);
  nor (_11682_, _11681_, _11680_);
  and (_11683_, _11682_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_11684_, _11683_, _11679_);
  or (_11685_, _11684_, _11671_);
  nor (_11686_, _11685_, _11670_);
  or (_11687_, _11322_, _07671_);
  nor (_11688_, _11687_, _11117_);
  or (_11689_, _07605_, _07654_);
  nor (_11690_, _11689_, _07580_);
  nor (_11691_, _11690_, _07653_);
  nor (_11692_, _11691_, _11283_);
  and (_11693_, _11692_, _11688_);
  not (_11694_, _11693_);
  and (_11695_, _11694_, _11686_);
  not (_11696_, _11695_);
  and (_11697_, _07704_, _07551_);
  not (_11698_, _11697_);
  and (_11699_, _11698_, _07711_);
  nor (_11700_, _11699_, _11686_);
  and (_11701_, _11121_, _07605_);
  nor (_11702_, _11701_, _11049_);
  not (_11703_, _11702_);
  nor (_11704_, _11703_, _11700_);
  and (_11705_, _11704_, _11696_);
  nor (_11706_, _11705_, _07706_);
  not (_11707_, _11706_);
  nor (_11708_, _11108_, _07308_);
  nor (_11709_, _11708_, _07619_);
  and (_11710_, _11709_, _11707_);
  nor (_11711_, _08335_, _08329_);
  not (_11712_, _11711_);
  and (_11713_, _11712_, _07618_);
  not (_11714_, _08205_);
  nor (_11715_, _08215_, _11714_);
  and (_11716_, _11715_, _08281_);
  not (_11717_, _11716_);
  and (_11718_, _11717_, _11682_);
  nor (_11719_, _11718_, _11713_);
  not (_11720_, _11719_);
  nor (_11721_, _11720_, _11710_);
  not (_11722_, _11721_);
  nor (_11723_, _11722_, _11659_);
  and (_11724_, _11723_, _11654_);
  and (_11725_, _11724_, _11617_);
  and (_12700_, _11725_, _12493_);
  and (_12701_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _12493_);
  nor (_11726_, \oc8051_top_1.oc8051_memory_interface1.dstb_o , rst);
  and (_11727_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_11728_, _12695_, xram_data_in_reg[7]);
  or (_12702_[7], _11728_, _11727_);
  nor (_11729_, _07344_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_11730_, _11729_, _08951_);
  nor (_11731_, _11730_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_11732_, _11731_);
  and (_11733_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_11734_, _11733_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_11735_, _11734_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_11736_, _11735_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_11737_, _11736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_11738_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_11739_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_11740_, _11739_, _11738_);
  and (_11741_, _11740_, _11737_);
  and (_11742_, _11741_, _11732_);
  and (_11743_, _11742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_11744_, _11743_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_11745_, _11744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_11746_, _11745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_11747_, _11745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_11748_, _11747_, _11746_);
  or (_11749_, _11748_, _11724_);
  and (_11750_, _11749_, _12493_);
  nor (_11751_, _11687_, _11283_);
  nand (_11752_, _11751_, _11665_);
  nand (_11753_, _11752_, _07616_);
  and (_11754_, _11107_, _07727_);
  and (_11755_, _07651_, _07727_);
  or (_11756_, _11755_, _11754_);
  nor (_11757_, _11756_, _07620_);
  and (_11758_, _11757_, _11753_);
  and (_11759_, _11758_, _09086_);
  nand (_11760_, _11757_, _11753_);
  and (_11761_, _11760_, _11484_);
  nor (_11762_, _11761_, _11759_);
  and (_11763_, _11762_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_11764_, _11762_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_11765_, _11764_);
  and (_11766_, _11758_, _09244_);
  and (_11767_, _11760_, _11608_);
  nor (_11768_, _11767_, _11766_);
  and (_11769_, _11768_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_11770_, _11769_);
  nor (_11771_, _11768_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_11772_, _11771_, _11769_);
  and (_11773_, _11758_, _09014_);
  and (_11774_, _11760_, _11590_);
  nor (_11775_, _11774_, _11773_);
  nor (_11776_, _11775_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_11777_, _11775_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_11778_, _11758_, _09343_);
  and (_11779_, _11760_, _11572_);
  nor (_11780_, _11779_, _11778_);
  nand (_11781_, _11780_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_11782_, _11758_, _09189_);
  and (_11783_, _11760_, _11555_);
  nor (_11784_, _11783_, _11782_);
  nor (_11785_, _11784_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_11786_, _11784_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_11787_, _11760_, _08969_);
  not (_11788_, _11537_);
  or (_11789_, _11758_, _11788_);
  nand (_11790_, _11789_, _11787_);
  or (_11791_, _11790_, _05897_);
  or (_11792_, _11760_, _09295_);
  not (_11793_, _11519_);
  or (_11794_, _11758_, _11793_);
  and (_11795_, _11794_, _11792_);
  nand (_11796_, _11795_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_11797_, _11760_, _09141_);
  not (_11798_, _11502_);
  or (_11799_, _11758_, _11798_);
  and (_11800_, _11799_, _11797_);
  and (_11801_, _11800_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_11802_, _11795_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_11803_, _11802_, _11796_);
  and (_11804_, _11803_, _11801_);
  not (_11805_, _11804_);
  nand (_11806_, _11805_, _11796_);
  nand (_11807_, _11790_, _05897_);
  and (_11808_, _11807_, _11791_);
  and (_11809_, _11808_, _11806_);
  not (_11810_, _11809_);
  nand (_11811_, _11810_, _11791_);
  nor (_11812_, _11811_, _11786_);
  nor (_11813_, _11812_, _11785_);
  or (_11814_, _11780_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_11815_, _11814_, _11781_);
  nand (_11816_, _11815_, _11813_);
  nand (_11817_, _11816_, _11781_);
  nor (_11818_, _11817_, _11777_);
  nor (_11819_, _11818_, _11776_);
  nand (_11820_, _11819_, _11772_);
  nand (_11821_, _11820_, _11770_);
  and (_11822_, _11821_, _11765_);
  nor (_11823_, _11822_, _11763_);
  and (_11824_, _11823_, _07919_);
  nand (_11825_, _11824_, _07925_);
  or (_11826_, _11825_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_11827_, _11826_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_11828_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_11829_, _11828_, _11827_);
  nand (_11830_, _11829_, _07942_);
  and (_11831_, _11830_, _11762_);
  or (_11832_, _11822_, _11763_);
  and (_11833_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_11834_, _11833_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_11835_, _11834_, _11832_);
  and (_11836_, _11835_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_11837_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_11838_, _11837_, _11836_);
  and (_11839_, _11838_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_11840_, _11839_, _11762_);
  or (_11841_, _11840_, _11831_);
  nand (_11842_, _11841_, _07947_);
  or (_11843_, _11841_, _07947_);
  and (_11844_, _11843_, _11842_);
  and (_11845_, _07559_, _07727_);
  and (_11846_, _11845_, _07522_);
  nor (_11847_, _11283_, _07704_);
  and (_11848_, _11847_, _11702_);
  and (_11849_, _11688_, _11665_);
  and (_11850_, _11849_, _11848_);
  nor (_11851_, _11850_, _07706_);
  nor (_11852_, _11851_, _11846_);
  not (_11853_, _11846_);
  nor (_11854_, _11754_, _07702_);
  and (_11855_, _11854_, _11753_);
  and (_11856_, _11855_, _11853_);
  and (_11857_, _11701_, _07616_);
  nor (_11858_, _11857_, _11708_);
  not (_11859_, _11858_);
  and (_11860_, _11859_, _11856_);
  nor (_11861_, _11860_, _11852_);
  and (_11862_, _11861_, _11844_);
  nand (_11863_, _11651_, _06452_);
  or (_11864_, _11863_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_11865_, _07559_, _07526_);
  and (_11866_, _11865_, _07616_);
  and (_11867_, _11712_, _11866_);
  nor (_11868_, _11867_, _11710_);
  and (_11869_, _07705_, _07520_);
  and (_11870_, _11717_, _11869_);
  and (_11871_, _11666_, _07293_);
  and (_11872_, _11871_, _06777_);
  and (_11873_, _11872_, _11655_);
  nor (_11874_, _11873_, _11870_);
  and (_11875_, _11874_, _11868_);
  and (_11876_, _11875_, _11864_);
  and (_11877_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_11878_, _11877_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_11879_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_11880_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_11881_, _11880_, _11879_);
  and (_11882_, _11881_, _11878_);
  and (_11883_, _11882_, _11834_);
  and (_11884_, _11883_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_11885_, _11884_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_11886_, _11885_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_11887_, _11886_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_11888_, _11887_, _07947_);
  or (_11889_, _11887_, _07947_);
  and (_11890_, _11889_, _11888_);
  not (_11891_, _11851_);
  and (_11892_, _11860_, _11891_);
  and (_11893_, _11892_, _11890_);
  nor (_11894_, _07703_, _06770_);
  and (_11895_, _11857_, _07958_);
  and (_11896_, _11754_, _09087_);
  and (_11897_, _07616_, _07606_);
  nor (_11898_, _11897_, _11708_);
  and (_11899_, _11898_, _11758_);
  and (_11900_, _11899_, _11891_);
  and (_11901_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_11902_, _11901_, _11896_);
  or (_11903_, _11902_, _11895_);
  or (_11904_, _11903_, _11894_);
  nor (_11905_, _11904_, _11893_);
  nand (_11906_, _11905_, _11876_);
  or (_11907_, _11906_, _11862_);
  and (_12703_[15], _11907_, _11750_);
  and (_11908_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12493_);
  and (_11909_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_11910_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11911_, _07312_, _11910_);
  not (_11912_, _11911_);
  not (_11913_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_11914_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_11915_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_11916_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_11917_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_11918_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_11919_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_11920_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_11921_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_11922_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_11923_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_11924_, _11923_, _11922_);
  and (_11925_, _11924_, _11921_);
  and (_11926_, _11925_, _11920_);
  and (_11927_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_11928_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_11929_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_11930_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_11931_, _11930_, _11928_);
  and (_11932_, _11931_, _11929_);
  nor (_11933_, _11932_, _11928_);
  nor (_11934_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_11935_, _11934_, _11927_);
  not (_11936_, _11935_);
  nor (_11937_, _11936_, _11933_);
  nor (_11938_, _11937_, _11927_);
  and (_11939_, _11938_, _11926_);
  and (_11940_, _11939_, _11919_);
  and (_11941_, _11940_, _11918_);
  and (_11942_, _11941_, _11917_);
  and (_11943_, _11942_, _11916_);
  and (_11944_, _11943_, _11915_);
  and (_11945_, _11944_, _11914_);
  and (_11946_, _11945_, _11913_);
  nor (_11947_, _11946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_11948_, _11946_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_11949_, _11948_, _11947_);
  nor (_11950_, _11945_, _11913_);
  nor (_11951_, _11950_, _11946_);
  not (_11952_, _11951_);
  nor (_11953_, _11944_, _11914_);
  or (_11954_, _11953_, _11945_);
  nor (_11955_, _11943_, _11915_);
  nor (_11956_, _11955_, _11944_);
  not (_11957_, _11956_);
  nor (_11958_, _11942_, _11916_);
  nor (_11959_, _11958_, _11943_);
  not (_11960_, _11959_);
  nor (_11961_, _11941_, _11917_);
  nor (_11962_, _11961_, _11942_);
  not (_11963_, _11962_);
  nor (_11964_, _11940_, _11918_);
  or (_11965_, _11964_, _11941_);
  and (_11966_, _11938_, _11925_);
  nor (_11967_, _11966_, _11920_);
  or (_11968_, _11967_, _11939_);
  and (_11969_, _11938_, _11924_);
  nor (_11970_, _11969_, _11921_);
  nor (_11971_, _11970_, _11966_);
  not (_11972_, _11971_);
  and (_11973_, _11938_, _11923_);
  nor (_11974_, _11973_, _11922_);
  nor (_11975_, _11974_, _11969_);
  not (_11976_, _11975_);
  not (_11977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_11978_, _11938_, _11977_);
  nor (_11979_, _11938_, _11977_);
  nor (_11980_, _11979_, _11978_);
  not (_11981_, _11980_);
  and (_11982_, _11019_, _10993_);
  not (_11983_, _11982_);
  and (_11984_, _10996_, _10966_);
  and (_11985_, _11017_, _10958_);
  nor (_11986_, _11985_, _11984_);
  and (_11987_, _11986_, _11983_);
  not (_11988_, _10946_);
  nor (_11989_, _11025_, _10983_);
  nor (_11990_, _11989_, _11988_);
  not (_11991_, _10966_);
  and (_11992_, _10998_, _10952_);
  not (_11993_, _11992_);
  and (_11994_, _10982_, _07515_);
  nor (_11995_, _11027_, _11994_);
  and (_11996_, _11995_, _11993_);
  nor (_11997_, _11996_, _11991_);
  nor (_11998_, _11997_, _11990_);
  and (_11999_, _10952_, _10981_);
  and (_12000_, _11999_, _10958_);
  and (_12001_, _10982_, _10964_);
  nor (_12002_, _12001_, _10996_);
  nor (_12003_, _12002_, _11988_);
  nor (_12004_, _12003_, _12000_);
  and (_12005_, _12004_, _11998_);
  and (_12006_, _12005_, _11987_);
  and (_12007_, _12006_, _11022_);
  and (_12008_, _10990_, _10959_);
  not (_12009_, _12008_);
  and (_12010_, _10952_, _10953_);
  and (_12011_, _10955_, _07433_);
  and (_12012_, _12011_, _12010_);
  not (_12013_, _12012_);
  and (_12014_, _11012_, _10968_);
  and (_12015_, _12014_, _10971_);
  nor (_12016_, _12015_, _11004_);
  and (_12017_, _12016_, _12013_);
  and (_12018_, _12017_, _12009_);
  and (_12019_, _11012_, _10981_);
  nor (_12020_, _10985_, _10946_);
  not (_12021_, _12020_);
  and (_12022_, _12021_, _12019_);
  not (_12023_, _10986_);
  nor (_12024_, _11025_, _10965_);
  nor (_12025_, _11019_, _11002_);
  and (_12026_, _12025_, _12024_);
  nor (_12027_, _12026_, _12023_);
  nor (_12028_, _12027_, _12022_);
  and (_12029_, _12028_, _12018_);
  and (_12030_, _11999_, _10966_);
  nor (_12031_, _12001_, _11999_);
  nor (_12032_, _12031_, _12023_);
  nor (_12033_, _12032_, _12030_);
  nor (_12034_, _12010_, _11025_);
  nor (_12035_, _12034_, _07407_);
  nor (_12036_, _10999_, _10947_);
  nor (_12037_, _12036_, _12023_);
  nor (_12038_, _12037_, _12035_);
  and (_12039_, _12038_, _12033_);
  and (_12040_, _11025_, _10958_);
  nor (_12041_, _12040_, _10949_);
  and (_12042_, _12041_, _10976_);
  and (_12043_, _12042_, _12039_);
  and (_12044_, _12043_, _12029_);
  nand (_12045_, _10997_, _10956_);
  and (_12046_, _10996_, _10958_);
  and (_12047_, _12019_, _10993_);
  nor (_12048_, _12047_, _12046_);
  and (_12049_, _12048_, _12045_);
  and (_12050_, _12049_, _10988_);
  nor (_12051_, _10985_, _10945_);
  and (_12052_, _11019_, _07355_);
  nor (_12053_, _12052_, _11013_);
  nor (_12054_, _12053_, _12051_);
  and (_12055_, _10952_, _10946_);
  and (_12056_, _12055_, _10978_);
  and (_12057_, _10965_, _10946_);
  nor (_12058_, _12057_, _12056_);
  not (_12059_, _12058_);
  nor (_12060_, _12059_, _12054_);
  and (_12061_, _12060_, _12050_);
  and (_12062_, _12061_, _12044_);
  and (_12063_, _12062_, _12007_);
  not (_12064_, _12063_);
  nor (_12065_, _11931_, _11929_);
  nor (_12066_, _12065_, _11932_);
  nand (_12067_, _12066_, _12064_);
  or (_12068_, _11018_, _10975_);
  or (_12069_, _12030_, _10949_);
  nor (_12070_, _12024_, _12023_);
  and (_12071_, _11012_, _10953_);
  and (_12072_, _12071_, _10993_);
  or (_12073_, _12072_, _12070_);
  or (_12074_, _12073_, _12069_);
  nor (_12075_, _12074_, _12068_);
  nand (_12076_, _12075_, _12050_);
  nor (_12077_, _12076_, _12063_);
  not (_12078_, _12077_);
  nor (_12079_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_12080_, _12079_, _11929_);
  and (_12081_, _12080_, _12078_);
  or (_12082_, _12066_, _12064_);
  and (_12083_, _12082_, _12067_);
  nand (_12084_, _12083_, _12081_);
  and (_12085_, _12084_, _12067_);
  not (_12086_, _12085_);
  and (_12087_, _11936_, _11933_);
  nor (_12088_, _12087_, _11937_);
  and (_12089_, _12088_, _12086_);
  and (_12090_, _12089_, _11981_);
  not (_12091_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_12092_, _11978_, _12091_);
  or (_12093_, _12092_, _11973_);
  and (_12094_, _12093_, _12090_);
  and (_12095_, _12094_, _11976_);
  and (_12096_, _12095_, _11972_);
  and (_12097_, _12096_, _11968_);
  nor (_12098_, _11939_, _11919_);
  or (_12099_, _12098_, _11940_);
  and (_12100_, _12099_, _12097_);
  and (_12101_, _12100_, _11965_);
  and (_12102_, _12101_, _11963_);
  and (_12103_, _12102_, _11960_);
  and (_12104_, _12103_, _11957_);
  and (_12105_, _12104_, _11954_);
  and (_12106_, _12105_, _11952_);
  or (_12107_, _12106_, _11949_);
  nand (_12108_, _12106_, _11949_);
  and (_12109_, _12108_, _12107_);
  or (_12110_, _12109_, _11912_);
  or (_12111_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_12112_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_12113_, _12112_, _12111_);
  and (_12114_, _12113_, _12110_);
  or (_12704_[15], _12114_, _11909_);
  nor (_12115_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_12705_, _12115_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_12706_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _12493_);
  and (_12116_, \oc8051_top_1.oc8051_rom1.ea_int , _07309_);
  nand (_12117_, _12116_, _07312_);
  and (_12707_, _12117_, _12706_);
  and (_12708_[7], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _12493_);
  nor (_12118_, _11731_, _08951_);
  or (_12119_, _12063_, _07327_);
  nor (_12120_, _12077_, _07322_);
  nand (_12121_, _12063_, _07327_);
  and (_12122_, _12121_, _12119_);
  nand (_12123_, _12122_, _12120_);
  and (_12124_, _12123_, _12119_);
  nor (_12125_, _12124_, _08951_);
  and (_12126_, _12125_, _07321_);
  nor (_12127_, _12125_, _07321_);
  nor (_12128_, _12127_, _12126_);
  nor (_12129_, _12128_, _12118_);
  and (_12130_, _07328_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_12131_, _12130_, _12118_);
  and (_12132_, _12131_, _12076_);
  or (_12133_, _12132_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_12134_, _12133_, _12129_);
  and (_12709_[2], _12134_, _12493_);
  and (_12135_, _07427_, _07375_);
  and (_12136_, _07540_, _07456_);
  and (_12137_, _12136_, _12135_);
  and (_12138_, _07313_, _12493_);
  and (_12139_, _12138_, _07482_);
  and (_12140_, _12139_, _07510_);
  and (_12141_, _07402_, _07350_);
  and (_12142_, _12141_, _12140_);
  and (_12712_, _12142_, _12137_);
  not (_12143_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_12144_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_12145_, _12144_, _12143_);
  or (_12146_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_12147_, _12146_, _12493_);
  and (_12713_[7], _12147_, _12145_);
  and (_12714_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _12493_);
  not (_12148_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_12149_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_12150_, _12149_, _12148_);
  and (_12151_, _12149_, _12148_);
  nor (_12152_, _12151_, _12150_);
  not (_12153_, _12152_);
  and (_12154_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_12155_, _12154_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_12156_, _12154_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_12157_, _12156_, _12155_);
  or (_12158_, _12157_, _12149_);
  and (_12159_, _12158_, _12153_);
  nor (_12160_, _12150_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_12161_, _12150_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_12162_, _12161_, _12160_);
  or (_12163_, _12155_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_12716_[3], _12163_, _12493_);
  and (_12164_, _12716_[3], _12162_);
  and (_12715_, _12164_, _12159_);
  not (_12165_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_12166_, _11731_, _12165_);
  and (_12167_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_12168_, _12166_);
  and (_12169_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_12170_, _12169_, _12167_);
  and (_12717_[31], _12170_, _12493_);
  and (_12171_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_12172_, _12166_, _09077_);
  or (_12173_, _12172_, _12171_);
  and (_12718_[31], _12173_, _12493_);
  not (_12174_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  nor (_12175_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  nor (_12176_, _12175_, _12174_);
  and (_12177_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_12178_, _12177_, _12175_);
  or (_12179_, _12178_, _12176_);
  and (_12719_[7], _12179_, _12493_);
  and (_12180_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  not (_12181_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_12182_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _12181_);
  or (_12183_, _12182_, _12180_);
  and (_12720_, _12183_, _11726_);
  and (_12721_, _12175_, _12493_);
  not (_12184_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  nor (_12185_, _12175_, _12184_);
  not (_12186_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_12187_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_12188_, _12187_, _12175_);
  or (_12189_, _12188_, _12185_);
  and (_12722_[15], _12189_, _12493_);
  or (_12190_, _12181_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_12723_, _12190_, _11726_);
  nor (_12191_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_12192_, _12191_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_12193_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_12194_, _12193_, _12192_);
  and (_12724_, _12194_, _12493_);
  and (_12195_, _12165_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_12196_, _12195_, _12192_);
  and (_12725_, _12196_, _12493_);
  not (_12197_, _12192_);
  or (_12198_, _12197_, _07958_);
  or (_12199_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_12200_, _12199_, _12493_);
  and (_12726_[15], _12200_, _12198_);
  and (_12727_, _07734_, _08870_);
  or (_12201_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_12202_, _11609_, _05929_);
  and (_12203_, _12202_, _12493_);
  and (_12692_[0], _12203_, _12201_);
  or (_12204_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_12205_, _11609_, _05879_);
  and (_12206_, _12205_, _12493_);
  and (_12692_[1], _12206_, _12204_);
  or (_12207_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_12208_, _11609_, _05897_);
  and (_12209_, _12208_, _12493_);
  and (_12692_[2], _12209_, _12207_);
  or (_12210_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_12211_, _11609_, _05782_);
  and (_12212_, _12211_, _12493_);
  and (_12692_[3], _12212_, _12210_);
  or (_12213_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_12214_, _11609_, _05633_);
  and (_12215_, _12214_, _12493_);
  and (_12692_[4], _12215_, _12213_);
  or (_12216_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_12217_, _11609_, _05800_);
  and (_12218_, _12217_, _12493_);
  and (_12692_[5], _12218_, _12216_);
  or (_12219_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_12220_, _11609_, _05821_);
  and (_12221_, _12220_, _12493_);
  and (_12692_[6], _12221_, _12219_);
  or (_12222_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_12223_, _11609_, _05852_);
  and (_12224_, _12223_, _12493_);
  and (_12692_[7], _12224_, _12222_);
  or (_12225_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_12226_, _11609_, _07919_);
  and (_12227_, _12226_, _12493_);
  and (_12692_[8], _12227_, _12225_);
  or (_12228_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_12229_, _11609_, _07925_);
  and (_12230_, _12229_, _12493_);
  and (_12692_[9], _12230_, _12228_);
  or (_12231_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_12232_, _11609_, _07930_);
  and (_12233_, _12232_, _12493_);
  and (_12692_[10], _12233_, _12231_);
  or (_12234_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_12235_, _11609_, _07915_);
  and (_12236_, _12235_, _12493_);
  and (_12692_[11], _12236_, _12234_);
  or (_12237_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_12238_, _11609_, _07936_);
  and (_12239_, _12238_, _12493_);
  and (_12692_[12], _12239_, _12237_);
  or (_12240_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_12241_, _11609_, _07911_);
  and (_12242_, _12241_, _12493_);
  and (_12692_[13], _12242_, _12240_);
  or (_12243_, _11609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_12244_, _11609_, _07942_);
  and (_12245_, _12244_, _12493_);
  and (_12692_[14], _12245_, _12243_);
  or (_12246_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_12247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _12493_);
  or (_12248_, _12247_, _00002_);
  and (_12693_[0], _12248_, _12246_);
  or (_12249_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_12250_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _12493_);
  or (_12251_, _12250_, _00002_);
  and (_12693_[1], _12251_, _12249_);
  or (_12252_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_12253_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _12493_);
  or (_12254_, _12253_, _00002_);
  and (_12693_[2], _12254_, _12252_);
  or (_12255_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_12256_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _12493_);
  or (_12257_, _12256_, _00002_);
  and (_12693_[3], _12257_, _12255_);
  or (_12258_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_12259_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _12493_);
  or (_12260_, _12259_, _00002_);
  and (_12693_[4], _12260_, _12258_);
  or (_12261_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_12262_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _12493_);
  or (_12263_, _12262_, _00002_);
  and (_12693_[5], _12263_, _12261_);
  or (_12264_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_12265_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _12493_);
  or (_12266_, _12265_, _00002_);
  and (_12693_[6], _12266_, _12264_);
  or (_12267_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_12268_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _12493_);
  or (_12269_, _12268_, _00002_);
  and (_12693_[7], _12269_, _12267_);
  or (_12270_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_12271_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _12493_);
  or (_12272_, _12271_, _00002_);
  and (_12693_[8], _12272_, _12270_);
  or (_12273_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_12274_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _12493_);
  or (_12275_, _12274_, _00002_);
  and (_12693_[9], _12275_, _12273_);
  or (_12276_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_12277_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _12493_);
  or (_12278_, _12277_, _00002_);
  and (_12693_[10], _12278_, _12276_);
  or (_12279_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_12280_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _12493_);
  or (_12281_, _12280_, _00002_);
  and (_12693_[11], _12281_, _12279_);
  or (_12282_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_12283_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _12493_);
  or (_12284_, _12283_, _00002_);
  and (_12693_[12], _12284_, _12282_);
  or (_12285_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_12286_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _12493_);
  or (_12287_, _12286_, _00002_);
  and (_12693_[13], _12287_, _12285_);
  or (_12288_, _11613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_12289_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _12493_);
  or (_12290_, _12289_, _00002_);
  and (_12693_[14], _12290_, _12288_);
  and (_12291_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nor (_12292_, _12166_, _11494_);
  or (_12293_, _12292_, _12291_);
  and (_12717_[0], _12293_, _12493_);
  and (_12294_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_12295_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_12296_, _12295_, _12166_);
  or (_12297_, _12296_, _12294_);
  and (_12717_[1], _12297_, _12493_);
  nor (_12298_, _12166_, _11529_);
  and (_12299_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_12300_, _12299_, _12166_);
  or (_12301_, _12300_, _12298_);
  and (_12717_[2], _12301_, _12493_);
  nor (_12302_, _12166_, _11547_);
  and (_12303_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_12304_, _12303_, _12166_);
  or (_12305_, _12304_, _12302_);
  and (_12717_[3], _12305_, _12493_);
  and (_12306_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_12307_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_12308_, _12307_, _12166_);
  or (_12309_, _12308_, _12306_);
  and (_12717_[4], _12309_, _12493_);
  and (_12310_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nor (_12311_, _12166_, _11582_);
  or (_12312_, _12311_, _12310_);
  and (_12717_[5], _12312_, _12493_);
  and (_12313_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nor (_12314_, _12166_, _11597_);
  or (_12315_, _12314_, _12313_);
  and (_12717_[6], _12315_, _12493_);
  nor (_12316_, _12166_, _11476_);
  and (_12317_, _12166_, _12144_);
  or (_12318_, _12317_, _12316_);
  and (_12717_[7], _12318_, _12493_);
  and (_12319_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_12320_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_12321_, _12320_, _12319_);
  and (_12717_[8], _12321_, _12493_);
  and (_12322_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_12323_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_12324_, _12323_, _12322_);
  and (_12717_[9], _12324_, _12493_);
  and (_12325_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_12326_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_12327_, _12326_, _12325_);
  and (_12717_[10], _12327_, _12493_);
  and (_12328_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_12329_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_12330_, _12329_, _12328_);
  and (_12717_[11], _12330_, _12493_);
  and (_12331_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_12332_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_12333_, _12332_, _12331_);
  and (_12717_[12], _12333_, _12493_);
  and (_12334_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_12335_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_12336_, _12335_, _12334_);
  and (_12717_[13], _12336_, _12493_);
  and (_12337_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_12338_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_12339_, _12338_, _12337_);
  and (_12717_[14], _12339_, _12493_);
  and (_12340_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_12341_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_12342_, _12341_, _12340_);
  and (_12717_[15], _12342_, _12493_);
  and (_12343_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_12344_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_12345_, _12344_, _12343_);
  and (_12717_[16], _12345_, _12493_);
  and (_12346_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_12347_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_12348_, _12347_, _12346_);
  and (_12717_[17], _12348_, _12493_);
  and (_12349_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_12350_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_12351_, _12350_, _12349_);
  and (_12717_[18], _12351_, _12493_);
  and (_12352_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_12353_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_12354_, _12353_, _12352_);
  and (_12717_[19], _12354_, _12493_);
  and (_12355_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_12356_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_12357_, _12356_, _12355_);
  and (_12717_[20], _12357_, _12493_);
  and (_12358_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_12359_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_12360_, _12359_, _12358_);
  and (_12717_[21], _12360_, _12493_);
  and (_12361_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_12362_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_12363_, _12362_, _12361_);
  and (_12717_[22], _12363_, _12493_);
  and (_12364_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_12365_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_12366_, _12365_, _12364_);
  and (_12717_[23], _12366_, _12493_);
  and (_12367_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_12368_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_12369_, _12368_, _12367_);
  and (_12717_[24], _12369_, _12493_);
  and (_12370_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_12371_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_12372_, _12371_, _12370_);
  and (_12717_[25], _12372_, _12493_);
  and (_12373_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_12374_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_12375_, _12374_, _12373_);
  and (_12717_[26], _12375_, _12493_);
  and (_12376_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_12377_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_12378_, _12377_, _12376_);
  and (_12717_[27], _12378_, _12493_);
  and (_12379_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_12380_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_12381_, _12380_, _12379_);
  and (_12717_[28], _12381_, _12493_);
  and (_12382_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_12383_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_12384_, _12383_, _12382_);
  and (_12717_[29], _12384_, _12493_);
  and (_12385_, _12166_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_12386_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_12387_, _12386_, _12385_);
  and (_12717_[30], _12387_, _12493_);
  nor (_12696_[0], _07360_, rst);
  nor (_12696_[1], _07438_, rst);
  nor (_12696_[2], _07386_, rst);
  nor (_12696_[3], _08883_, rst);
  and (_12697_[0], _09119_, _12493_);
  and (_12697_[1], _09279_, _12493_);
  and (_12697_[2], _08939_, _12493_);
  and (_12697_[3], _09167_, _12493_);
  and (_12697_[4], _09327_, _12493_);
  and (_12697_[5], _08996_, _12493_);
  and (_12697_[6], _09226_, _12493_);
  and (_12388_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0]);
  and (_12389_, _12695_, xram_data_in_reg[0]);
  or (_12702_[0], _12389_, _12388_);
  and (_12390_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1]);
  and (_12391_, _12695_, xram_data_in_reg[1]);
  or (_12702_[1], _12391_, _12390_);
  and (_12392_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2]);
  and (_12393_, _12695_, xram_data_in_reg[2]);
  or (_12702_[2], _12393_, _12392_);
  and (_12394_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3]);
  and (_12395_, _12695_, xram_data_in_reg[3]);
  or (_12702_[3], _12395_, _12394_);
  and (_12396_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4]);
  and (_12397_, _12695_, xram_data_in_reg[4]);
  or (_12702_[4], _12397_, _12396_);
  and (_12398_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5]);
  and (_12399_, _12695_, xram_data_in_reg[5]);
  or (_12702_[5], _12399_, _12398_);
  and (_12400_, _11726_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6]);
  and (_12401_, _12695_, xram_data_in_reg[6]);
  or (_12702_[6], _12401_, _12400_);
  or (_12402_, _11900_, _11897_);
  and (_12403_, _12402_, _06878_);
  and (_12404_, _07702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_12405_, _11754_, _11798_);
  and (_12406_, _11892_, _09141_);
  or (_12407_, _12406_, _12405_);
  or (_12408_, _12407_, _12404_);
  nor (_12409_, _11800_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_12410_, _12409_, _11801_);
  and (_12411_, _12410_, _11861_);
  or (_12412_, _12411_, _12408_);
  nor (_12413_, _12412_, _12403_);
  nand (_12414_, _12413_, _11876_);
  or (_12415_, _11876_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_12416_, _12415_, _12493_);
  and (_12703_[0], _12416_, _12414_);
  not (_12417_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_12418_, _11725_, _12417_);
  and (_12419_, _12402_, _06940_);
  or (_12420_, _11803_, _11801_);
  nor (_12421_, _11851_, _11755_);
  nor (_12422_, _11898_, _11760_);
  nor (_12423_, _12422_, _12421_);
  and (_12424_, _12423_, _11805_);
  and (_12425_, _12424_, _12420_);
  and (_12426_, _11754_, _11793_);
  and (_12427_, _12422_, _11891_);
  and (_12428_, _12427_, _09295_);
  or (_12429_, _12428_, _12426_);
  or (_12430_, _12429_, _12425_);
  or (_12431_, _12430_, _12419_);
  and (_12432_, _12431_, _11876_);
  or (_12433_, _12432_, _12418_);
  and (_12703_[1], _12433_, _12493_);
  not (_12434_, _11724_);
  not (_12435_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_12436_, _11731_, _12435_);
  and (_12437_, _11731_, _12435_);
  nor (_12438_, _12437_, _12436_);
  and (_12439_, _12438_, _12434_);
  and (_12440_, _12402_, _07001_);
  or (_12441_, _11808_, _11806_);
  and (_12442_, _12423_, _11810_);
  and (_12443_, _12442_, _12441_);
  and (_12444_, _11754_, _11788_);
  and (_12445_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_12446_, _12427_, _08969_);
  or (_12447_, _12446_, _12445_);
  or (_12448_, _12447_, _12444_);
  or (_12449_, _12448_, _12443_);
  or (_12450_, _12449_, _12440_);
  and (_12451_, _12450_, _11724_);
  or (_12452_, _12451_, _12439_);
  and (_12703_[2], _12452_, _12493_);
  and (_12453_, _12436_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_12454_, _12436_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_12455_, _12454_, _12453_);
  and (_12456_, _12455_, _12434_);
  and (_12457_, _12402_, _07065_);
  not (_12458_, _11811_);
  or (_12459_, _11785_, _11786_);
  nand (_12460_, _12459_, _12458_);
  or (_12461_, _12459_, _12458_);
  and (_12462_, _12461_, _12423_);
  and (_12463_, _12462_, _12460_);
  not (_12464_, _11555_);
  and (_12465_, _11754_, _12464_);
  and (_12466_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_12467_, _12427_, _09190_);
  or (_12468_, _12467_, _12466_);
  or (_12469_, _12468_, _12465_);
  or (_12470_, _12469_, _12463_);
  or (_12472_, _12470_, _12457_);
  and (_12474_, _12472_, _11724_);
  or (_12476_, _12474_, _12456_);
  and (_12703_[3], _12476_, _12493_);
  and (_12479_, _12436_, _11733_);
  nor (_12481_, _12453_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_12483_, _12481_, _12479_);
  nor (_12484_, _12483_, _11724_);
  and (_12485_, _12402_, _07135_);
  or (_12486_, _11815_, _11813_);
  and (_12487_, _12423_, _11816_);
  and (_12488_, _12487_, _12486_);
  not (_12489_, _11572_);
  and (_12491_, _11754_, _12489_);
  and (_12492_, _12427_, _09344_);
  and (_12494_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_12495_, _12494_, _12492_);
  or (_12496_, _12495_, _12491_);
  or (_12498_, _12496_, _12488_);
  or (_12499_, _12498_, _12485_);
  and (_12500_, _12499_, _11724_);
  or (_12502_, _12500_, _12484_);
  and (_12703_[4], _12502_, _12493_);
  and (_12503_, _12479_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12505_, _12479_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_12506_, _12505_, _12503_);
  nor (_12507_, _12506_, _11724_);
  and (_12509_, _12402_, _07213_);
  or (_12510_, _11776_, _11777_);
  and (_12511_, _12510_, _11817_);
  nor (_12513_, _12510_, _11817_);
  or (_12514_, _12513_, _12511_);
  and (_12515_, _12514_, _12423_);
  not (_12517_, _11590_);
  and (_12518_, _11754_, _12517_);
  and (_12519_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12521_, _12427_, _09015_);
  or (_12522_, _12521_, _12519_);
  or (_12523_, _12522_, _12518_);
  or (_12524_, _12523_, _12515_);
  or (_12525_, _12524_, _12509_);
  and (_12526_, _12525_, _11724_);
  or (_12527_, _12526_, _12507_);
  and (_12703_[5], _12527_, _12493_);
  and (_12528_, _12503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_12529_, _12503_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_12530_, _12529_, _12528_);
  nor (_12531_, _12530_, _11724_);
  and (_12532_, _12402_, _07286_);
  or (_12533_, _11819_, _11772_);
  and (_12534_, _12423_, _11820_);
  and (_12535_, _12534_, _12533_);
  not (_12536_, _11608_);
  and (_12537_, _11754_, _12536_);
  and (_12538_, _07620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12539_, _12427_, _09245_);
  or (_12540_, _12539_, _12538_);
  or (_12542_, _12540_, _12537_);
  or (_12543_, _12542_, _12535_);
  or (_12545_, _12543_, _12532_);
  and (_12546_, _12545_, _11724_);
  or (_12547_, _12546_, _12531_);
  and (_12703_[6], _12547_, _12493_);
  and (_12549_, _11737_, _11732_);
  nor (_12550_, _12528_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_12552_, _12550_, _12549_);
  nor (_12553_, _12552_, _11724_);
  or (_12554_, _11763_, _11764_);
  and (_12556_, _12554_, _11821_);
  nor (_12557_, _12554_, _11821_);
  or (_12558_, _12557_, _12556_);
  and (_12560_, _12558_, _11861_);
  and (_12561_, _12402_, _06771_);
  and (_12562_, _07702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_12564_, _11484_);
  and (_12565_, _11754_, _12564_);
  and (_12566_, _11892_, _09087_);
  or (_12568_, _12566_, _12565_);
  or (_12569_, _12568_, _12562_);
  or (_12570_, _12569_, _12561_);
  or (_12572_, _12570_, _12560_);
  and (_12573_, _12572_, _11724_);
  or (_12574_, _12573_, _12553_);
  and (_12703_[7], _12574_, _12493_);
  and (_12575_, _12549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_12576_, _12549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_12577_, _12576_, _12575_);
  or (_12578_, _12577_, _11724_);
  and (_12579_, _12578_, _12493_);
  and (_12580_, _11832_, _07919_);
  and (_12581_, _11823_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_12582_, _12581_, _12580_);
  nor (_12583_, _12582_, _11762_);
  and (_12584_, _12582_, _11762_);
  or (_12585_, _12584_, _12583_);
  and (_12586_, _12585_, _11861_);
  and (_12587_, _11897_, _07994_);
  and (_12588_, _11754_, _09141_);
  and (_12589_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12590_, _12427_, _10968_);
  or (_12591_, _12590_, _12589_);
  or (_12593_, _12591_, _12588_);
  or (_12594_, _12593_, _12587_);
  nor (_12596_, _07703_, _06877_);
  or (_12597_, _12596_, _12594_);
  nor (_12598_, _12597_, _12586_);
  nand (_12600_, _12598_, _11876_);
  and (_12703_[8], _12600_, _12579_);
  and (_12601_, _12575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_12603_, _12575_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_12604_, _12603_, _12601_);
  or (_12605_, _12604_, _11724_);
  and (_12607_, _12605_, _12493_);
  not (_12608_, _11762_);
  and (_00011_, _11832_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00013_, _00011_, _12608_);
  and (_00014_, _11824_, _11762_);
  nor (_00015_, _00014_, _00013_);
  nand (_00017_, _00015_, _07925_);
  or (_00018_, _00015_, _07925_);
  and (_00019_, _00018_, _12423_);
  and (_00021_, _00019_, _00017_);
  nor (_00022_, _11617_, _06939_);
  not (_00023_, _08024_);
  nand (_00025_, _11897_, _00023_);
  and (_00026_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_00027_, _11754_, _09295_);
  or (_00028_, _00027_, _00026_);
  and (_00029_, _12427_, _11011_);
  nor (_00030_, _00029_, _00028_);
  and (_00031_, _00030_, _00025_);
  nand (_00032_, _00031_, _11724_);
  or (_00033_, _00032_, _00022_);
  or (_00034_, _00033_, _00021_);
  and (_12703_[9], _00034_, _12607_);
  nor (_00035_, _12601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00036_, _12601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00037_, _00036_, _00035_);
  or (_00038_, _00037_, _11724_);
  and (_00039_, _00038_, _12493_);
  and (_00040_, _00014_, _07925_);
  and (_00041_, _00013_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_00042_, _00041_, _00040_);
  nand (_00043_, _00042_, _07930_);
  or (_00044_, _00042_, _07930_);
  and (_00046_, _00044_, _12423_);
  and (_00047_, _00046_, _00043_);
  nor (_00049_, _11617_, _07000_);
  not (_00050_, _11897_);
  or (_00051_, _00050_, _08055_);
  and (_00053_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_00054_, _11754_, _08969_);
  and (_00055_, _12427_, _10951_);
  or (_00057_, _00055_, _00054_);
  nor (_00058_, _00057_, _00053_);
  and (_00059_, _00058_, _00051_);
  nand (_00061_, _00059_, _11724_);
  or (_00062_, _00061_, _00049_);
  or (_00063_, _00062_, _00047_);
  and (_12703_[10], _00063_, _00039_);
  nand (_00065_, _12601_, _11738_);
  or (_00066_, _00036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_00068_, _00066_, _00065_);
  or (_00069_, _00068_, _11724_);
  and (_00070_, _00069_, _12493_);
  and (_00072_, _11835_, _12608_);
  not (_00073_, _00072_);
  or (_00074_, _11826_, _12608_);
  and (_00076_, _00074_, _00073_);
  or (_00077_, _00076_, _07915_);
  nand (_00078_, _00076_, _07915_);
  and (_00079_, _00078_, _12423_);
  and (_00080_, _00079_, _00077_);
  and (_00081_, _07620_, _07065_);
  or (_00082_, _00050_, _08085_);
  and (_00083_, _11754_, _09190_);
  and (_00084_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_00085_, _11883_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_00086_, _00085_, _11884_);
  and (_00087_, _00086_, _12427_);
  or (_00088_, _00087_, _00084_);
  nor (_00089_, _00088_, _00083_);
  and (_00090_, _00089_, _00082_);
  nand (_00091_, _00090_, _11724_);
  or (_00092_, _00091_, _00081_);
  or (_00093_, _00092_, _00080_);
  and (_12703_[11], _00093_, _00070_);
  nor (_00094_, _11742_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00095_, _00094_, _11743_);
  or (_00097_, _00095_, _11724_);
  and (_00098_, _00097_, _12493_);
  and (_00100_, _11836_, _12608_);
  not (_00101_, _00100_);
  nand (_00102_, _11827_, _11762_);
  and (_00104_, _00102_, _00101_);
  nand (_00105_, _00104_, _07936_);
  or (_00106_, _00104_, _07936_);
  and (_00108_, _00106_, _12423_);
  and (_00109_, _00108_, _00105_);
  nor (_00110_, _11617_, _07134_);
  or (_00112_, _00050_, _08117_);
  and (_00113_, _11754_, _09344_);
  and (_00114_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_00116_, _11884_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_00117_, _00116_, _11885_);
  and (_00118_, _00117_, _12427_);
  or (_00120_, _00118_, _00114_);
  nor (_00121_, _00120_, _00113_);
  and (_00122_, _00121_, _00112_);
  nand (_00124_, _00122_, _11724_);
  or (_00125_, _00124_, _00110_);
  or (_00126_, _00125_, _00109_);
  and (_12703_[12], _00126_, _00098_);
  not (_00128_, _11876_);
  nand (_00129_, _00100_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_00130_, _00102_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_00131_, _00130_, _00129_);
  and (_00132_, _00131_, _07911_);
  nor (_00133_, _00131_, _07911_);
  or (_00134_, _00133_, _00132_);
  and (_00135_, _00134_, _12423_);
  and (_00136_, _07620_, _07213_);
  nor (_00137_, _00050_, _08150_);
  and (_00138_, _11754_, _09015_);
  and (_00139_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00140_, _11885_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00141_, _00140_, _11886_);
  and (_00142_, _00141_, _12427_);
  or (_00143_, _00142_, _00139_);
  or (_00144_, _00143_, _00138_);
  or (_00145_, _00144_, _00137_);
  or (_00146_, _00145_, _00136_);
  or (_00147_, _00146_, _00135_);
  or (_00149_, _00147_, _00128_);
  nor (_00150_, _11743_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_00152_, _00150_, _11744_);
  or (_00153_, _00152_, _11876_);
  and (_00154_, _00153_, _12493_);
  and (_12703_[13], _00154_, _00149_);
  nor (_00156_, _11617_, _07285_);
  nor (_00157_, _00050_, _08180_);
  and (_00159_, _11900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_00160_, _11754_, _09245_);
  or (_00161_, _00160_, _00159_);
  or (_00163_, _11886_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00164_, _00163_, _11887_);
  and (_00165_, _00164_, _12427_);
  or (_00167_, _00165_, _00161_);
  or (_00168_, _00167_, _00157_);
  or (_00169_, _00168_, _00156_);
  nor (_00171_, _11762_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00172_, _11762_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_00173_, _00172_, _00171_);
  and (_00175_, _00173_, _00131_);
  nor (_00176_, _00175_, _07942_);
  and (_00177_, _00175_, _07942_);
  or (_00179_, _00177_, _00176_);
  and (_00180_, _00179_, _12423_);
  or (_00181_, _00180_, _00169_);
  or (_00182_, _00181_, _00128_);
  nor (_00183_, _11744_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_00184_, _00183_, _11745_);
  or (_00185_, _00184_, _11876_);
  and (_00186_, _00185_, _12493_);
  and (_12703_[14], _00186_, _00182_);
  and (_00187_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_00188_, _12080_, _12078_);
  nor (_00189_, _00188_, _12081_);
  or (_00190_, _00189_, _11912_);
  or (_00191_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_00192_, _00191_, _12112_);
  and (_00193_, _00192_, _00190_);
  or (_12704_[0], _00193_, _00187_);
  and (_00194_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00195_, _12083_, _12081_);
  and (_00196_, _00195_, _12084_);
  or (_00197_, _00196_, _11912_);
  or (_00199_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00200_, _00199_, _12112_);
  and (_00202_, _00200_, _00197_);
  or (_12704_[1], _00202_, _00194_);
  and (_00203_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00205_, _12088_, _12086_);
  nor (_00206_, _00205_, _12089_);
  or (_00207_, _00206_, _11912_);
  or (_00209_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00210_, _00209_, _12112_);
  and (_00211_, _00210_, _00207_);
  or (_12704_[2], _00211_, _00203_);
  nor (_00213_, _12089_, _11981_);
  nor (_00214_, _00213_, _12090_);
  or (_00216_, _00214_, _11912_);
  or (_00217_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00218_, _00217_, _12112_);
  and (_00220_, _00218_, _00216_);
  and (_00221_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_12704_[3], _00221_, _00220_);
  nor (_00223_, _12093_, _12090_);
  nor (_00224_, _00223_, _12094_);
  or (_00225_, _00224_, _11912_);
  or (_00227_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00228_, _00227_, _12112_);
  and (_00229_, _00228_, _00225_);
  and (_00230_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_12704_[4], _00230_, _00229_);
  and (_00231_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00232_, _12094_, _11976_);
  nor (_00233_, _00232_, _12095_);
  or (_00234_, _00233_, _11912_);
  or (_00235_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00236_, _00235_, _12112_);
  and (_00237_, _00236_, _00234_);
  or (_12704_[5], _00237_, _00231_);
  and (_00238_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00239_, _12095_, _11972_);
  nor (_00240_, _00239_, _12096_);
  or (_00241_, _00240_, _11912_);
  or (_00242_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00243_, _00242_, _12112_);
  and (_00244_, _00243_, _00241_);
  or (_12704_[6], _00244_, _00238_);
  or (_00246_, _12096_, _11968_);
  nor (_00247_, _12097_, _11912_);
  and (_00249_, _00247_, _00246_);
  nor (_00250_, _11911_, _05852_);
  or (_00251_, _00250_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00253_, _00251_, _00249_);
  or (_00254_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _07309_);
  and (_00255_, _00254_, _12493_);
  and (_12704_[7], _00255_, _00253_);
  nor (_00257_, _12099_, _12097_);
  nor (_00258_, _00257_, _12100_);
  or (_00260_, _00258_, _11912_);
  or (_00261_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00262_, _00261_, _12112_);
  and (_00264_, _00262_, _00260_);
  and (_00265_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_12704_[8], _00265_, _00264_);
  nor (_00267_, _12100_, _11965_);
  nor (_00268_, _00267_, _12101_);
  or (_00269_, _00268_, _11912_);
  or (_00271_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00272_, _00271_, _12112_);
  and (_00273_, _00272_, _00269_);
  and (_00275_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_12704_[9], _00275_, _00273_);
  nor (_00276_, _12101_, _11963_);
  nor (_00277_, _00276_, _12102_);
  or (_00278_, _00277_, _11912_);
  or (_00279_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00280_, _00279_, _12112_);
  and (_00281_, _00280_, _00278_);
  and (_00282_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_12704_[10], _00282_, _00281_);
  nor (_00283_, _12102_, _11960_);
  nor (_00284_, _00283_, _12103_);
  or (_00285_, _00284_, _11912_);
  or (_00286_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00287_, _00286_, _12112_);
  and (_00288_, _00287_, _00285_);
  and (_00289_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_12704_[11], _00289_, _00288_);
  nor (_00290_, _12103_, _11957_);
  nor (_00291_, _00290_, _12104_);
  or (_00292_, _00291_, _11912_);
  or (_00294_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00295_, _00294_, _12112_);
  and (_00297_, _00295_, _00292_);
  and (_00298_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_12704_[12], _00298_, _00297_);
  nor (_00300_, _12104_, _11954_);
  nor (_00301_, _00300_, _12105_);
  or (_00302_, _00301_, _11912_);
  or (_00304_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00305_, _00304_, _12112_);
  and (_00306_, _00305_, _00302_);
  and (_00308_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_12704_[13], _00308_, _00306_);
  nor (_00309_, _12105_, _11952_);
  nor (_00311_, _00309_, _12106_);
  or (_00312_, _00311_, _11912_);
  or (_00313_, _11911_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_00315_, _00313_, _12112_);
  and (_00316_, _00315_, _00312_);
  and (_00317_, _11908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_12704_[14], _00317_, _00316_);
  and (_12708_[0], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12493_);
  and (_12708_[1], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12493_);
  and (_12708_[2], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _12493_);
  and (_12708_[3], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12493_);
  and (_12708_[4], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12493_);
  and (_12708_[5], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _12493_);
  and (_12708_[6], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _12493_);
  nor (_00320_, _12077_, _08951_);
  nand (_00321_, _00320_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00322_, _00320_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00323_, _00322_, _12112_);
  and (_12709_[0], _00323_, _00321_);
  or (_00324_, _12122_, _12120_);
  and (_00325_, _00324_, _12123_);
  or (_00326_, _00325_, _08951_);
  or (_00327_, _07312_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00328_, _00327_, _12112_);
  and (_12709_[1], _00328_, _00326_);
  and (_00329_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_00330_, _00329_, _12143_);
  or (_00331_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00332_, _00331_, _12493_);
  and (_12713_[0], _00332_, _00330_);
  or (_00334_, _12295_, _12143_);
  or (_00335_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00337_, _00335_, _12493_);
  and (_12713_[1], _00337_, _00334_);
  or (_00338_, _12299_, _12143_);
  or (_00340_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00341_, _00340_, _12493_);
  and (_12713_[2], _00341_, _00338_);
  or (_00343_, _12303_, _12143_);
  or (_00344_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00345_, _00344_, _12493_);
  and (_12713_[3], _00345_, _00343_);
  or (_00347_, _12307_, _12143_);
  or (_00348_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00350_, _00348_, _12493_);
  and (_12713_[4], _00350_, _00347_);
  and (_00351_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_00353_, _00351_, _12143_);
  or (_00354_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00355_, _00354_, _12493_);
  and (_12713_[5], _00355_, _00353_);
  and (_00357_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_00358_, _00357_, _12143_);
  or (_00360_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00361_, _00360_, _12493_);
  and (_12713_[6], _00361_, _00358_);
  and (_12716_[0], _12152_, _12493_);
  nor (_12716_[1], _12162_, rst);
  and (_12716_[2], _12158_, _12493_);
  or (_00362_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand (_00363_, _12166_, _11494_);
  and (_00364_, _00363_, _12493_);
  and (_12718_[0], _00364_, _00362_);
  and (_00365_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00366_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00367_, _00366_, _00365_);
  and (_12718_[1], _00367_, _12493_);
  or (_00368_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_00369_, _12166_, _11529_);
  and (_00370_, _00369_, _12493_);
  and (_12718_[2], _00370_, _00368_);
  or (_00371_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_00372_, _12166_, _11547_);
  and (_00373_, _00372_, _12493_);
  and (_12718_[3], _00373_, _00371_);
  and (_00375_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00377_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00378_, _00377_, _00375_);
  and (_12718_[4], _00378_, _12493_);
  or (_00380_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_00381_, _12166_, _11582_);
  and (_00382_, _00381_, _12493_);
  and (_12718_[5], _00382_, _00380_);
  or (_00384_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_00385_, _12166_, _11597_);
  and (_00387_, _00385_, _12493_);
  and (_12718_[6], _00387_, _00384_);
  or (_00388_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_00390_, _12166_, _11476_);
  and (_00391_, _00390_, _12493_);
  and (_12718_[7], _00391_, _00388_);
  and (_00393_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_00394_, _12166_, _07326_);
  or (_00395_, _00394_, _00393_);
  and (_12718_[8], _00395_, _12493_);
  and (_00397_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00398_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00400_, _00398_, _00397_);
  and (_12718_[9], _00400_, _12493_);
  and (_00401_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_00402_, _12166_, _07363_);
  or (_00403_, _00402_, _00401_);
  and (_12718_[10], _00403_, _12493_);
  and (_00404_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_00405_, _12166_, _07391_);
  or (_00406_, _00405_, _00404_);
  and (_12718_[11], _00406_, _12493_);
  and (_00407_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00408_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00409_, _00408_, _00407_);
  and (_12718_[12], _00409_, _12493_);
  and (_00410_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_00411_, _12166_, _07505_);
  or (_00412_, _00411_, _00410_);
  and (_12718_[13], _00412_, _12493_);
  and (_00413_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_00414_, _12166_, _07471_);
  or (_00415_, _00414_, _00413_);
  and (_12718_[14], _00415_, _12493_);
  and (_00417_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_00419_, _12166_, _07445_);
  or (_00420_, _00419_, _00417_);
  and (_12718_[15], _00420_, _12493_);
  and (_00422_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_00423_, _12166_, _07320_);
  or (_00424_, _00423_, _00422_);
  and (_12718_[16], _00424_, _12493_);
  and (_00426_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00427_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00429_, _00427_, _00426_);
  and (_12718_[17], _00429_, _12493_);
  and (_00430_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_00432_, _12166_, _07365_);
  or (_00433_, _00432_, _00430_);
  and (_12718_[18], _00433_, _12493_);
  and (_00435_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_00436_, _12166_, _07389_);
  or (_00437_, _00436_, _00435_);
  and (_12718_[19], _00437_, _12493_);
  and (_00439_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_00440_, _12166_, _07530_);
  or (_00442_, _00440_, _00439_);
  and (_12718_[20], _00442_, _12493_);
  and (_00443_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_00444_, _12166_, _07498_);
  or (_00445_, _00444_, _00443_);
  and (_12718_[21], _00445_, _12493_);
  and (_00446_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_00447_, _12166_, _07475_);
  or (_00448_, _00447_, _00446_);
  and (_12718_[22], _00448_, _12493_);
  and (_00449_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_00450_, _12166_, _07449_);
  or (_00451_, _00450_, _00449_);
  and (_12718_[23], _00451_, _12493_);
  and (_00452_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_00453_, _12166_, _09130_);
  or (_00454_, _00453_, _00452_);
  and (_12718_[24], _00454_, _12493_);
  and (_00455_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00456_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00457_, _00456_, _00455_);
  and (_12718_[25], _00457_, _12493_);
  and (_00459_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor (_00461_, _12166_, _08959_);
  or (_00462_, _00461_, _00459_);
  and (_12718_[26], _00462_, _12493_);
  and (_00464_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_00465_, _12166_, _09177_);
  or (_00466_, _00465_, _00464_);
  and (_12718_[27], _00466_, _12493_);
  and (_00468_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00469_, _12168_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00471_, _00469_, _00468_);
  and (_12718_[28], _00471_, _12493_);
  and (_00472_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_00474_, _12166_, _09008_);
  or (_00475_, _00474_, _00472_);
  and (_12718_[29], _00475_, _12493_);
  and (_00477_, _12166_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_00478_, _12166_, _09238_);
  or (_00479_, _00478_, _00477_);
  and (_12718_[30], _00479_, _12493_);
  not (_00481_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  nor (_00482_, _12175_, _00481_);
  and (_00484_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00485_, _00484_, _12175_);
  or (_00486_, _00485_, _00482_);
  and (_12719_[0], _00486_, _12493_);
  not (_00487_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  nor (_00488_, _12175_, _00487_);
  and (_00489_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00490_, _00489_, _12175_);
  or (_00491_, _00490_, _00488_);
  and (_12719_[1], _00491_, _12493_);
  not (_00492_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  nor (_00493_, _12175_, _00492_);
  and (_00494_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00495_, _00494_, _12175_);
  or (_00496_, _00495_, _00493_);
  and (_12719_[2], _00496_, _12493_);
  not (_00497_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  nor (_00498_, _12175_, _00497_);
  and (_00499_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00500_, _00499_, _12175_);
  or (_00501_, _00500_, _00498_);
  and (_12719_[3], _00501_, _12493_);
  not (_00503_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  nor (_00505_, _12175_, _00503_);
  and (_00506_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00507_, _00506_, _12175_);
  or (_00509_, _00507_, _00505_);
  and (_12719_[4], _00509_, _12493_);
  not (_00510_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  nor (_00512_, _12175_, _00510_);
  and (_00513_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_00514_, _00513_, _12175_);
  or (_00516_, _00514_, _00512_);
  and (_12719_[5], _00516_, _12493_);
  not (_00517_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  nor (_00519_, _12175_, _00517_);
  and (_00520_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00521_, _00520_, _12175_);
  or (_00523_, _00521_, _00519_);
  and (_12719_[6], _00523_, _12493_);
  not (_00524_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  nor (_00526_, _12175_, _00524_);
  or (_00527_, _09119_, _12186_);
  or (_00528_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00530_, _00528_, _12175_);
  and (_00531_, _00530_, _00527_);
  or (_00532_, _00531_, _00526_);
  and (_12722_[0], _00532_, _12493_);
  not (_00533_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  nor (_00534_, _12175_, _00533_);
  or (_00535_, _09279_, _12186_);
  or (_00536_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00537_, _00536_, _12175_);
  and (_00538_, _00537_, _00535_);
  or (_00539_, _00538_, _00534_);
  and (_12722_[1], _00539_, _12493_);
  not (_00540_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  nor (_00541_, _12175_, _00540_);
  or (_00542_, _08939_, _12186_);
  or (_00543_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00544_, _00543_, _12175_);
  and (_00545_, _00544_, _00542_);
  or (_00546_, _00545_, _00541_);
  and (_12722_[2], _00546_, _12493_);
  not (_00547_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  nor (_00548_, _12175_, _00547_);
  or (_00549_, _09167_, _12186_);
  or (_00551_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00552_, _00551_, _12175_);
  and (_00553_, _00552_, _00549_);
  or (_00554_, _00553_, _00548_);
  and (_12722_[3], _00554_, _12493_);
  not (_00555_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  nor (_00556_, _12175_, _00555_);
  or (_00557_, _09327_, _12186_);
  or (_00558_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00559_, _00558_, _12175_);
  and (_00560_, _00559_, _00557_);
  or (_00561_, _00560_, _00556_);
  and (_12722_[4], _00561_, _12493_);
  not (_00562_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  nor (_00563_, _12175_, _00562_);
  or (_00564_, _08996_, _12186_);
  or (_00565_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00566_, _00565_, _12175_);
  and (_00567_, _00566_, _00564_);
  or (_00568_, _00567_, _00563_);
  and (_12722_[5], _00568_, _12493_);
  not (_00569_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  nor (_00570_, _12175_, _00569_);
  or (_00571_, _09226_, _12186_);
  or (_00572_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00573_, _00572_, _12175_);
  and (_00574_, _00573_, _00571_);
  or (_00575_, _00574_, _00570_);
  and (_12722_[6], _00575_, _12493_);
  not (_00576_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  nor (_00577_, _12175_, _00576_);
  or (_00578_, _09069_, _12186_);
  or (_00579_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00580_, _00579_, _12175_);
  and (_00581_, _00580_, _00578_);
  or (_00582_, _00581_, _00577_);
  and (_12722_[7], _00582_, _12493_);
  not (_00583_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  nor (_00584_, _12175_, _00583_);
  and (_00585_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_00586_, _00585_, _12175_);
  or (_00587_, _00586_, _00584_);
  and (_12722_[8], _00587_, _12493_);
  not (_00588_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  nor (_00589_, _12175_, _00588_);
  and (_00590_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_00591_, _00590_, _12175_);
  or (_00592_, _00591_, _00589_);
  and (_12722_[9], _00592_, _12493_);
  not (_00593_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  nor (_00594_, _12175_, _00593_);
  and (_00595_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_00596_, _00595_, _12175_);
  or (_00597_, _00596_, _00594_);
  and (_12722_[10], _00597_, _12493_);
  not (_00598_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  nor (_00599_, _12175_, _00598_);
  and (_00600_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_00601_, _00600_, _12175_);
  or (_00602_, _00601_, _00599_);
  and (_12722_[11], _00602_, _12493_);
  not (_00603_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  nor (_00604_, _12175_, _00603_);
  and (_00605_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_00606_, _00605_, _12175_);
  or (_00607_, _00606_, _00604_);
  and (_12722_[12], _00607_, _12493_);
  not (_00608_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  nor (_00609_, _12175_, _00608_);
  and (_00610_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_00611_, _00610_, _12175_);
  or (_00612_, _00611_, _00609_);
  and (_12722_[13], _00612_, _12493_);
  not (_00613_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  nor (_00614_, _12175_, _00613_);
  and (_00615_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_00616_, _00615_, _12175_);
  or (_00617_, _00616_, _00614_);
  and (_12722_[14], _00617_, _12493_);
  nand (_00618_, _12192_, _06877_);
  or (_00619_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00620_, _00619_, _12493_);
  and (_12726_[0], _00620_, _00618_);
  nand (_00621_, _12192_, _06939_);
  or (_00622_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00623_, _00622_, _12493_);
  and (_12726_[1], _00623_, _00621_);
  nand (_00624_, _12192_, _07000_);
  or (_00625_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00626_, _00625_, _12493_);
  and (_12726_[2], _00626_, _00624_);
  or (_00627_, _12197_, _07065_);
  or (_00628_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00629_, _00628_, _12493_);
  and (_12726_[3], _00629_, _00627_);
  nand (_00630_, _12192_, _07134_);
  or (_00631_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00632_, _00631_, _12493_);
  and (_12726_[4], _00632_, _00630_);
  or (_00633_, _12197_, _07213_);
  or (_00634_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00635_, _00634_, _12493_);
  and (_12726_[5], _00635_, _00633_);
  nand (_00636_, _12192_, _07285_);
  or (_00637_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00638_, _00637_, _12493_);
  and (_12726_[6], _00638_, _00636_);
  nand (_00639_, _12192_, _06770_);
  or (_00640_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00641_, _00640_, _12493_);
  and (_12726_[7], _00641_, _00639_);
  or (_00642_, _12197_, _07994_);
  or (_00643_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00644_, _00643_, _12493_);
  and (_12726_[8], _00644_, _00642_);
  nand (_00645_, _12192_, _08024_);
  or (_00646_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00647_, _00646_, _12493_);
  and (_12726_[9], _00647_, _00645_);
  nand (_00648_, _12192_, _08055_);
  or (_00649_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00650_, _00649_, _12493_);
  and (_12726_[10], _00650_, _00648_);
  nand (_00651_, _12192_, _08085_);
  or (_00652_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00653_, _00652_, _12493_);
  and (_12726_[11], _00653_, _00651_);
  nand (_00654_, _12192_, _08117_);
  or (_00655_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00656_, _00655_, _12493_);
  and (_12726_[12], _00656_, _00654_);
  nand (_00657_, _12192_, _08150_);
  or (_00658_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00659_, _00658_, _12493_);
  and (_12726_[13], _00659_, _00657_);
  nand (_00660_, _12192_, _08180_);
  or (_00661_, _12192_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00662_, _00661_, _12493_);
  and (_12726_[14], _00662_, _00660_);
  nor (_12691_, _08868_, rst);
  nor (_00663_, _09250_, _09092_);
  and (_00664_, _09355_, _09023_);
  and (_00665_, _00664_, _09194_);
  and (_00666_, _00665_, _00663_);
  not (_00667_, _08973_);
  or (_00668_, _08365_, _08353_);
  nand (_00669_, _08365_, _08353_);
  nand (_00670_, _00669_, _00668_);
  nand (_00671_, _08376_, _08374_);
  nand (_00672_, _08394_, _00671_);
  or (_00673_, _08394_, _00671_);
  and (_00674_, _00673_, _00672_);
  nand (_00675_, _00674_, _00670_);
  or (_00676_, _00674_, _00670_);
  nand (_00677_, _00676_, _00675_);
  nand (_00678_, _08419_, _08406_);
  or (_00679_, _08419_, _08406_);
  nand (_00680_, _00679_, _00678_);
  nand (_00681_, _08341_, _08340_);
  or (_00682_, _08431_, _00681_);
  nand (_00683_, _08430_, _08428_);
  or (_00684_, _00683_, _08342_);
  and (_00685_, _00684_, _00682_);
  nand (_00686_, _00685_, _00680_);
  or (_00687_, _00685_, _00680_);
  nand (_00688_, _00687_, _00686_);
  nand (_00689_, _00688_, _00677_);
  or (_00690_, _00688_, _00677_);
  and (_00691_, _00690_, _00689_);
  or (_00692_, _00691_, _00667_);
  and (_00693_, _09145_, _09304_);
  or (_00694_, _08973_, _08287_);
  and (_00695_, _00694_, _00693_);
  and (_00696_, _00695_, _00692_);
  nor (_00697_, _09145_, _09304_);
  and (_00698_, _00697_, _00667_);
  and (_00699_, _00698_, _08225_);
  and (_00700_, _00697_, _08973_);
  and (_00701_, _00700_, _08276_);
  or (_00702_, _08973_, _08296_);
  not (_00703_, _09145_);
  and (_00704_, _00703_, _09304_);
  or (_00705_, _00667_, _08233_);
  and (_00706_, _00705_, _00704_);
  and (_00707_, _00706_, _00702_);
  or (_00708_, _00707_, _00701_);
  or (_00709_, _00708_, _00699_);
  or (_00710_, _00667_, _08269_);
  nor (_00711_, _00703_, _09304_);
  or (_00712_, _08973_, _08312_);
  and (_00713_, _00712_, _00711_);
  and (_00714_, _00713_, _00710_);
  or (_00715_, _00714_, _00709_);
  or (_00716_, _00715_, _00696_);
  and (_00717_, _00716_, _00666_);
  and (_00718_, _07579_, _07643_);
  not (_00719_, _00718_);
  nor (_00720_, _11085_, _07642_);
  and (_00721_, _00720_, _00719_);
  nor (_00722_, _07690_, _07686_);
  and (_00723_, _00722_, _00721_);
  nor (_00724_, _11151_, _11086_);
  and (_00725_, _00724_, _00723_);
  and (_00726_, _07555_, _07525_);
  not (_00727_, _00726_);
  and (_00728_, _07637_, _07643_);
  nor (_00729_, _11261_, _00728_);
  and (_00730_, _00729_, _00727_);
  and (_00731_, _00730_, _11429_);
  and (_00732_, _00731_, _00725_);
  and (_00733_, _00732_, _07682_);
  nor (_00734_, _00733_, _07308_);
  or (_00735_, _11609_, p2in_reg[6]);
  or (_00736_, _11613_, p2_in[6]);
  and (_00737_, _00736_, _00735_);
  or (_00738_, _00737_, _00734_);
  not (_00739_, _00734_);
  or (_00740_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_00741_, _00740_, _00738_);
  and (_00742_, _00741_, _00667_);
  or (_00743_, _11609_, p2in_reg[2]);
  or (_00744_, _11613_, p2_in[2]);
  and (_00745_, _00744_, _00743_);
  or (_00746_, _00745_, _00734_);
  nand (_00747_, _00734_, _08703_);
  and (_00748_, _00747_, _00746_);
  and (_00749_, _00748_, _08973_);
  or (_00750_, _00749_, _00742_);
  and (_00751_, _00750_, _00711_);
  or (_00752_, _11609_, p2in_reg[3]);
  or (_00753_, _11613_, p2_in[3]);
  and (_00754_, _00753_, _00752_);
  or (_00755_, _00754_, _00734_);
  or (_00756_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00757_, _00756_, _00755_);
  and (_00758_, _00757_, _00700_);
  or (_00759_, _00758_, _00751_);
  or (_00760_, _11609_, p2in_reg[7]);
  or (_00761_, _11613_, p2_in[7]);
  and (_00762_, _00761_, _00760_);
  or (_00763_, _00762_, _00734_);
  nand (_00764_, _00734_, _08473_);
  and (_00765_, _00764_, _00763_);
  and (_00766_, _00765_, _00698_);
  or (_00767_, _11609_, p2in_reg[5]);
  or (_00768_, _11613_, p2_in[5]);
  and (_00769_, _00768_, _00767_);
  or (_00770_, _00769_, _00734_);
  or (_00771_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00772_, _00771_, _00770_);
  and (_00773_, _00772_, _00667_);
  or (_00774_, _11609_, p2in_reg[1]);
  or (_00775_, _11613_, p2_in[1]);
  and (_00776_, _00775_, _00774_);
  or (_00777_, _00776_, _00734_);
  or (_00778_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_00779_, _00778_, _00777_);
  and (_00780_, _00779_, _08973_);
  or (_00781_, _00780_, _00773_);
  and (_00782_, _00781_, _00704_);
  or (_00783_, _11609_, p2in_reg[4]);
  or (_00784_, _11613_, p2_in[4]);
  and (_00785_, _00784_, _00783_);
  or (_00786_, _00785_, _00734_);
  or (_00787_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00788_, _00787_, _00786_);
  or (_00789_, _00788_, _08973_);
  or (_00790_, _11609_, p2in_reg[0]);
  or (_00791_, _11613_, p2_in[0]);
  and (_00792_, _00791_, _00790_);
  or (_00793_, _00792_, _00734_);
  or (_00794_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_00795_, _00794_, _00793_);
  or (_00796_, _00795_, _00667_);
  and (_00797_, _00796_, _00693_);
  and (_00798_, _00797_, _00789_);
  or (_00799_, _00798_, _00782_);
  or (_00800_, _00799_, _00766_);
  or (_00801_, _00800_, _00759_);
  nor (_00802_, _09195_, _09092_);
  and (_00803_, _00802_, _09354_);
  not (_00804_, _09250_);
  nor (_00805_, _00804_, _09023_);
  and (_00806_, _00805_, _00803_);
  and (_00807_, _00806_, _00801_);
  nor (_00808_, _09250_, _09023_);
  and (_00809_, _00802_, _09355_);
  and (_00810_, _00809_, _00808_);
  or (_00811_, _08973_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_00812_, _08973_, _06880_);
  and (_00813_, _00812_, _00693_);
  and (_00814_, _00813_, _00811_);
  and (_00815_, _00700_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00816_, _00815_, _00814_);
  and (_00817_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_00818_, _08973_, _07288_);
  and (_00819_, _08973_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00820_, _00819_, _00818_);
  and (_00821_, _00820_, _00711_);
  nor (_00822_, _08973_, _07215_);
  and (_00823_, _08973_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00824_, _00823_, _00822_);
  and (_00825_, _00824_, _00704_);
  or (_00826_, _00825_, _00821_);
  or (_00827_, _00826_, _00817_);
  or (_00828_, _00827_, _00816_);
  and (_00829_, _00828_, _00810_);
  or (_00830_, _11609_, p1in_reg[5]);
  or (_00831_, _11613_, p1_in[5]);
  and (_00832_, _00831_, _00830_);
  or (_00833_, _00832_, _00734_);
  or (_00834_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00835_, _00834_, _00833_);
  and (_00836_, _00835_, _00667_);
  or (_00837_, _11609_, p1in_reg[1]);
  or (_00838_, _11613_, p1_in[1]);
  and (_00839_, _00838_, _00837_);
  or (_00840_, _00839_, _00734_);
  or (_00841_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_00842_, _00841_, _00840_);
  and (_00843_, _00842_, _08973_);
  or (_00844_, _00843_, _00836_);
  and (_00845_, _00844_, _00704_);
  or (_00846_, _11609_, p1in_reg[4]);
  or (_00847_, _11613_, p1_in[4]);
  and (_00848_, _00847_, _00846_);
  or (_00849_, _00848_, _00734_);
  or (_00850_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00851_, _00850_, _00849_);
  or (_00852_, _00851_, _08973_);
  or (_00853_, _11609_, p1in_reg[0]);
  or (_00854_, _11613_, p1_in[0]);
  and (_00855_, _00854_, _00853_);
  or (_00856_, _00855_, _00734_);
  or (_00857_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_00858_, _00857_, _00856_);
  or (_00859_, _00858_, _00667_);
  and (_00860_, _00859_, _00693_);
  and (_00861_, _00860_, _00852_);
  or (_00862_, _00861_, _00845_);
  or (_00863_, _11609_, p1in_reg[6]);
  or (_00864_, _11613_, p1_in[6]);
  and (_00865_, _00864_, _00863_);
  or (_00866_, _00865_, _00734_);
  or (_00867_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_00868_, _00867_, _00866_);
  and (_00869_, _00868_, _00667_);
  or (_00870_, _11609_, p1in_reg[2]);
  or (_00871_, _11613_, p1_in[2]);
  and (_00872_, _00871_, _00870_);
  or (_00873_, _00872_, _00734_);
  nand (_00874_, _00734_, _08618_);
  and (_00875_, _00874_, _00873_);
  and (_00876_, _00875_, _08973_);
  or (_00877_, _00876_, _00869_);
  and (_00878_, _00877_, _00711_);
  or (_00879_, _11609_, p1in_reg[7]);
  or (_00880_, _11613_, p1_in[7]);
  and (_00881_, _00880_, _00879_);
  or (_00882_, _00881_, _00734_);
  nand (_00883_, _00734_, _08453_);
  and (_00884_, _00883_, _00882_);
  and (_00885_, _00884_, _00698_);
  or (_00886_, _11609_, p1in_reg[3]);
  or (_00887_, _11613_, p1_in[3]);
  and (_00888_, _00887_, _00886_);
  or (_00889_, _00888_, _00734_);
  or (_00890_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00891_, _00890_, _00889_);
  and (_00892_, _00891_, _00700_);
  or (_00893_, _00892_, _00885_);
  or (_00894_, _00893_, _00878_);
  or (_00895_, _00894_, _00862_);
  nor (_00896_, _00804_, _09092_);
  and (_00897_, _00896_, _00665_);
  and (_00898_, _00897_, _00895_);
  or (_00899_, _00898_, _00829_);
  or (_00900_, _00899_, _00807_);
  or (_00901_, _11609_, p3in_reg[6]);
  or (_00902_, _11613_, p3_in[6]);
  and (_00903_, _00902_, _00901_);
  or (_00904_, _00903_, _00734_);
  or (_00905_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_00906_, _00905_, _00904_);
  and (_00907_, _00906_, _00667_);
  or (_00908_, _11609_, p3in_reg[2]);
  or (_00909_, _11613_, p3_in[2]);
  and (_00910_, _00909_, _00908_);
  or (_00911_, _00910_, _00734_);
  nand (_00912_, _00734_, _08787_);
  and (_00913_, _00912_, _00911_);
  and (_00914_, _00913_, _08973_);
  or (_00915_, _00914_, _00907_);
  and (_00916_, _00915_, _00711_);
  or (_00917_, _11609_, p3in_reg[3]);
  or (_00918_, _11613_, p3_in[3]);
  and (_00919_, _00918_, _00917_);
  or (_00920_, _00919_, _00734_);
  or (_00921_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00922_, _00921_, _00920_);
  and (_00923_, _00922_, _00700_);
  or (_00924_, _00923_, _00916_);
  or (_00925_, _11609_, p3in_reg[4]);
  or (_00926_, _11613_, p3_in[4]);
  and (_00927_, _00926_, _00925_);
  or (_00928_, _00927_, _00734_);
  or (_00929_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_00930_, _00929_, _00928_);
  or (_00931_, _00930_, _08973_);
  or (_00932_, _11609_, p3in_reg[0]);
  or (_00933_, _11613_, p3_in[0]);
  and (_00934_, _00933_, _00932_);
  or (_00935_, _00934_, _00734_);
  or (_00936_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_00937_, _00936_, _00935_);
  or (_00938_, _00937_, _00667_);
  and (_00939_, _00938_, _00693_);
  and (_00940_, _00939_, _00931_);
  or (_00941_, _11609_, p3in_reg[5]);
  or (_00942_, _11613_, p3_in[5]);
  and (_00943_, _00942_, _00941_);
  or (_00944_, _00943_, _00734_);
  or (_00945_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00946_, _00945_, _00944_);
  and (_00947_, _00946_, _00667_);
  or (_00948_, _11609_, p3in_reg[1]);
  or (_00949_, _11613_, p3_in[1]);
  and (_00950_, _00949_, _00948_);
  or (_00951_, _00950_, _00734_);
  or (_00952_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_00953_, _00952_, _00951_);
  and (_00954_, _00953_, _08973_);
  or (_00955_, _00954_, _00947_);
  and (_00956_, _00955_, _00704_);
  or (_00957_, _11609_, p3in_reg[7]);
  or (_00958_, _11613_, p3_in[7]);
  and (_00959_, _00958_, _00957_);
  or (_00960_, _00959_, _00734_);
  nand (_00961_, _00734_, _08481_);
  and (_00962_, _00961_, _00960_);
  and (_00963_, _00962_, _00698_);
  or (_00964_, _00963_, _00956_);
  or (_00965_, _00964_, _00940_);
  or (_00966_, _00965_, _00924_);
  and (_00967_, _00809_, _00805_);
  and (_00968_, _00967_, _00966_);
  and (_00969_, _00693_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00970_, _00969_, _08973_);
  and (_00971_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00972_, _00711_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_00973_, _00704_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00974_, _00973_, _00972_);
  or (_00975_, _00974_, _00971_);
  or (_00976_, _00975_, _00970_);
  and (_00977_, _00808_, _00803_);
  and (_00978_, _00693_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00979_, _00978_, _00667_);
  and (_00980_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00981_, _00711_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_00982_, _00704_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00983_, _00982_, _00981_);
  or (_00984_, _00983_, _00980_);
  or (_00985_, _00984_, _00979_);
  and (_00986_, _00985_, _00977_);
  and (_00987_, _00986_, _00976_);
  or (_00988_, _00987_, _00968_);
  or (_00989_, _11609_, p0in_reg[4]);
  or (_00990_, _11613_, p0_in[4]);
  and (_00991_, _00990_, _00989_);
  or (_00992_, _00991_, _00734_);
  or (_00993_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_00994_, _00993_, _00992_);
  or (_00995_, _00994_, _08973_);
  or (_00996_, _11609_, p0in_reg[0]);
  or (_00997_, _11613_, p0_in[0]);
  and (_00998_, _00997_, _00996_);
  or (_00999_, _00998_, _00734_);
  or (_01000_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00667_);
  and (_01003_, _01002_, _00693_);
  and (_01004_, _01003_, _00995_);
  or (_01005_, _11609_, p0in_reg[3]);
  or (_01006_, _11613_, p0_in[3]);
  and (_01007_, _01006_, _01005_);
  or (_01008_, _01007_, _00734_);
  or (_01009_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_01010_, _01009_, _01008_);
  and (_01011_, _01010_, _00700_);
  or (_01012_, _01011_, _01004_);
  or (_01013_, _11609_, p0in_reg[6]);
  or (_01014_, _11613_, p0_in[6]);
  and (_01015_, _01014_, _01013_);
  or (_01017_, _01015_, _00734_);
  nand (_01018_, _00734_, _08577_);
  and (_01019_, _01018_, _01017_);
  and (_01020_, _01019_, _00667_);
  or (_01021_, _11609_, p0in_reg[2]);
  or (_01022_, _11613_, p0_in[2]);
  and (_01023_, _01022_, _01021_);
  or (_01024_, _01023_, _00734_);
  nand (_01025_, _00734_, _08533_);
  and (_01026_, _01025_, _01024_);
  and (_01027_, _01026_, _08973_);
  or (_01028_, _01027_, _01020_);
  and (_01029_, _01028_, _00711_);
  or (_01030_, _11609_, p0in_reg[5]);
  or (_01031_, _11613_, p0_in[5]);
  and (_01032_, _01031_, _01030_);
  or (_01033_, _01032_, _00734_);
  or (_01034_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01035_, _01034_, _01033_);
  and (_01036_, _01035_, _00667_);
  or (_01037_, _11609_, p0in_reg[1]);
  or (_01038_, _11613_, p0_in[1]);
  and (_01039_, _01038_, _01037_);
  or (_01040_, _01039_, _00734_);
  or (_01041_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01042_, _01041_, _01040_);
  and (_01043_, _01042_, _08973_);
  or (_01044_, _01043_, _01036_);
  and (_01045_, _01044_, _00704_);
  or (_01046_, _01045_, _01029_);
  or (_01048_, _11609_, p0in_reg[7]);
  or (_01049_, _11613_, p0_in[7]);
  and (_01050_, _01049_, _01048_);
  or (_01051_, _01050_, _00734_);
  nand (_01052_, _00734_, _08443_);
  and (_01053_, _01052_, _01051_);
  and (_01054_, _01053_, _00698_);
  or (_01055_, _01054_, _01046_);
  or (_01056_, _01055_, _01012_);
  and (_01057_, _09354_, _09023_);
  and (_01058_, _01057_, _00896_);
  and (_01059_, _01058_, _09194_);
  and (_01060_, _01059_, _01056_);
  and (_01061_, _00896_, _09194_);
  or (_01062_, _00810_, _00666_);
  or (_01063_, _01062_, _01061_);
  or (_01064_, _01063_, _00977_);
  and (_01065_, _01064_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_01066_, _01065_, _11651_);
  or (_01067_, _01066_, _01060_);
  or (_01069_, _01067_, _00988_);
  or (_01070_, _01069_, _00900_);
  or (_01071_, _01070_, _00717_);
  and (_01072_, _00977_, _08315_);
  and (_01073_, _01066_, _06829_);
  nor (_01074_, _01073_, _01072_);
  and (_01075_, _01074_, _01071_);
  not (_01076_, _08214_);
  and (_01077_, _01061_, _00739_);
  nor (_01078_, _01077_, _01076_);
  and (_01079_, _01078_, _01064_);
  nand (_01080_, _01079_, _11655_);
  nand (_01081_, _00697_, _08342_);
  nand (_01082_, _00704_, _08419_);
  and (_01083_, _01082_, _00667_);
  nand (_01084_, _00693_, _08406_);
  nand (_01085_, _00711_, _08431_);
  and (_01086_, _01085_, _01084_);
  and (_01087_, _01086_, _01083_);
  and (_01088_, _01087_, _01081_);
  and (_01089_, _00693_, _08353_);
  and (_01090_, _00704_, _08365_);
  or (_01091_, _01090_, _00667_);
  and (_01092_, _00711_, _08377_);
  and (_01093_, _00697_, _08394_);
  or (_01094_, _01093_, _01092_);
  or (_01095_, _01094_, _01091_);
  or (_01096_, _01095_, _01089_);
  nand (_01097_, _01096_, _01072_);
  or (_01098_, _01097_, _01088_);
  nand (_01099_, _01098_, _01080_);
  or (_01100_, _01099_, _01075_);
  not (_01101_, _07818_);
  and (_01102_, _00698_, _01101_);
  or (_01103_, _08973_, _09205_);
  nand (_01104_, _08973_, _07783_);
  and (_01105_, _01104_, _00711_);
  and (_01106_, _01105_, _01103_);
  nand (_01107_, _00667_, _07768_);
  nand (_01108_, _08973_, _07797_);
  and (_01109_, _01108_, _00693_);
  and (_01110_, _01109_, _01107_);
  or (_01111_, _01110_, _01106_);
  nand (_01112_, _00667_, _07761_);
  nand (_01113_, _08973_, _07790_);
  and (_01114_, _01113_, _00704_);
  and (_01115_, _01114_, _01112_);
  and (_01116_, _00700_, _09147_);
  or (_01117_, _01116_, _01115_);
  or (_01118_, _01117_, _01111_);
  or (_01119_, _01118_, _01102_);
  or (_01120_, _01119_, _01080_);
  and (_01121_, _01120_, _12493_);
  and (_12732_, _01121_, _01100_);
  and (_01122_, _09194_, _08973_);
  and (_01123_, _01122_, _00697_);
  and (_01124_, _01123_, _01058_);
  and (_01125_, _01124_, _07869_);
  not (_01126_, _01125_);
  and (_01127_, _01122_, _00693_);
  and (_01128_, _01127_, _00663_);
  and (_01129_, _01128_, _00664_);
  nand (_01130_, _01129_, _11714_);
  and (_01131_, _01130_, _01126_);
  nor (_01132_, _01131_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_01133_, _00698_, _08328_);
  and (_01134_, _01133_, _11655_);
  or (_01135_, _08325_, _08315_);
  and (_01136_, _09354_, _09024_);
  and (_01137_, _01136_, _01128_);
  and (_01138_, _01137_, _01135_);
  or (_01139_, _01138_, _01134_);
  or (_01140_, _01139_, _11653_);
  or (_01141_, _01140_, _01132_);
  and (_01142_, _01122_, _00711_);
  and (_01143_, _01142_, _01058_);
  and (_01144_, _01143_, _07869_);
  nor (_01145_, _01144_, rst);
  and (_12733_, _01145_, _01141_);
  not (_01146_, _01141_);
  or (_01147_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_01148_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_01149_, _01127_, _00896_);
  and (_01150_, _01149_, _01136_);
  and (_01151_, _01150_, _00765_);
  or (_01152_, _01151_, _01148_);
  nor (_01153_, _09354_, _09023_);
  and (_01154_, _01153_, _01128_);
  and (_01155_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_01156_, _01149_, _00664_);
  and (_01157_, _01156_, _00884_);
  or (_01158_, _01157_, _01155_);
  or (_01159_, _01158_, _01152_);
  and (_01160_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_01161_, _01122_, _00704_);
  and (_01162_, _01161_, _01058_);
  and (_01163_, _01162_, _07820_);
  or (_01164_, _01163_, _01160_);
  and (_01165_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_01166_, _01127_, _01058_);
  and (_01167_, _01166_, _01053_);
  or (_01168_, _01167_, _01165_);
  or (_01169_, _01168_, _01164_);
  and (_01170_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01171_, _01153_, _01149_);
  and (_01172_, _01171_, _00962_);
  or (_01173_, _01172_, _01170_);
  or (_01174_, _01173_, _01169_);
  or (_01175_, _01174_, _01159_);
  or (_01176_, _01175_, _01141_);
  and (_01177_, _01176_, _01147_);
  or (_01178_, _01177_, _01144_);
  nand (_01179_, _01144_, _06770_);
  and (_01180_, _01179_, _12493_);
  and (_12734_[7], _01180_, _01178_);
  and (_01181_, _01129_, _00691_);
  and (_01182_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01183_, _01150_, _00795_);
  and (_01184_, _01156_, _00858_);
  or (_01185_, _01184_, _01183_);
  or (_01186_, _01185_, _01182_);
  and (_01187_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_01188_, _01162_, _09122_);
  or (_01189_, _01188_, _01187_);
  and (_01190_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01191_, _01166_, _01001_);
  or (_01192_, _01191_, _01190_);
  or (_01193_, _01192_, _01189_);
  and (_01194_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_01195_, _01171_, _00937_);
  or (_01196_, _01195_, _01194_);
  or (_01197_, _01196_, _01193_);
  or (_01198_, _01197_, _01186_);
  or (_01199_, _01198_, _01141_);
  or (_01200_, _01199_, _01181_);
  or (_01201_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_01202_, _01201_, _01200_);
  or (_01203_, _01202_, _01144_);
  nand (_01204_, _01144_, _06877_);
  and (_01205_, _01204_, _12493_);
  and (_12734_[0], _01205_, _01203_);
  or (_01206_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_01207_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_01208_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_01209_, _01208_, _01207_);
  and (_01210_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01211_, _01156_, _00842_);
  or (_01212_, _01211_, _01210_);
  or (_01213_, _01212_, _01209_);
  and (_01214_, _01150_, _00779_);
  and (_01215_, _01171_, _00953_);
  or (_01216_, _01215_, _01214_);
  and (_01217_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_01218_, _01162_, _09298_);
  or (_01219_, _01218_, _01217_);
  and (_01220_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_01221_, _01166_, _01042_);
  or (_01222_, _01221_, _01220_);
  or (_01223_, _01222_, _01219_);
  or (_01224_, _01223_, _01216_);
  or (_01225_, _01224_, _01213_);
  or (_01226_, _01225_, _01141_);
  and (_01227_, _01226_, _01206_);
  or (_01228_, _01227_, _01144_);
  nand (_01229_, _01144_, _06939_);
  and (_01230_, _01229_, _12493_);
  and (_12734_[1], _01230_, _01228_);
  or (_01231_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_01232_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01233_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_01234_, _01233_, _01232_);
  and (_01235_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01236_, _01156_, _00875_);
  or (_01237_, _01236_, _01235_);
  or (_01238_, _01237_, _01234_);
  and (_01239_, _01150_, _00748_);
  and (_01240_, _01171_, _00913_);
  or (_01241_, _01240_, _01239_);
  and (_01242_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_01243_, _01166_, _01026_);
  or (_01244_, _01243_, _01242_);
  and (_01245_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_01246_, _01162_, _08943_);
  or (_01247_, _01246_, _01245_);
  or (_01248_, _01247_, _01244_);
  or (_01249_, _01248_, _01241_);
  or (_01250_, _01249_, _01238_);
  or (_01251_, _01250_, _01141_);
  and (_01252_, _01251_, _01231_);
  or (_01253_, _01252_, _01144_);
  nand (_01254_, _01144_, _07000_);
  and (_01255_, _01254_, _12493_);
  and (_12734_[2], _01255_, _01253_);
  or (_01256_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_01257_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01258_, _01156_, _00891_);
  or (_01259_, _01258_, _01257_);
  and (_01260_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01261_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_01262_, _01261_, _01260_);
  or (_01263_, _01262_, _01259_);
  and (_01264_, _01150_, _00757_);
  and (_01265_, _01171_, _00922_);
  or (_01266_, _01265_, _01264_);
  and (_01267_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_01268_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_01269_, _01268_, _01267_);
  and (_01270_, _01162_, _09170_);
  and (_01271_, _01166_, _01010_);
  or (_01272_, _01271_, _01270_);
  or (_01273_, _01272_, _01269_);
  or (_01274_, _01273_, _01266_);
  or (_01275_, _01274_, _01263_);
  or (_01276_, _01275_, _01141_);
  and (_01277_, _01276_, _01256_);
  or (_01278_, _01277_, _01144_);
  nand (_01279_, _01144_, _08058_);
  and (_01280_, _01279_, _12493_);
  and (_12734_[3], _01280_, _01278_);
  or (_01281_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_01282_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01283_, _01156_, _00851_);
  or (_01284_, _01283_, _01282_);
  and (_01285_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01286_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_01287_, _01286_, _01285_);
  or (_01288_, _01287_, _01284_);
  and (_01289_, _01150_, _00788_);
  and (_01290_, _01171_, _00930_);
  or (_01291_, _01290_, _01289_);
  and (_01292_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_01293_, _01166_, _00994_);
  or (_01294_, _01293_, _01292_);
  and (_01295_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  not (_01296_, _07852_);
  and (_01297_, _01162_, _01296_);
  or (_01298_, _01297_, _01295_);
  or (_01299_, _01298_, _01294_);
  or (_01300_, _01299_, _01291_);
  or (_01301_, _01300_, _01288_);
  or (_01302_, _01301_, _01141_);
  and (_01303_, _01302_, _01281_);
  or (_01304_, _01303_, _01144_);
  nand (_01305_, _01144_, _07134_);
  and (_01306_, _01305_, _12493_);
  and (_12734_[4], _01306_, _01304_);
  or (_01307_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_01308_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_01309_, _01156_, _00835_);
  or (_01310_, _01309_, _01308_);
  and (_01311_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01312_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_01313_, _01312_, _01311_);
  or (_01314_, _01313_, _01310_);
  and (_01315_, _01150_, _00772_);
  and (_01316_, _01171_, _00946_);
  or (_01317_, _01316_, _01315_);
  and (_01318_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01319_, _01166_, _01035_);
  or (_01320_, _01319_, _01318_);
  and (_01321_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  not (_01322_, _07858_);
  and (_01323_, _01162_, _01322_);
  or (_01324_, _01323_, _01321_);
  or (_01325_, _01324_, _01320_);
  or (_01326_, _01325_, _01317_);
  or (_01327_, _01326_, _01314_);
  or (_01328_, _01327_, _01141_);
  and (_01329_, _01328_, _01307_);
  or (_01330_, _01329_, _01144_);
  nand (_01331_, _01144_, _08120_);
  and (_01332_, _01331_, _12493_);
  and (_12734_[5], _01332_, _01330_);
  or (_01333_, _01146_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_01334_, _01154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01335_, _01137_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_01336_, _01335_, _01334_);
  and (_01337_, _01129_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01338_, _01156_, _00868_);
  or (_01339_, _01338_, _01337_);
  or (_01340_, _01339_, _01336_);
  and (_01341_, _01150_, _00741_);
  and (_01342_, _01171_, _00906_);
  or (_01343_, _01342_, _01341_);
  and (_01344_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01345_, _01124_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01346_, _01345_, _01344_);
  not (_01347_, _07864_);
  and (_01348_, _01162_, _01347_);
  and (_01349_, _01166_, _01019_);
  or (_01350_, _01349_, _01348_);
  or (_01351_, _01350_, _01346_);
  or (_01352_, _01351_, _01343_);
  or (_01353_, _01352_, _01340_);
  or (_01354_, _01353_, _01141_);
  and (_01355_, _01354_, _01333_);
  or (_01356_, _01355_, _01144_);
  nand (_01357_, _01144_, _07285_);
  and (_01358_, _01357_, _12493_);
  and (_12734_[6], _01358_, _01356_);
  and (_12728_, _09367_, _12493_);
  and (_12729_[7], _09056_, _12493_);
  nor (_12731_[2], _08973_, rst);
  and (_12729_[0], _09106_, _12493_);
  and (_12729_[1], _09266_, _12493_);
  and (_12729_[2], _08923_, _12493_);
  and (_12729_[3], _09155_, _12493_);
  and (_12729_[4], _09314_, _12493_);
  and (_12729_[5], _08983_, _12493_);
  and (_12729_[6], _09214_, _12493_);
  nor (_12731_[0], _09145_, rst);
  nor (_12731_[1], _09304_, rst);
  nor (_01359_, _12455_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01360_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _12143_);
  nor (_01361_, _01360_, _01359_);
  not (_01362_, _01361_);
  nor (_01363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01364_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _12143_);
  nor (_01365_, _01364_, _01363_);
  nor (_01366_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _12143_);
  nor (_01368_, _01367_, _01366_);
  nor (_01369_, _01368_, _01365_);
  not (_01370_, _01369_);
  nor (_01371_, _12438_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01372_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _12143_);
  nor (_01373_, _01372_, _01371_);
  and (_01374_, _01373_, _01370_);
  nor (_01375_, _01373_, _01370_);
  nor (_01376_, _01375_, _01374_);
  and (_01377_, _01376_, _01362_);
  and (_01378_, _01368_, _01365_);
  and (_01379_, _01378_, _01377_);
  and (_01380_, _01379_, _10416_);
  not (_01381_, _01365_);
  nor (_01382_, _01368_, _01381_);
  or (_01383_, _01361_, _01375_);
  or (_01384_, _01362_, _01374_);
  and (_01385_, _01384_, _01383_);
  and (_01386_, _01385_, _01382_);
  and (_01387_, _01386_, _10161_);
  or (_01388_, _01387_, _01380_);
  and (_01389_, _01382_, _01377_);
  and (_01390_, _01389_, _10325_);
  and (_01391_, _01376_, _01361_);
  and (_01392_, _01391_, _01382_);
  and (_01393_, _01392_, _10756_);
  or (_01394_, _01393_, _01390_);
  or (_01395_, _01394_, _01388_);
  and (_01396_, _01368_, _01381_);
  and (_01397_, _01396_, _01377_);
  and (_01398_, _01397_, _10366_);
  and (_01399_, _01385_, _01378_);
  and (_01400_, _01399_, _10243_);
  or (_01401_, _01400_, _01398_);
  and (_01402_, _01396_, _01385_);
  and (_01403_, _01402_, _10202_);
  and (_01404_, _01391_, _01378_);
  and (_01405_, _01404_, _10862_);
  or (_01406_, _01405_, _01403_);
  or (_01407_, _01406_, _01401_);
  and (_01408_, _01362_, _01373_);
  and (_01409_, _01408_, _01382_);
  and (_01410_, _01409_, _10528_);
  and (_01411_, _01408_, _01378_);
  and (_01412_, _01411_, _10642_);
  and (_01413_, _01408_, _01396_);
  and (_01414_, _01413_, _10586_);
  or (_01415_, _01414_, _01412_);
  or (_01416_, _01415_, _01410_);
  and (_01417_, _01396_, _01391_);
  and (_01418_, _01417_, _10814_);
  and (_01419_, _01373_, _01369_);
  and (_01420_, _01419_, _01361_);
  and (_01421_, _01420_, _10903_);
  and (_01422_, _01361_, _01375_);
  and (_01423_, _01422_, _10699_);
  or (_01424_, _01423_, _01421_);
  and (_01425_, _01362_, _01375_);
  and (_01426_, _01425_, _10284_);
  and (_01427_, _01419_, _01362_);
  and (_01428_, _01427_, _10472_);
  or (_01429_, _01428_, _01426_);
  or (_01430_, _01429_, _01424_);
  or (_01431_, _01430_, _01418_);
  or (_01432_, _01431_, _01416_);
  or (_01433_, _01432_, _01407_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01433_, _01395_);
  and (_01434_, _01379_, _10325_);
  and (_01435_, _01389_, _10243_);
  or (_01436_, _01435_, _01434_);
  and (_01437_, _01402_, _10903_);
  and (_01438_, _01399_, _10161_);
  or (_01439_, _01438_, _01437_);
  or (_01440_, _01439_, _01436_);
  and (_01441_, _01392_, _10642_);
  and (_01442_, _01417_, _10699_);
  or (_01443_, _01442_, _01441_);
  and (_01444_, _01397_, _10284_);
  and (_01445_, _01404_, _10756_);
  or (_01446_, _01445_, _01444_);
  or (_01447_, _01446_, _01443_);
  and (_01448_, _01413_, _10472_);
  and (_01449_, _01409_, _10416_);
  and (_01450_, _01411_, _10528_);
  or (_01451_, _01450_, _01449_);
  or (_01452_, _01451_, _01448_);
  and (_01453_, _01386_, _10862_);
  and (_01454_, _01422_, _10586_);
  and (_01455_, _01420_, _10814_);
  or (_01456_, _01455_, _01454_);
  and (_01457_, _01427_, _10366_);
  and (_01458_, _01425_, _10202_);
  or (_01459_, _01458_, _01457_);
  or (_01460_, _01459_, _01456_);
  or (_01461_, _01460_, _01453_);
  or (_01462_, _01461_, _01452_);
  or (_01463_, _01462_, _01447_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01463_, _01440_);
  and (_01464_, _01404_, _10814_);
  and (_01465_, _01402_, _10161_);
  or (_01466_, _01465_, _01464_);
  and (_01467_, _01399_, _10202_);
  and (_01468_, _01379_, _10366_);
  or (_01469_, _01468_, _01467_);
  or (_01470_, _01469_, _01466_);
  and (_01471_, _01386_, _10903_);
  and (_01472_, _01417_, _10756_);
  or (_01473_, _01472_, _01471_);
  and (_01474_, _01392_, _10699_);
  and (_01475_, _01397_, _10325_);
  or (_01476_, _01475_, _01474_);
  or (_01477_, _01476_, _01473_);
  and (_01478_, _01409_, _10472_);
  and (_01479_, _01411_, _10586_);
  and (_01480_, _01413_, _10528_);
  or (_01481_, _01480_, _01479_);
  or (_01482_, _01481_, _01478_);
  and (_01483_, _01389_, _10284_);
  and (_01484_, _01420_, _10862_);
  and (_01485_, _01422_, _10642_);
  or (_01486_, _01485_, _01484_);
  and (_01487_, _01425_, _10243_);
  and (_01488_, _01427_, _10416_);
  or (_01489_, _01488_, _01487_);
  or (_01490_, _01489_, _01486_);
  or (_01491_, _01490_, _01483_);
  or (_01492_, _01491_, _01482_);
  or (_01493_, _01492_, _01477_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01493_, _01470_);
  and (_01494_, _01392_, _10586_);
  and (_01495_, _01386_, _10814_);
  or (_01496_, _01495_, _01494_);
  and (_01497_, _01397_, _10243_);
  and (_01498_, _01404_, _10699_);
  or (_01499_, _01498_, _01497_);
  or (_01500_, _01499_, _01496_);
  and (_01501_, _01399_, _10903_);
  and (_01502_, _01417_, _10642_);
  or (_01503_, _01502_, _01501_);
  and (_01504_, _01389_, _10202_);
  and (_01505_, _01379_, _10284_);
  or (_01506_, _01505_, _01504_);
  or (_01507_, _01506_, _01503_);
  and (_01508_, _01409_, _10366_);
  and (_01509_, _01413_, _10416_);
  and (_01510_, _01411_, _10472_);
  or (_01511_, _01510_, _01509_);
  or (_01512_, _01511_, _01508_);
  and (_01513_, _01402_, _10862_);
  and (_01514_, _01427_, _10325_);
  and (_01515_, _01420_, _10756_);
  or (_01516_, _01515_, _01514_);
  and (_01517_, _01425_, _10161_);
  and (_01518_, _01422_, _10528_);
  or (_01519_, _01518_, _01517_);
  or (_01520_, _01519_, _01516_);
  or (_01521_, _01520_, _01513_);
  or (_01522_, _01521_, _01512_);
  or (_01523_, _01522_, _01507_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01523_, _01500_);
  and (_01524_, _01397_, _10371_);
  and (_01525_, _01399_, _10248_);
  or (_01526_, _01525_, _01524_);
  and (_01527_, _01402_, _10207_);
  and (_01528_, _01404_, _10867_);
  or (_01529_, _01528_, _01527_);
  or (_01530_, _01529_, _01526_);
  and (_01531_, _01379_, _10423_);
  and (_01532_, _01389_, _10330_);
  or (_01533_, _01532_, _01531_);
  and (_01534_, _01386_, _10166_);
  and (_01535_, _01392_, _10763_);
  or (_01536_, _01535_, _01534_);
  or (_01537_, _01536_, _01533_);
  and (_01538_, _01411_, _10649_);
  and (_01539_, _01413_, _10592_);
  or (_01540_, _01539_, _01538_);
  and (_01541_, _01409_, _10535_);
  or (_01542_, _01541_, _01540_);
  and (_01543_, _01417_, _10820_);
  and (_01544_, _01420_, _10908_);
  and (_01545_, _01425_, _10289_);
  or (_01546_, _01545_, _01544_);
  and (_01547_, _01427_, _10479_);
  and (_01548_, _01422_, _10706_);
  or (_01549_, _01548_, _01547_);
  or (_01550_, _01549_, _01546_);
  or (_01551_, _01550_, _01543_);
  or (_01552_, _01551_, _01542_);
  or (_01553_, _01552_, _01537_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01553_, _01530_);
  and (_01554_, _01404_, _10872_);
  and (_01555_, _01397_, _10377_);
  or (_01556_, _01555_, _01554_);
  and (_01557_, _01392_, _10770_);
  and (_01558_, _01402_, _10212_);
  or (_01559_, _01558_, _01557_);
  or (_01560_, _01559_, _01556_);
  and (_01561_, _01386_, _10171_);
  and (_01562_, _01389_, _10335_);
  or (_01563_, _01562_, _01561_);
  and (_01564_, _01417_, _10827_);
  and (_01565_, _01379_, _10430_);
  or (_01566_, _01565_, _01564_);
  or (_01567_, _01566_, _01563_);
  and (_01568_, _01409_, _10542_);
  and (_01569_, _01413_, _10599_);
  and (_01570_, _01411_, _10656_);
  or (_01571_, _01570_, _01569_);
  or (_01572_, _01571_, _01568_);
  and (_01573_, _01399_, _10253_);
  and (_01574_, _01420_, _10913_);
  and (_01575_, _01422_, _10713_);
  or (_01576_, _01575_, _01574_);
  and (_01577_, _01427_, _10486_);
  and (_01578_, _01425_, _10294_);
  or (_01579_, _01578_, _01577_);
  or (_01580_, _01579_, _01576_);
  or (_01581_, _01580_, _01573_);
  or (_01582_, _01581_, _01572_);
  or (_01583_, _01582_, _01567_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01583_, _01560_);
  and (_01584_, _01402_, _10217_);
  and (_01585_, _01404_, _10877_);
  or (_01586_, _01585_, _01584_);
  and (_01587_, _01397_, _10383_);
  and (_01588_, _01386_, _10176_);
  or (_01589_, _01588_, _01587_);
  or (_01590_, _01589_, _01586_);
  and (_01591_, _01399_, _10258_);
  and (_01592_, _01417_, _10834_);
  or (_01593_, _01592_, _01591_);
  and (_01594_, _01389_, _10340_);
  and (_01595_, _01392_, _10777_);
  or (_01596_, _01595_, _01594_);
  or (_01597_, _01596_, _01593_);
  and (_01598_, _01409_, _10549_);
  and (_01599_, _01413_, _10606_);
  and (_01600_, _01411_, _10663_);
  or (_01601_, _01600_, _01599_);
  or (_01602_, _01601_, _01598_);
  and (_01603_, _01379_, _10437_);
  and (_01604_, _01420_, _10918_);
  and (_01605_, _01425_, _10299_);
  or (_01606_, _01605_, _01604_);
  and (_01607_, _01427_, _10493_);
  and (_01608_, _01422_, _10720_);
  or (_01609_, _01608_, _01607_);
  or (_01610_, _01609_, _01606_);
  or (_01611_, _01610_, _01603_);
  or (_01612_, _01611_, _01602_);
  or (_01613_, _01612_, _01597_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01613_, _01590_);
  and (_01614_, _01386_, _10181_);
  and (_01615_, _01379_, _10443_);
  or (_01616_, _01615_, _01614_);
  and (_01617_, _01392_, _10784_);
  and (_01618_, _01389_, _10345_);
  or (_01619_, _01618_, _01617_);
  or (_01620_, _01619_, _01616_);
  and (_01621_, _01417_, _10841_);
  and (_01622_, _01402_, _10222_);
  or (_01623_, _01622_, _01621_);
  and (_01624_, _01399_, _10263_);
  and (_01625_, _01397_, _10389_);
  or (_01626_, _01625_, _01624_);
  or (_01627_, _01626_, _01623_);
  and (_01628_, _01409_, _10556_);
  and (_01629_, _01411_, _10670_);
  and (_01630_, _01413_, _10614_);
  or (_01631_, _01630_, _01629_);
  or (_01632_, _01631_, _01628_);
  and (_01633_, _01404_, _10882_);
  and (_01634_, _01420_, _10923_);
  and (_01635_, _01422_, _10727_);
  or (_01636_, _01635_, _01634_);
  and (_01637_, _01427_, _10500_);
  and (_01638_, _01425_, _10304_);
  or (_01639_, _01638_, _01637_);
  or (_01640_, _01639_, _01636_);
  or (_01641_, _01640_, _01633_);
  or (_01642_, _01641_, _01632_);
  or (_01643_, _01642_, _01627_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01643_, _01620_);
  and (_01644_, _01417_, _10846_);
  and (_01645_, _01402_, _10227_);
  or (_01646_, _01645_, _01644_);
  and (_01647_, _01404_, _10887_);
  and (_01648_, _01397_, _10396_);
  or (_01649_, _01648_, _01647_);
  or (_01650_, _01649_, _01646_);
  and (_01651_, _01392_, _10791_);
  and (_01652_, _01399_, _10268_);
  or (_01653_, _01652_, _01651_);
  and (_01654_, _01386_, _10186_);
  and (_01655_, _01389_, _10350_);
  or (_01656_, _01655_, _01654_);
  or (_01657_, _01656_, _01653_);
  and (_01658_, _01409_, _10563_);
  and (_01659_, _01413_, _10619_);
  and (_01660_, _01411_, _10677_);
  or (_01661_, _01660_, _01659_);
  or (_01662_, _01661_, _01658_);
  and (_01663_, _01379_, _10450_);
  and (_01664_, _01420_, _10928_);
  and (_01665_, _01425_, _10309_);
  or (_01666_, _01665_, _01664_);
  and (_01667_, _01427_, _10506_);
  and (_01668_, _01422_, _10734_);
  or (_01669_, _01668_, _01667_);
  or (_01670_, _01669_, _01666_);
  or (_01671_, _01670_, _01663_);
  or (_01672_, _01671_, _01662_);
  or (_01673_, _01672_, _01657_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01673_, _01650_);
  and (_01674_, _01417_, _10851_);
  and (_01675_, _01386_, _10191_);
  or (_01676_, _01675_, _01674_);
  and (_01677_, _01389_, _10355_);
  and (_01678_, _01399_, _10273_);
  or (_01679_, _01678_, _01677_);
  or (_01680_, _01679_, _01676_);
  and (_01681_, _01392_, _10798_);
  and (_01682_, _01397_, _10402_);
  or (_01683_, _01682_, _01681_);
  and (_01684_, _01404_, _10892_);
  and (_01685_, _01402_, _10232_);
  or (_01686_, _01685_, _01684_);
  or (_01687_, _01686_, _01683_);
  and (_01688_, _01409_, _10570_);
  and (_01689_, _01411_, _10684_);
  and (_01690_, _01413_, _10626_);
  or (_01691_, _01690_, _01689_);
  or (_01692_, _01691_, _01688_);
  and (_01693_, _01379_, _10457_);
  and (_01694_, _01420_, _10933_);
  and (_01695_, _01422_, _10741_);
  or (_01696_, _01695_, _01694_);
  and (_01697_, _01427_, _10513_);
  and (_01698_, _01425_, _10314_);
  or (_01699_, _01698_, _01697_);
  or (_01700_, _01699_, _01696_);
  or (_01701_, _01700_, _01693_);
  or (_01702_, _01701_, _01692_);
  or (_01703_, _01702_, _01687_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01703_, _01680_);
  and (_01704_, _01404_, _10897_);
  and (_01705_, _01397_, _10409_);
  or (_01706_, _01705_, _01704_);
  and (_01707_, _01392_, _10805_);
  and (_01708_, _01402_, _10237_);
  or (_01709_, _01708_, _01707_);
  or (_01710_, _01709_, _01706_);
  and (_01711_, _01386_, _10196_);
  and (_01712_, _01389_, _10360_);
  or (_01713_, _01712_, _01711_);
  and (_01714_, _01417_, _10856_);
  and (_01715_, _01379_, _10464_);
  or (_01716_, _01715_, _01714_);
  or (_01717_, _01716_, _01713_);
  and (_01718_, _01409_, _10577_);
  and (_01719_, _01413_, _10633_);
  and (_01720_, _01411_, _10691_);
  or (_01721_, _01720_, _01719_);
  or (_01722_, _01721_, _01718_);
  and (_01723_, _01399_, _10278_);
  and (_01724_, _01420_, _10938_);
  and (_01725_, _01422_, _10748_);
  or (_01726_, _01725_, _01724_);
  and (_01727_, _01427_, _10520_);
  and (_01728_, _01425_, _10319_);
  or (_01729_, _01728_, _01727_);
  or (_01730_, _01729_, _01726_);
  or (_01731_, _01730_, _01723_);
  or (_01732_, _01731_, _01722_);
  or (_01733_, _01732_, _01717_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01733_, _01710_);
  and (_01734_, _01389_, _10248_);
  and (_01735_, _01379_, _10330_);
  or (_01736_, _01735_, _01734_);
  and (_01737_, _01402_, _10908_);
  and (_01738_, _01399_, _10166_);
  or (_01739_, _01738_, _01737_);
  or (_01740_, _01739_, _01736_);
  and (_01741_, _01392_, _10649_);
  and (_01742_, _01417_, _10706_);
  or (_01743_, _01742_, _01741_);
  and (_01744_, _01397_, _10289_);
  and (_01745_, _01404_, _10763_);
  or (_01746_, _01745_, _01744_);
  or (_01747_, _01746_, _01743_);
  and (_01748_, _01413_, _10479_);
  and (_01749_, _01409_, _10423_);
  and (_01750_, _01411_, _10535_);
  or (_01751_, _01750_, _01749_);
  or (_01752_, _01751_, _01748_);
  and (_01753_, _01386_, _10867_);
  and (_01754_, _01422_, _10592_);
  and (_01755_, _01420_, _10820_);
  or (_01756_, _01755_, _01754_);
  and (_01757_, _01425_, _10207_);
  and (_01758_, _01427_, _10371_);
  or (_01759_, _01758_, _01757_);
  or (_01760_, _01759_, _01756_);
  or (_01761_, _01760_, _01753_);
  or (_01762_, _01761_, _01752_);
  or (_01763_, _01762_, _01747_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01763_, _01740_);
  and (_01764_, _01379_, _10335_);
  and (_01765_, _01389_, _10253_);
  or (_01766_, _01765_, _01764_);
  and (_01767_, _01402_, _10913_);
  and (_01768_, _01399_, _10171_);
  or (_01769_, _01768_, _01767_);
  or (_01770_, _01769_, _01766_);
  and (_01771_, _01392_, _10656_);
  and (_01772_, _01417_, _10713_);
  or (_01773_, _01772_, _01771_);
  and (_01774_, _01397_, _10294_);
  and (_01775_, _01404_, _10770_);
  or (_01776_, _01775_, _01774_);
  or (_01777_, _01776_, _01773_);
  and (_01778_, _01413_, _10486_);
  and (_01779_, _01409_, _10430_);
  and (_01780_, _01411_, _10542_);
  or (_01781_, _01780_, _01779_);
  or (_01782_, _01781_, _01778_);
  and (_01783_, _01386_, _10872_);
  and (_01784_, _01422_, _10599_);
  and (_01785_, _01420_, _10827_);
  or (_01786_, _01785_, _01784_);
  and (_01787_, _01427_, _10377_);
  and (_01788_, _01425_, _10212_);
  or (_01789_, _01788_, _01787_);
  or (_01790_, _01789_, _01786_);
  or (_01791_, _01790_, _01783_);
  or (_01792_, _01791_, _01782_);
  or (_01793_, _01792_, _01777_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01793_, _01770_);
  and (_01794_, _01389_, _10258_);
  and (_01795_, _01404_, _10777_);
  or (_01796_, _01795_, _01794_);
  and (_01797_, _01399_, _10176_);
  and (_01798_, _01386_, _10877_);
  or (_01799_, _01798_, _01797_);
  or (_01800_, _01799_, _01796_);
  and (_01801_, _01379_, _10340_);
  and (_01802_, _01397_, _10299_);
  or (_01803_, _01802_, _01801_);
  and (_01804_, _01402_, _10918_);
  and (_01805_, _01417_, _10720_);
  or (_01806_, _01805_, _01804_);
  or (_01807_, _01806_, _01803_);
  and (_01808_, _01411_, _10549_);
  and (_01809_, _01409_, _10437_);
  and (_01810_, _01413_, _10493_);
  or (_01811_, _01810_, _01809_);
  or (_01812_, _01811_, _01808_);
  and (_01813_, _01392_, _10663_);
  and (_01814_, _01422_, _10606_);
  and (_01815_, _01420_, _10834_);
  or (_01816_, _01815_, _01814_);
  and (_01817_, _01427_, _10383_);
  and (_01818_, _01425_, _10217_);
  or (_01819_, _01818_, _01817_);
  or (_01820_, _01819_, _01816_);
  or (_01821_, _01820_, _01813_);
  or (_01822_, _01821_, _01812_);
  or (_01823_, _01822_, _01807_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01823_, _01800_);
  and (_01824_, _01397_, _10304_);
  and (_01825_, _01389_, _10263_);
  or (_01826_, _01825_, _01824_);
  and (_01827_, _01402_, _10923_);
  and (_01828_, _01379_, _10345_);
  or (_01829_, _01828_, _01827_);
  or (_01830_, _01829_, _01826_);
  and (_01831_, _01392_, _10670_);
  and (_01832_, _01417_, _10727_);
  or (_01833_, _01832_, _01831_);
  and (_01834_, _01399_, _10181_);
  and (_01835_, _01404_, _10784_);
  or (_01836_, _01835_, _01834_);
  or (_01837_, _01836_, _01833_);
  and (_01838_, _01413_, _10500_);
  and (_01839_, _01409_, _10443_);
  and (_01840_, _01411_, _10556_);
  or (_01841_, _01840_, _01839_);
  or (_01842_, _01841_, _01838_);
  and (_01843_, _01386_, _10882_);
  and (_01844_, _01422_, _10614_);
  and (_01845_, _01420_, _10841_);
  or (_01846_, _01845_, _01844_);
  and (_01847_, _01427_, _10389_);
  and (_01848_, _01425_, _10222_);
  or (_01849_, _01848_, _01847_);
  or (_01850_, _01849_, _01846_);
  or (_01851_, _01850_, _01843_);
  or (_01852_, _01851_, _01842_);
  or (_01853_, _01852_, _01837_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01853_, _01830_);
  and (_01854_, _01389_, _10268_);
  and (_01855_, _01379_, _10350_);
  or (_01856_, _01855_, _01854_);
  and (_01857_, _01402_, _10928_);
  and (_01858_, _01399_, _10186_);
  or (_01859_, _01858_, _01857_);
  or (_01860_, _01859_, _01856_);
  and (_01861_, _01392_, _10677_);
  and (_01862_, _01417_, _10734_);
  or (_01863_, _01862_, _01861_);
  and (_01864_, _01397_, _10309_);
  and (_01865_, _01404_, _10791_);
  or (_01866_, _01865_, _01864_);
  or (_01867_, _01866_, _01863_);
  and (_01868_, _01413_, _10506_);
  and (_01869_, _01409_, _10450_);
  and (_01870_, _01411_, _10563_);
  or (_01871_, _01870_, _01869_);
  or (_01872_, _01871_, _01868_);
  and (_01873_, _01386_, _10887_);
  and (_01874_, _01422_, _10619_);
  and (_01875_, _01420_, _10846_);
  or (_01876_, _01875_, _01874_);
  and (_01877_, _01425_, _10227_);
  and (_01878_, _01427_, _10396_);
  or (_01879_, _01878_, _01877_);
  or (_01880_, _01879_, _01876_);
  or (_01881_, _01880_, _01873_);
  or (_01882_, _01881_, _01872_);
  or (_01883_, _01882_, _01867_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01883_, _01860_);
  and (_01884_, _01402_, _10933_);
  and (_01885_, _01417_, _10741_);
  or (_01886_, _01885_, _01884_);
  and (_01887_, _01389_, _10273_);
  and (_01888_, _01386_, _10892_);
  or (_01889_, _01888_, _01887_);
  or (_01890_, _01889_, _01886_);
  and (_01891_, _01379_, _10355_);
  and (_01892_, _01397_, _10314_);
  or (_01893_, _01892_, _01891_);
  and (_01894_, _01392_, _10684_);
  and (_01895_, _01404_, _10798_);
  or (_01896_, _01895_, _01894_);
  or (_01897_, _01896_, _01893_);
  and (_01898_, _01413_, _10513_);
  and (_01899_, _01409_, _10457_);
  and (_01900_, _01411_, _10570_);
  or (_01901_, _01900_, _01899_);
  or (_01902_, _01901_, _01898_);
  and (_01903_, _01399_, _10191_);
  and (_01904_, _01425_, _10232_);
  and (_01905_, _01420_, _10851_);
  or (_01906_, _01905_, _01904_);
  and (_01907_, _01427_, _10402_);
  and (_01908_, _01422_, _10626_);
  or (_01909_, _01908_, _01907_);
  or (_01910_, _01909_, _01906_);
  or (_01911_, _01910_, _01903_);
  or (_01912_, _01911_, _01902_);
  or (_01913_, _01912_, _01897_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01913_, _01890_);
  and (_01914_, _01379_, _10360_);
  and (_01915_, _01389_, _10278_);
  or (_01916_, _01915_, _01914_);
  and (_01917_, _01402_, _10938_);
  and (_01918_, _01399_, _10196_);
  or (_01919_, _01918_, _01917_);
  or (_01920_, _01919_, _01916_);
  and (_01921_, _01392_, _10691_);
  and (_01922_, _01417_, _10748_);
  or (_01923_, _01922_, _01921_);
  and (_01924_, _01397_, _10319_);
  and (_01925_, _01404_, _10805_);
  or (_01926_, _01925_, _01924_);
  or (_01927_, _01926_, _01923_);
  and (_01928_, _01413_, _10520_);
  and (_01929_, _01409_, _10464_);
  and (_01930_, _01411_, _10577_);
  or (_01931_, _01930_, _01929_);
  or (_01932_, _01931_, _01928_);
  and (_01933_, _01386_, _10897_);
  and (_01934_, _01422_, _10633_);
  and (_01935_, _01420_, _10856_);
  or (_01936_, _01935_, _01934_);
  and (_01937_, _01427_, _10409_);
  and (_01938_, _01425_, _10237_);
  or (_01939_, _01938_, _01937_);
  or (_01940_, _01939_, _01936_);
  or (_01941_, _01940_, _01933_);
  or (_01942_, _01941_, _01932_);
  or (_01943_, _01942_, _01927_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01943_, _01920_);
  and (_01944_, _01392_, _10706_);
  and (_01945_, _01397_, _10330_);
  or (_01946_, _01945_, _01944_);
  and (_01947_, _01399_, _10207_);
  and (_01948_, _01379_, _10371_);
  or (_01949_, _01948_, _01947_);
  or (_01950_, _01949_, _01946_);
  and (_01951_, _01386_, _10908_);
  and (_01952_, _01417_, _10763_);
  or (_01953_, _01952_, _01951_);
  and (_01954_, _01404_, _10820_);
  and (_01955_, _01389_, _10289_);
  or (_01956_, _01955_, _01954_);
  or (_01957_, _01956_, _01953_);
  and (_01958_, _01413_, _10535_);
  and (_01959_, _01409_, _10479_);
  or (_01960_, _01959_, _01958_);
  and (_01961_, _01411_, _10592_);
  or (_01962_, _01961_, _01960_);
  and (_01963_, _01402_, _10166_);
  and (_01964_, _01420_, _10867_);
  and (_01965_, _01425_, _10248_);
  or (_01966_, _01965_, _01964_);
  and (_01967_, _01422_, _10649_);
  and (_01968_, _01427_, _10423_);
  or (_01969_, _01968_, _01967_);
  or (_01970_, _01969_, _01966_);
  or (_01971_, _01970_, _01963_);
  or (_01972_, _01971_, _01962_);
  or (_01973_, _01972_, _01957_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01973_, _01950_);
  and (_01974_, _01392_, _10713_);
  and (_01975_, _01389_, _10294_);
  or (_01976_, _01975_, _01974_);
  and (_01977_, _01397_, _10335_);
  and (_01978_, _01402_, _10171_);
  or (_01979_, _01978_, _01977_);
  or (_01980_, _01979_, _01976_);
  and (_01981_, _01386_, _10913_);
  and (_01982_, _01417_, _10770_);
  or (_01983_, _01982_, _01981_);
  and (_01984_, _01404_, _10827_);
  and (_01985_, _01399_, _10212_);
  or (_01986_, _01985_, _01984_);
  or (_01987_, _01986_, _01983_);
  and (_01988_, _01409_, _10486_);
  and (_01989_, _01411_, _10599_);
  and (_01990_, _01413_, _10542_);
  or (_01991_, _01990_, _01989_);
  or (_01992_, _01991_, _01988_);
  and (_01993_, _01379_, _10377_);
  and (_01994_, _01420_, _10872_);
  and (_01995_, _01427_, _10430_);
  or (_01996_, _01995_, _01994_);
  and (_01997_, _01422_, _10656_);
  and (_01998_, _01425_, _10253_);
  or (_01999_, _01998_, _01997_);
  or (_02000_, _01999_, _01996_);
  or (_02001_, _02000_, _01993_);
  or (_02002_, _02001_, _01992_);
  or (_02003_, _02002_, _01987_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _02003_, _01980_);
  and (_02004_, _01389_, _10299_);
  and (_02005_, _01417_, _10777_);
  or (_02006_, _02005_, _02004_);
  and (_02007_, _01386_, _10918_);
  and (_02008_, _01402_, _10176_);
  or (_02009_, _02008_, _02007_);
  or (_02010_, _02009_, _02006_);
  and (_02011_, _01379_, _10383_);
  and (_02012_, _01399_, _10217_);
  or (_02013_, _02012_, _02011_);
  and (_02014_, _01397_, _10340_);
  and (_02015_, _01392_, _10720_);
  or (_02016_, _02015_, _02014_);
  or (_02017_, _02016_, _02013_);
  and (_02018_, _01409_, _10493_);
  and (_02019_, _01411_, _10606_);
  and (_02020_, _01413_, _10549_);
  or (_02021_, _02020_, _02019_);
  or (_02022_, _02021_, _02018_);
  and (_02023_, _01404_, _10834_);
  and (_02024_, _01427_, _10437_);
  and (_02025_, _01420_, _10877_);
  or (_02026_, _02025_, _02024_);
  and (_02027_, _01425_, _10258_);
  and (_02028_, _01422_, _10663_);
  or (_02029_, _02028_, _02027_);
  or (_02030_, _02029_, _02026_);
  or (_02031_, _02030_, _02023_);
  or (_02032_, _02031_, _02022_);
  or (_02033_, _02032_, _02017_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _02033_, _02010_);
  and (_02034_, _01399_, _10222_);
  and (_02035_, _01397_, _10345_);
  or (_02036_, _02035_, _02034_);
  and (_02037_, _01417_, _10784_);
  and (_02038_, _01402_, _10181_);
  or (_02039_, _02038_, _02037_);
  or (_02040_, _02039_, _02036_);
  and (_02041_, _01404_, _10841_);
  and (_02042_, _01392_, _10727_);
  or (_02043_, _02042_, _02041_);
  and (_02044_, _01379_, _10389_);
  and (_02045_, _01389_, _10304_);
  or (_02046_, _02045_, _02044_);
  or (_02047_, _02046_, _02043_);
  and (_02048_, _01413_, _10556_);
  and (_02049_, _01409_, _10500_);
  or (_02050_, _02049_, _02048_);
  and (_02051_, _01411_, _10614_);
  or (_02052_, _02051_, _02050_);
  and (_02053_, _01386_, _10923_);
  and (_02054_, _01420_, _10882_);
  and (_02055_, _01422_, _10670_);
  or (_02056_, _02055_, _02054_);
  and (_02057_, _01425_, _10263_);
  and (_02058_, _01427_, _10443_);
  or (_02059_, _02058_, _02057_);
  or (_02060_, _02059_, _02056_);
  or (_02061_, _02060_, _02053_);
  or (_02062_, _02061_, _02052_);
  or (_02063_, _02062_, _02047_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _02063_, _02040_);
  and (_02064_, _01404_, _10846_);
  and (_02065_, _01417_, _10791_);
  or (_02066_, _02065_, _02064_);
  and (_02067_, _01386_, _10928_);
  and (_02068_, _01397_, _10350_);
  or (_02069_, _02068_, _02067_);
  or (_02070_, _02069_, _02066_);
  and (_02071_, _01389_, _10309_);
  and (_02072_, _01402_, _10186_);
  or (_02073_, _02072_, _02071_);
  and (_02074_, _01399_, _10227_);
  and (_02075_, _01392_, _10734_);
  or (_02076_, _02075_, _02074_);
  or (_02077_, _02076_, _02073_);
  and (_02078_, _01413_, _10563_);
  and (_02079_, _01409_, _10506_);
  or (_02080_, _02079_, _02078_);
  and (_02081_, _01411_, _10619_);
  or (_02082_, _02081_, _02080_);
  and (_02083_, _01379_, _10396_);
  and (_02084_, _01427_, _10450_);
  and (_02085_, _01420_, _10887_);
  or (_02086_, _02085_, _02084_);
  and (_02087_, _01425_, _10268_);
  and (_02088_, _01422_, _10677_);
  or (_02089_, _02088_, _02087_);
  or (_02090_, _02089_, _02086_);
  or (_02091_, _02090_, _02083_);
  or (_02092_, _02091_, _02082_);
  or (_02093_, _02092_, _02077_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _02093_, _02070_);
  and (_02094_, _01386_, _10933_);
  and (_02095_, _01404_, _10851_);
  or (_02096_, _02095_, _02094_);
  and (_02097_, _01399_, _10232_);
  and (_02098_, _01417_, _10798_);
  or (_02099_, _02098_, _02097_);
  or (_02100_, _02099_, _02096_);
  and (_02101_, _01397_, _10355_);
  and (_02102_, _01402_, _10191_);
  or (_02103_, _02102_, _02101_);
  and (_02104_, _01389_, _10314_);
  and (_02105_, _01392_, _10741_);
  or (_02106_, _02105_, _02104_);
  or (_02107_, _02106_, _02103_);
  and (_02108_, _01409_, _10513_);
  and (_02109_, _01413_, _10570_);
  or (_02110_, _02109_, _02108_);
  and (_02111_, _01411_, _10626_);
  or (_02112_, _02111_, _02110_);
  and (_02113_, _01379_, _10402_);
  and (_02114_, _01422_, _10684_);
  and (_02115_, _01420_, _10892_);
  or (_02116_, _02115_, _02114_);
  and (_02117_, _01427_, _10457_);
  and (_02118_, _01425_, _10273_);
  or (_02119_, _02118_, _02117_);
  or (_02120_, _02119_, _02116_);
  or (_02121_, _02120_, _02113_);
  or (_02122_, _02121_, _02112_);
  or (_02123_, _02122_, _02107_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _02123_, _02100_);
  and (_02124_, _01404_, _10856_);
  and (_02125_, _01417_, _10805_);
  or (_02126_, _02125_, _02124_);
  and (_02127_, _01386_, _10938_);
  and (_02128_, _01397_, _10360_);
  or (_02129_, _02128_, _02127_);
  or (_02130_, _02129_, _02126_);
  and (_02131_, _01389_, _10319_);
  and (_02132_, _01402_, _10196_);
  or (_02133_, _02132_, _02131_);
  and (_02134_, _01399_, _10237_);
  and (_02135_, _01392_, _10748_);
  or (_02136_, _02135_, _02134_);
  or (_02137_, _02136_, _02133_);
  and (_02138_, _01413_, _10577_);
  and (_02139_, _01409_, _10520_);
  or (_02140_, _02139_, _02138_);
  and (_02141_, _01411_, _10633_);
  or (_02142_, _02141_, _02140_);
  and (_02143_, _01379_, _10409_);
  and (_02144_, _01427_, _10464_);
  and (_02145_, _01420_, _10897_);
  or (_02146_, _02145_, _02144_);
  and (_02147_, _01425_, _10278_);
  and (_02148_, _01422_, _10691_);
  or (_02149_, _02148_, _02147_);
  or (_02150_, _02149_, _02146_);
  or (_02151_, _02150_, _02143_);
  or (_02152_, _02151_, _02142_);
  or (_02153_, _02152_, _02137_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _02153_, _02130_);
  and (_02154_, _01392_, _10592_);
  and (_02155_, _01386_, _10820_);
  or (_02156_, _02155_, _02154_);
  and (_02157_, _01379_, _10289_);
  and (_02158_, _01404_, _10706_);
  or (_02159_, _02158_, _02157_);
  or (_02160_, _02159_, _02156_);
  and (_02161_, _01397_, _10248_);
  and (_02162_, _01417_, _10649_);
  or (_02163_, _02162_, _02161_);
  and (_02164_, _01399_, _10908_);
  and (_02165_, _01389_, _10207_);
  or (_02166_, _02165_, _02164_);
  or (_02167_, _02166_, _02163_);
  and (_02168_, _01409_, _10371_);
  and (_02169_, _01413_, _10423_);
  and (_02170_, _01411_, _10479_);
  or (_02171_, _02170_, _02169_);
  or (_02172_, _02171_, _02168_);
  and (_02173_, _01402_, _10867_);
  and (_02174_, _01422_, _10535_);
  and (_02175_, _01420_, _10763_);
  or (_02176_, _02175_, _02174_);
  and (_02177_, _01427_, _10330_);
  and (_02178_, _01425_, _10166_);
  or (_02179_, _02178_, _02177_);
  or (_02180_, _02179_, _02176_);
  or (_02181_, _02180_, _02173_);
  or (_02182_, _02181_, _02172_);
  or (_02183_, _02182_, _02167_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02183_, _02160_);
  and (_02184_, _01389_, _10212_);
  and (_02185_, _01386_, _10827_);
  or (_02186_, _02185_, _02184_);
  and (_02187_, _01399_, _10913_);
  and (_02188_, _01379_, _10294_);
  or (_02189_, _02188_, _02187_);
  or (_02190_, _02189_, _02186_);
  and (_02191_, _01392_, _10599_);
  and (_02192_, _01417_, _10656_);
  or (_02193_, _02192_, _02191_);
  and (_02194_, _01397_, _10253_);
  and (_02195_, _01404_, _10713_);
  or (_02196_, _02195_, _02194_);
  or (_02197_, _02196_, _02193_);
  and (_02198_, _01413_, _10430_);
  and (_02199_, _01409_, _10377_);
  and (_02200_, _01411_, _10486_);
  or (_02201_, _02200_, _02199_);
  or (_02202_, _02201_, _02198_);
  and (_02203_, _01402_, _10872_);
  and (_02204_, _01422_, _10542_);
  and (_02205_, _01420_, _10770_);
  or (_02206_, _02205_, _02204_);
  and (_02207_, _01425_, _10171_);
  and (_02208_, _01427_, _10335_);
  or (_02209_, _02208_, _02207_);
  or (_02210_, _02209_, _02206_);
  or (_02211_, _02210_, _02203_);
  or (_02212_, _02211_, _02202_);
  or (_02213_, _02212_, _02197_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02213_, _02190_);
  and (_02214_, _01379_, _10299_);
  and (_02215_, _01404_, _10720_);
  or (_02216_, _02215_, _02214_);
  and (_02217_, _01417_, _10663_);
  and (_02218_, _01386_, _10834_);
  or (_02219_, _02218_, _02217_);
  or (_02220_, _02219_, _02216_);
  and (_02221_, _01399_, _10918_);
  and (_02222_, _01389_, _10217_);
  or (_02223_, _02222_, _02221_);
  and (_02224_, _01397_, _10258_);
  and (_02225_, _01392_, _10606_);
  or (_02226_, _02225_, _02224_);
  or (_02227_, _02226_, _02223_);
  and (_02228_, _01413_, _10437_);
  and (_02229_, _01409_, _10383_);
  or (_02230_, _02229_, _02228_);
  and (_02231_, _01411_, _10493_);
  or (_02232_, _02231_, _02230_);
  and (_02233_, _01402_, _10877_);
  and (_02234_, _01427_, _10340_);
  and (_02235_, _01422_, _10549_);
  or (_02236_, _02235_, _02234_);
  and (_02237_, _01425_, _10176_);
  and (_02238_, _01420_, _10777_);
  or (_02239_, _02238_, _02237_);
  or (_02240_, _02239_, _02236_);
  or (_02241_, _02240_, _02233_);
  or (_02242_, _02241_, _02232_);
  or (_02243_, _02242_, _02227_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02243_, _02220_);
  and (_02244_, _01392_, _10614_);
  and (_02245_, _01386_, _10841_);
  or (_02246_, _02245_, _02244_);
  and (_02247_, _01397_, _10263_);
  and (_02248_, _01404_, _10727_);
  or (_02249_, _02248_, _02247_);
  or (_02250_, _02249_, _02246_);
  and (_02251_, _01379_, _10304_);
  and (_02252_, _01417_, _10670_);
  or (_02253_, _02252_, _02251_);
  and (_02254_, _01399_, _10923_);
  and (_02255_, _01389_, _10222_);
  or (_02256_, _02255_, _02254_);
  or (_02257_, _02256_, _02253_);
  and (_02258_, _01413_, _10443_);
  and (_02259_, _01409_, _10389_);
  and (_02260_, _01411_, _10500_);
  or (_02261_, _02260_, _02259_);
  or (_02262_, _02261_, _02258_);
  and (_02263_, _01402_, _10882_);
  and (_02264_, _01422_, _10556_);
  and (_02265_, _01420_, _10784_);
  or (_02266_, _02265_, _02264_);
  and (_02267_, _01427_, _10345_);
  and (_02268_, _01425_, _10181_);
  or (_02269_, _02268_, _02267_);
  or (_02270_, _02269_, _02266_);
  or (_02271_, _02270_, _02263_);
  or (_02272_, _02271_, _02262_);
  or (_02273_, _02272_, _02257_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02273_, _02250_);
  and (_02274_, _01379_, _10309_);
  and (_02275_, _01386_, _10846_);
  or (_02276_, _02275_, _02274_);
  and (_02277_, _01399_, _10928_);
  and (_02278_, _01397_, _10268_);
  or (_02279_, _02278_, _02277_);
  or (_02280_, _02279_, _02276_);
  and (_02281_, _01417_, _10677_);
  and (_02282_, _01404_, _10734_);
  or (_02283_, _02282_, _02281_);
  and (_02284_, _01389_, _10227_);
  and (_02285_, _01392_, _10619_);
  or (_02286_, _02285_, _02284_);
  or (_02287_, _02286_, _02283_);
  and (_02288_, _01409_, _10396_);
  and (_02289_, _01413_, _10450_);
  and (_02290_, _01411_, _10506_);
  or (_02291_, _02290_, _02289_);
  or (_02292_, _02291_, _02288_);
  and (_02293_, _01402_, _10887_);
  and (_02294_, _01422_, _10563_);
  and (_02295_, _01420_, _10791_);
  or (_02296_, _02295_, _02294_);
  and (_02297_, _01427_, _10350_);
  and (_02298_, _01425_, _10186_);
  or (_02299_, _02298_, _02297_);
  or (_02300_, _02299_, _02296_);
  or (_02301_, _02300_, _02293_);
  or (_02302_, _02301_, _02292_);
  or (_02303_, _02302_, _02287_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02303_, _02280_);
  and (_02304_, _01417_, _10684_);
  and (_02305_, _01402_, _10892_);
  or (_02306_, _02305_, _02304_);
  and (_02307_, _01397_, _10273_);
  and (_02308_, _01404_, _10741_);
  or (_02309_, _02308_, _02307_);
  or (_02310_, _02309_, _02306_);
  and (_02311_, _01379_, _10314_);
  and (_02312_, _01386_, _10851_);
  or (_02313_, _02312_, _02311_);
  and (_02314_, _01399_, _10933_);
  and (_02315_, _01392_, _10626_);
  or (_02316_, _02315_, _02314_);
  or (_02317_, _02316_, _02313_);
  and (_02318_, _01413_, _10457_);
  and (_02319_, _01409_, _10402_);
  or (_02320_, _02319_, _02318_);
  and (_02321_, _01411_, _10513_);
  or (_02322_, _02321_, _02320_);
  and (_02323_, _01389_, _10232_);
  and (_02324_, _01425_, _10191_);
  and (_02325_, _01420_, _10798_);
  or (_02326_, _02325_, _02324_);
  and (_02327_, _01427_, _10355_);
  and (_02328_, _01422_, _10570_);
  or (_02329_, _02328_, _02327_);
  or (_02330_, _02329_, _02326_);
  or (_02331_, _02330_, _02323_);
  or (_02332_, _02331_, _02322_);
  or (_02333_, _02332_, _02317_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02333_, _02310_);
  and (_02334_, _01417_, _10691_);
  and (_02335_, _01402_, _10897_);
  or (_02336_, _02335_, _02334_);
  and (_02337_, _01397_, _10278_);
  and (_02338_, _01404_, _10748_);
  or (_02339_, _02338_, _02337_);
  or (_02340_, _02339_, _02336_);
  and (_02341_, _01389_, _10237_);
  and (_02342_, _01386_, _10856_);
  or (_02343_, _02342_, _02341_);
  and (_02344_, _01399_, _10938_);
  and (_02345_, _01392_, _10633_);
  or (_02346_, _02345_, _02344_);
  or (_02347_, _02346_, _02343_);
  and (_02348_, _01409_, _10409_);
  and (_02349_, _01413_, _10464_);
  or (_02350_, _02349_, _02348_);
  and (_02351_, _01411_, _10520_);
  or (_02352_, _02351_, _02350_);
  and (_02353_, _01379_, _10319_);
  and (_02354_, _01425_, _10196_);
  and (_02355_, _01420_, _10805_);
  or (_02356_, _02355_, _02354_);
  and (_02357_, _01427_, _10360_);
  and (_02358_, _01422_, _10577_);
  or (_02359_, _02358_, _02357_);
  or (_02360_, _02359_, _02356_);
  or (_02361_, _02360_, _02353_);
  or (_02362_, _02361_, _02352_);
  or (_02363_, _02362_, _02347_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02363_, _02340_);
  not (_02364_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_02365_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_02366_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_02367_, _02366_, _02365_);
  and (_02368_, _02367_, _10923_);
  not (_02369_, \oc8051_golden_model_1.PC [0]);
  nor (_02370_, \oc8051_golden_model_1.PC [1], _02369_);
  not (_02371_, \oc8051_golden_model_1.PC [3]);
  and (_02372_, \oc8051_golden_model_1.PC [2], _02371_);
  and (_02373_, _02372_, _02370_);
  and (_02374_, _02373_, _10389_);
  nor (_02375_, _02374_, _02368_);
  nor (_02376_, \oc8051_golden_model_1.PC [2], _02371_);
  and (_02377_, _02376_, _02365_);
  and (_02378_, _02377_, _10727_);
  and (_02379_, _02376_, _02370_);
  and (_02380_, _02379_, _10614_);
  nor (_02381_, _02380_, _02378_);
  and (_02382_, _02381_, _02375_);
  and (_02383_, \oc8051_golden_model_1.PC [1], _02369_);
  and (_02384_, _02383_, _02366_);
  and (_02385_, _02384_, _10882_);
  nor (_02386_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  and (_02387_, _02372_, _02386_);
  and (_02388_, _02387_, _10345_);
  nor (_02389_, _02388_, _02385_);
  and (_02390_, _02365_, \oc8051_golden_model_1.PC [2]);
  and (_02391_, _02390_, _02371_);
  and (_02392_, _02391_, _10500_);
  and (_02393_, _02372_, _02383_);
  and (_02394_, _02393_, _10443_);
  nor (_02395_, _02394_, _02392_);
  and (_02396_, _02395_, _02389_);
  and (_02397_, _02396_, _02382_);
  nor (_02398_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  and (_02399_, _02398_, _02383_);
  and (_02400_, _02399_, _10263_);
  and (_02401_, _02398_, _02370_);
  and (_02402_, _02401_, _10222_);
  nor (_02403_, _02402_, _02400_);
  and (_02404_, _02376_, _02383_);
  and (_02405_, _02404_, _10670_);
  and (_02406_, _02386_, _02376_);
  and (_02407_, _02406_, _10556_);
  nor (_02408_, _02407_, _02405_);
  and (_02409_, _02408_, _02403_);
  and (_02410_, _02370_, _02366_);
  and (_02411_, _02410_, _10841_);
  and (_02412_, _02398_, _02386_);
  and (_02413_, _02412_, _10181_);
  nor (_02414_, _02413_, _02411_);
  and (_02415_, _02386_, _02366_);
  and (_02416_, _02415_, _10784_);
  and (_02417_, _02398_, _02365_);
  and (_02418_, _02417_, _10304_);
  nor (_02419_, _02418_, _02416_);
  and (_02420_, _02419_, _02414_);
  and (_02421_, _02420_, _02409_);
  and (_02422_, _02421_, _02397_);
  not (_02423_, _02422_);
  and (_02424_, _02373_, _10383_);
  and (_02425_, _02412_, _10176_);
  nor (_02426_, _02425_, _02424_);
  and (_02427_, _02417_, _10299_);
  and (_02428_, _02401_, _10217_);
  nor (_02429_, _02428_, _02427_);
  and (_02430_, _02429_, _02426_);
  and (_02431_, _02410_, _10834_);
  and (_02432_, _02384_, _10877_);
  nor (_02433_, _02432_, _02431_);
  and (_02434_, _02367_, _10918_);
  and (_02435_, _02406_, _10549_);
  nor (_02436_, _02435_, _02434_);
  and (_02437_, _02436_, _02433_);
  and (_02438_, _02437_, _02430_);
  and (_02439_, _02415_, _10777_);
  and (_02440_, _02377_, _10720_);
  nor (_02441_, _02440_, _02439_);
  and (_02442_, _02379_, _10606_);
  and (_02443_, _02387_, _10340_);
  nor (_02444_, _02443_, _02442_);
  and (_02445_, _02444_, _02441_);
  and (_02446_, _02391_, _10493_);
  and (_02447_, _02393_, _10437_);
  nor (_02448_, _02447_, _02446_);
  and (_02449_, _02404_, _10663_);
  and (_02450_, _02399_, _10258_);
  nor (_02451_, _02450_, _02449_);
  and (_02452_, _02451_, _02448_);
  and (_02453_, _02452_, _02445_);
  and (_02454_, _02453_, _02438_);
  and (_02455_, _02454_, _02423_);
  and (_02456_, _02404_, _10691_);
  and (_02457_, _02401_, _10237_);
  nor (_02458_, _02457_, _02456_);
  and (_02459_, _02377_, _10748_);
  and (_02460_, _02399_, _10278_);
  nor (_02461_, _02460_, _02459_);
  and (_02462_, _02461_, _02458_);
  and (_02463_, _02384_, _10897_);
  and (_02464_, _02387_, _10360_);
  nor (_02465_, _02464_, _02463_);
  and (_02466_, _02367_, _10938_);
  and (_02467_, _02410_, _10856_);
  nor (_02468_, _02467_, _02466_);
  and (_02469_, _02468_, _02465_);
  and (_02470_, _02469_, _02462_);
  and (_02471_, _02373_, _10409_);
  and (_02472_, _02417_, _10319_);
  nor (_02473_, _02472_, _02471_);
  and (_02474_, _02415_, _10805_);
  and (_02475_, _02406_, _10577_);
  nor (_02476_, _02475_, _02474_);
  and (_02477_, _02476_, _02473_);
  and (_02478_, _02391_, _10520_);
  and (_02479_, _02412_, _10196_);
  nor (_02480_, _02479_, _02478_);
  and (_02481_, _02379_, _10633_);
  and (_02482_, _02393_, _10464_);
  nor (_02483_, _02482_, _02481_);
  and (_02484_, _02483_, _02480_);
  and (_02485_, _02484_, _02477_);
  and (_02486_, _02485_, _02470_);
  not (_02487_, _02486_);
  and (_02488_, _02377_, _10699_);
  and (_02489_, _02391_, _10472_);
  nor (_02490_, _02489_, _02488_);
  and (_02491_, _02417_, _10284_);
  and (_02492_, _02401_, _10202_);
  nor (_02493_, _02492_, _02491_);
  and (_02494_, _02493_, _02490_);
  and (_02495_, _02410_, _10814_);
  and (_02496_, _02404_, _10642_);
  nor (_02497_, _02496_, _02495_);
  and (_02498_, _02367_, _10903_);
  and (_02499_, _02379_, _10586_);
  nor (_02500_, _02499_, _02498_);
  and (_02501_, _02500_, _02497_);
  and (_02502_, _02501_, _02494_);
  and (_02503_, _02393_, _10416_);
  and (_02504_, _02387_, _10325_);
  nor (_02505_, _02504_, _02503_);
  and (_02506_, _02412_, _10161_);
  and (_02507_, _02399_, _10243_);
  nor (_02508_, _02507_, _02506_);
  and (_02509_, _02508_, _02505_);
  and (_02510_, _02384_, _10862_);
  and (_02511_, _02415_, _10756_);
  nor (_02512_, _02511_, _02510_);
  and (_02513_, _02406_, _10528_);
  and (_02514_, _02373_, _10366_);
  nor (_02515_, _02514_, _02513_);
  and (_02516_, _02515_, _02512_);
  and (_02517_, _02516_, _02509_);
  and (_02518_, _02517_, _02502_);
  and (_02519_, _02518_, _02487_);
  and (_02520_, _02519_, _02455_);
  and (_02521_, _02406_, _10535_);
  and (_02522_, _02417_, _10289_);
  nor (_02523_, _02522_, _02521_);
  and (_02524_, _02377_, _10706_);
  and (_02525_, _02379_, _10592_);
  nor (_02526_, _02525_, _02524_);
  and (_02527_, _02526_, _02523_);
  and (_02528_, _02415_, _10763_);
  and (_02529_, _02393_, _10423_);
  nor (_02530_, _02529_, _02528_);
  and (_02531_, _02391_, _10479_);
  and (_02532_, _02373_, _10371_);
  nor (_02533_, _02532_, _02531_);
  and (_02534_, _02533_, _02530_);
  and (_02535_, _02534_, _02527_);
  and (_02536_, _02410_, _10820_);
  and (_02537_, _02399_, _10248_);
  nor (_02538_, _02537_, _02536_);
  and (_02539_, _02387_, _10330_);
  and (_02540_, _02412_, _10166_);
  nor (_02541_, _02540_, _02539_);
  and (_02542_, _02541_, _02538_);
  and (_02543_, _02367_, _10908_);
  and (_02544_, _02401_, _10207_);
  nor (_02545_, _02544_, _02543_);
  and (_02546_, _02384_, _10867_);
  and (_02547_, _02404_, _10649_);
  nor (_02548_, _02547_, _02546_);
  and (_02549_, _02548_, _02545_);
  and (_02550_, _02549_, _02542_);
  and (_02551_, _02550_, _02535_);
  not (_02552_, _02551_);
  and (_02553_, _02410_, _10827_);
  and (_02554_, _02391_, _10486_);
  nor (_02555_, _02554_, _02553_);
  and (_02556_, _02377_, _10713_);
  and (_02557_, _02399_, _10253_);
  nor (_02558_, _02557_, _02556_);
  and (_02559_, _02558_, _02555_);
  and (_02560_, _02415_, _10770_);
  and (_02561_, _02393_, _10430_);
  nor (_02562_, _02561_, _02560_);
  and (_02563_, _02367_, _10913_);
  and (_02564_, _02384_, _10872_);
  nor (_02565_, _02564_, _02563_);
  and (_02566_, _02565_, _02562_);
  and (_02567_, _02566_, _02559_);
  and (_02568_, _02404_, _10656_);
  and (_02569_, _02379_, _10599_);
  nor (_02570_, _02569_, _02568_);
  and (_02571_, _02417_, _10294_);
  and (_02572_, _02412_, _10171_);
  nor (_02573_, _02572_, _02571_);
  and (_02574_, _02573_, _02570_);
  and (_02575_, _02406_, _10542_);
  and (_02576_, _02373_, _10377_);
  nor (_02577_, _02576_, _02575_);
  and (_02578_, _02387_, _10335_);
  and (_02579_, _02401_, _10212_);
  nor (_02580_, _02579_, _02578_);
  and (_02581_, _02580_, _02577_);
  and (_02582_, _02581_, _02574_);
  and (_02583_, _02582_, _02567_);
  and (_02584_, _02583_, _02552_);
  and (_02585_, _02406_, _10563_);
  and (_02586_, _02417_, _10309_);
  nor (_02587_, _02586_, _02585_);
  and (_02588_, _02377_, _10734_);
  and (_02589_, _02379_, _10619_);
  nor (_02590_, _02589_, _02588_);
  and (_02591_, _02590_, _02587_);
  and (_02592_, _02415_, _10791_);
  and (_02593_, _02393_, _10450_);
  nor (_02594_, _02593_, _02592_);
  and (_02595_, _02391_, _10506_);
  and (_02596_, _02373_, _10396_);
  nor (_02597_, _02596_, _02595_);
  and (_02598_, _02597_, _02594_);
  and (_02599_, _02598_, _02591_);
  and (_02600_, _02410_, _10846_);
  and (_02601_, _02399_, _10268_);
  nor (_02602_, _02601_, _02600_);
  and (_02603_, _02387_, _10350_);
  and (_02604_, _02412_, _10186_);
  nor (_02605_, _02604_, _02603_);
  and (_02606_, _02605_, _02602_);
  and (_02607_, _02367_, _10928_);
  and (_02608_, _02401_, _10227_);
  nor (_02609_, _02608_, _02607_);
  and (_02610_, _02384_, _10887_);
  and (_02611_, _02404_, _10677_);
  nor (_02612_, _02611_, _02610_);
  and (_02613_, _02612_, _02609_);
  and (_02614_, _02613_, _02606_);
  and (_02615_, _02614_, _02599_);
  and (_02616_, _02410_, _10851_);
  and (_02617_, _02391_, _10513_);
  nor (_02618_, _02617_, _02616_);
  and (_02619_, _02377_, _10741_);
  and (_02620_, _02399_, _10273_);
  nor (_02621_, _02620_, _02619_);
  and (_02622_, _02621_, _02618_);
  and (_02623_, _02415_, _10798_);
  and (_02624_, _02393_, _10457_);
  nor (_02625_, _02624_, _02623_);
  and (_02626_, _02367_, _10933_);
  and (_02627_, _02384_, _10892_);
  nor (_02628_, _02627_, _02626_);
  and (_02629_, _02628_, _02625_);
  and (_02630_, _02629_, _02622_);
  and (_02631_, _02404_, _10684_);
  and (_02632_, _02379_, _10626_);
  nor (_02633_, _02632_, _02631_);
  and (_02634_, _02417_, _10314_);
  and (_02635_, _02412_, _10191_);
  nor (_02636_, _02635_, _02634_);
  and (_02637_, _02636_, _02633_);
  and (_02638_, _02406_, _10570_);
  and (_02639_, _02373_, _10402_);
  nor (_02640_, _02639_, _02638_);
  and (_02641_, _02387_, _10355_);
  and (_02642_, _02401_, _10232_);
  nor (_02643_, _02642_, _02641_);
  and (_02644_, _02643_, _02640_);
  and (_02645_, _02644_, _02637_);
  and (_02646_, _02645_, _02630_);
  and (_02647_, _02646_, _02615_);
  and (_02648_, _02647_, _02584_);
  and (_02649_, _02648_, _02520_);
  nand (_02650_, _00002_, WR_COND_ABSTR_IRAM_0);
  nor (_02651_, _02650_, _02649_);
  and (_02652_, _02651_, WR_ADDR_ABSTR_IRAM_0[2]);
  and (_02653_, _02652_, WR_ADDR_ABSTR_IRAM_0[3]);
  and (_02654_, _02651_, WR_ADDR_ABSTR_IRAM_0[1]);
  and (_02655_, _02654_, WR_ADDR_ABSTR_IRAM_0[0]);
  and (_02656_, _02655_, _02653_);
  nor (_02657_, _02656_, _02364_);
  and (_02658_, _02651_, WR_DATA_ABSTR_IRAM_0[7]);
  and (_02659_, _02658_, _02656_);
  or (_02660_, _02659_, _02657_);
  nand (_02661_, _00002_, WR_COND_ABSTR_IRAM_1);
  nor (_02662_, _02661_, _02649_);
  and (_02663_, _02662_, WR_ADDR_ABSTR_IRAM_1[1]);
  and (_02664_, _02663_, WR_ADDR_ABSTR_IRAM_1[0]);
  and (_02665_, _02662_, WR_ADDR_ABSTR_IRAM_1[2]);
  and (_02666_, _02665_, WR_ADDR_ABSTR_IRAM_1[3]);
  and (_02667_, _02666_, _02664_);
  not (_02668_, _02667_);
  and (_02669_, _02668_, _02660_);
  and (_02670_, _02662_, WR_DATA_ABSTR_IRAM_1[7]);
  and (_02671_, _02670_, _02667_);
  or (_12667_[7], _02671_, _02669_);
  not (_02672_, _02649_);
  and (_02673_, _02672_, XRAM_DATA_OUT_abstr[7]);
  or (_02674_, _02673_, _11613_);
  or (_02675_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [7]);
  and (_02676_, _02675_, _12493_);
  and (_12635_[7], _02676_, _02674_);
  and (_02677_, _02367_, \oc8051_golden_model_1.PC [4]);
  and (_02678_, _02677_, \oc8051_golden_model_1.PC [5]);
  and (_02679_, _02678_, \oc8051_golden_model_1.PC [6]);
  and (_02680_, _02679_, \oc8051_golden_model_1.PC [7]);
  and (_02681_, _02680_, \oc8051_golden_model_1.PC [8]);
  and (_02682_, _02681_, \oc8051_golden_model_1.PC [9]);
  and (_02683_, _02682_, \oc8051_golden_model_1.PC [10]);
  and (_02684_, _02683_, \oc8051_golden_model_1.PC [11]);
  and (_02685_, _02684_, \oc8051_golden_model_1.PC [12]);
  and (_02686_, _02685_, \oc8051_golden_model_1.PC [13]);
  and (_02687_, _02686_, \oc8051_golden_model_1.PC [14]);
  nor (_02688_, _02687_, \oc8051_golden_model_1.PC [15]);
  and (_02689_, _02687_, \oc8051_golden_model_1.PC [15]);
  or (_02690_, _02689_, _02688_);
  nor (_02691_, _02690_, _02672_);
  and (_02692_, _02672_, PC_abstr[15]);
  nor (_02693_, _02692_, _02691_);
  nand (_02694_, _02693_, _11609_);
  or (_02695_, _11609_, \oc8051_golden_model_1.PC [15]);
  and (_02696_, _02695_, _12493_);
  and (_12623_[15], _02696_, _02694_);
  and (_02697_, _02672_, XRAM_ADDR_abstr[15]);
  or (_02698_, _02697_, _11613_);
  or (_02699_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [15]);
  and (_02700_, _02699_, _12493_);
  and (_12634_[15], _02700_, _02698_);
  and (_12633_[7], \oc8051_golden_model_1.TMOD [7], _12493_);
  and (_12632_[7], \oc8051_golden_model_1.TL1 [7], _12493_);
  and (_12631_[7], \oc8051_golden_model_1.TL0 [7], _12493_);
  and (_12630_[7], \oc8051_golden_model_1.TH1 [7], _12493_);
  and (_12629_[7], \oc8051_golden_model_1.TH0 [7], _12493_);
  and (_12628_[7], \oc8051_golden_model_1.TCON [7], _12493_);
  nor (_02701_, _02649_, _11613_);
  and (_02702_, _02701_, SP_abstr[7]);
  not (_02703_, \oc8051_golden_model_1.SP [7]);
  nor (_02704_, _02701_, _02703_);
  or (_02705_, _02704_, _02702_);
  and (_12627_[7], _02705_, _12493_);
  and (_12626_[7], \oc8051_golden_model_1.SCON [7], _12493_);
  and (_12625_[7], \oc8051_golden_model_1.SBUF [7], _12493_);
  and (_12622_[7], \oc8051_golden_model_1.PCON [7], _12493_);
  not (_02706_, \oc8051_golden_model_1.PSW [7]);
  nor (_02707_, _02701_, _02706_);
  and (_02708_, _02701_, PSW_abstr[7]);
  or (_02709_, _02708_, _02707_);
  and (_12624_[7], _02709_, _12493_);
  and (_02710_, _02701_, P3_abstr[7]);
  not (_02711_, \oc8051_golden_model_1.P3 [7]);
  nor (_02712_, _02701_, _02711_);
  or (_02713_, _02712_, rst);
  or (_12621_[7], _02713_, _02710_);
  and (_02714_, _02701_, P2_abstr[7]);
  not (_02715_, \oc8051_golden_model_1.P2 [7]);
  nor (_02716_, _02701_, _02715_);
  or (_02717_, _02716_, rst);
  or (_12620_[7], _02717_, _02714_);
  and (_02718_, _02701_, P1_abstr[7]);
  not (_02719_, \oc8051_golden_model_1.P1 [7]);
  nor (_02720_, _02701_, _02719_);
  or (_02721_, _02720_, rst);
  or (_12619_[7], _02721_, _02718_);
  and (_02722_, _02701_, P0_abstr[7]);
  not (_02723_, \oc8051_golden_model_1.P0 [7]);
  nor (_02724_, _02701_, _02723_);
  or (_02725_, _02724_, rst);
  or (_12618_[7], _02725_, _02722_);
  and (_12617_[7], \oc8051_golden_model_1.IP [7], _12493_);
  and (_12616_[7], \oc8051_golden_model_1.IE [7], _12493_);
  and (_02726_, _02701_, DPH_abstr[7]);
  not (_02727_, \oc8051_golden_model_1.DPH [7]);
  nor (_02728_, _02701_, _02727_);
  or (_02729_, _02728_, _02726_);
  and (_12614_[7], _02729_, _12493_);
  and (_02730_, _02701_, DPL_abstr[7]);
  not (_02731_, \oc8051_golden_model_1.DPL [7]);
  nor (_02733_, _02701_, _02731_);
  or (_02734_, _02733_, _02730_);
  and (_12615_[7], _02734_, _12493_);
  not (_02735_, \oc8051_golden_model_1.ACC [7]);
  nor (_02736_, _11609_, _02735_);
  and (_02737_, _02672_, RD_IRAM_0_ABSTR_ADDR[2]);
  nor (_02738_, _02649_, RD_IRAM_0_ABSTR_ADDR[0]);
  not (_02739_, _02738_);
  or (_02740_, _02739_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_02741_, _02672_, RD_IRAM_0_ABSTR_ADDR[1]);
  nor (_02742_, _02738_, \oc8051_golden_model_1.IRAM[5] [7]);
  nor (_02743_, _02742_, _02741_);
  and (_02744_, _02743_, _02740_);
  and (_02745_, _02738_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_02746_, _02739_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_02747_, _02746_, _02745_);
  and (_02748_, _02747_, _02741_);
  nor (_02749_, _02748_, _02744_);
  nand (_02750_, _02749_, _02737_);
  and (_02751_, _02672_, RD_IRAM_0_ABSTR_ADDR[3]);
  and (_02752_, _02649_, \oc8051_golden_model_1.PSW [3]);
  nor (_02753_, _02752_, _02751_);
  not (_02754_, _02737_);
  or (_02755_, _02739_, \oc8051_golden_model_1.IRAM[0] [7]);
  nor (_02756_, _02738_, \oc8051_golden_model_1.IRAM[1] [7]);
  nor (_02757_, _02756_, _02741_);
  and (_02758_, _02757_, _02755_);
  and (_02759_, _02738_, \oc8051_golden_model_1.IRAM[2] [7]);
  not (_02760_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor (_02761_, _02738_, _02760_);
  or (_02762_, _02761_, _02759_);
  and (_02763_, _02762_, _02741_);
  nor (_02764_, _02763_, _02758_);
  nand (_02765_, _02764_, _02754_);
  and (_02766_, _02765_, _02753_);
  and (_02767_, _02766_, _02750_);
  not (_02768_, _02753_);
  or (_02769_, _02739_, \oc8051_golden_model_1.IRAM[8] [7]);
  nor (_02770_, _02738_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor (_02771_, _02770_, _02741_);
  and (_02772_, _02771_, _02769_);
  and (_02773_, _02738_, \oc8051_golden_model_1.IRAM[10] [7]);
  not (_02774_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_02775_, _02738_, _02774_);
  or (_02776_, _02775_, _02773_);
  and (_02777_, _02776_, _02741_);
  nor (_02778_, _02777_, _02772_);
  nor (_02779_, _02778_, _02737_);
  nor (_02780_, _02739_, \oc8051_golden_model_1.IRAM[12] [7]);
  nor (_02781_, _02738_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_02782_, _02781_, _02741_);
  nor (_02783_, _02782_, _02780_);
  and (_02784_, _02738_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_02785_, _02738_, _02364_);
  or (_02786_, _02785_, _02784_);
  and (_02787_, _02786_, _02741_);
  nor (_02788_, _02787_, _02783_);
  nor (_02789_, _02788_, _02754_);
  or (_02790_, _02789_, _02779_);
  and (_02791_, _02790_, _02768_);
  or (_02792_, _02791_, _02767_);
  nor (_02793_, _02792_, \oc8051_golden_model_1.ACC [7]);
  and (_02794_, _02793_, _02649_);
  or (_02795_, _02649_, ACC_abstr[7]);
  nand (_02796_, _02795_, _11609_);
  nor (_02797_, _02796_, _02794_);
  or (_02798_, _02797_, _02736_);
  and (_12612_[7], _02798_, _12493_);
  and (_02799_, _02701_, B_abstr[7]);
  not (_02800_, \oc8051_golden_model_1.B [7]);
  nor (_02801_, _02701_, _02800_);
  or (_02802_, _02801_, _02799_);
  and (_12613_[7], _02802_, _12493_);
  and (_02803_, _02662_, WR_ADDR_ABSTR_IRAM_1[0]);
  nor (_02804_, _02803_, _02663_);
  and (_02805_, _02662_, WR_ADDR_ABSTR_IRAM_1[3]);
  nor (_02806_, _02805_, _02665_);
  and (_02807_, _02806_, _02804_);
  and (_02808_, _02807_, _02662_);
  not (_02809_, _02808_);
  not (_02810_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_02811_, _02651_, WR_ADDR_ABSTR_IRAM_0[3]);
  nor (_02812_, _02811_, _02652_);
  and (_02813_, _02651_, WR_ADDR_ABSTR_IRAM_0[0]);
  nor (_02814_, _02813_, _02654_);
  and (_02815_, _02814_, _02812_);
  and (_02816_, _02815_, _02651_);
  nor (_02817_, _02816_, _02810_);
  and (_02818_, _02816_, WR_DATA_ABSTR_IRAM_0[0]);
  or (_02819_, _02818_, _02817_);
  and (_02820_, _02819_, _02809_);
  and (_02821_, _02808_, WR_DATA_ABSTR_IRAM_1[0]);
  or (_12636_, _02821_, _02820_);
  not (_02822_, \oc8051_golden_model_1.IRAM[0] [1]);
  nor (_02823_, _02816_, _02822_);
  and (_02824_, _02651_, WR_DATA_ABSTR_IRAM_0[1]);
  and (_02825_, _02824_, _02815_);
  or (_02826_, _02825_, _02823_);
  and (_02827_, _02826_, _02809_);
  and (_02828_, _02808_, WR_DATA_ABSTR_IRAM_1[1]);
  or (_12637_, _02828_, _02827_);
  not (_02829_, _02816_);
  and (_02830_, _02829_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_02831_, _02651_, WR_DATA_ABSTR_IRAM_0[2]);
  and (_02832_, _02831_, _02816_);
  or (_02833_, _02832_, _02830_);
  and (_02834_, _02833_, _02809_);
  and (_02835_, _02808_, WR_DATA_ABSTR_IRAM_1[2]);
  or (_12638_, _02835_, _02834_);
  or (_02836_, _02829_, WR_DATA_ABSTR_IRAM_0[3]);
  or (_02837_, _02816_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_02838_, _02837_, _02836_);
  or (_02839_, _02838_, _02808_);
  or (_02840_, _02809_, WR_DATA_ABSTR_IRAM_1[3]);
  and (_12639_, _02840_, _02839_);
  or (_02841_, _02829_, WR_DATA_ABSTR_IRAM_0[4]);
  or (_02842_, _02816_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_02843_, _02842_, _02841_);
  or (_02844_, _02843_, _02808_);
  or (_02845_, _02809_, WR_DATA_ABSTR_IRAM_1[4]);
  and (_12640_, _02845_, _02844_);
  or (_02846_, _02816_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_02847_, _02829_, WR_DATA_ABSTR_IRAM_0[5]);
  and (_02848_, _02847_, _02809_);
  and (_02849_, _02848_, _02846_);
  and (_02850_, _02662_, WR_DATA_ABSTR_IRAM_1[5]);
  and (_02851_, _02850_, _02807_);
  or (_12641_, _02851_, _02849_);
  or (_02852_, _02829_, WR_DATA_ABSTR_IRAM_0[6]);
  or (_02853_, _02816_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_02854_, _02853_, _02852_);
  or (_02855_, _02854_, _02808_);
  or (_02856_, _02809_, WR_DATA_ABSTR_IRAM_1[6]);
  and (_12642_, _02856_, _02855_);
  and (_02857_, _02807_, _02670_);
  or (_02858_, _02816_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_02859_, _02829_, WR_DATA_ABSTR_IRAM_0[7]);
  and (_02860_, _02859_, _02809_);
  and (_02861_, _02860_, _02858_);
  or (_12643_, _02861_, _02857_);
  not (_02862_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_02863_, WR_ADDR_ABSTR_IRAM_0[1]);
  and (_02864_, _02813_, _02863_);
  and (_02865_, _02864_, _02812_);
  nor (_02866_, _02865_, _02862_);
  and (_02867_, _02651_, WR_DATA_ABSTR_IRAM_0[0]);
  and (_02868_, _02867_, _02865_);
  nor (_02869_, _02868_, _02866_);
  not (_02870_, WR_ADDR_ABSTR_IRAM_1[1]);
  and (_02871_, _02803_, _02870_);
  and (_02872_, _02871_, _02806_);
  nor (_02873_, _02872_, _02869_);
  and (_02874_, _02662_, WR_DATA_ABSTR_IRAM_1[0]);
  and (_02875_, _02872_, _02874_);
  or (_12644_, _02875_, _02873_);
  and (_02876_, _02672_, WR_COND_ABSTR_IRAM_1);
  and (_02877_, _02876_, WR_ADDR_ABSTR_IRAM_1[2]);
  and (_02878_, _02877_, _11609_);
  and (_02879_, _02878_, _12493_);
  and (_02880_, _02876_, WR_ADDR_ABSTR_IRAM_1[3]);
  and (_02881_, _02880_, _11609_);
  and (_02882_, _02881_, _12493_);
  or (_02883_, _02882_, _02879_);
  and (_02884_, _02876_, WR_ADDR_ABSTR_IRAM_1[0]);
  and (_02885_, _02884_, _11609_);
  and (_02886_, _02885_, _12493_);
  and (_02887_, _02876_, WR_ADDR_ABSTR_IRAM_1[1]);
  and (_02888_, _02887_, _11609_);
  and (_02889_, _02888_, _12493_);
  not (_02890_, _02889_);
  nand (_02891_, _02890_, _02886_);
  or (_02892_, _02891_, _02883_);
  not (_02893_, _02865_);
  or (_02894_, _02893_, _02824_);
  or (_02895_, _02865_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_02896_, _02895_, _02894_);
  and (_02897_, _02896_, _02892_);
  and (_02898_, _02662_, WR_DATA_ABSTR_IRAM_1[1]);
  and (_02899_, _02872_, _02898_);
  or (_12645_, _02899_, _02897_);
  or (_02900_, _02893_, _02831_);
  or (_02901_, _02865_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_02902_, _02901_, _02900_);
  and (_02903_, _02902_, _02892_);
  and (_02904_, _02662_, WR_DATA_ABSTR_IRAM_1[2]);
  and (_02905_, _02904_, _02872_);
  or (_12646_, _02905_, _02903_);
  and (_02906_, _02651_, WR_DATA_ABSTR_IRAM_0[3]);
  or (_02907_, _02906_, _02893_);
  or (_02908_, _02865_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_02909_, _02908_, _02907_);
  and (_02910_, _02909_, _02892_);
  and (_02911_, _02662_, WR_DATA_ABSTR_IRAM_1[3]);
  and (_02912_, _02872_, _02911_);
  or (_12647_, _02912_, _02910_);
  and (_02913_, _02651_, WR_DATA_ABSTR_IRAM_0[4]);
  or (_02914_, _02913_, _02893_);
  or (_02915_, _02865_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_02916_, _02915_, _02914_);
  and (_02917_, _02916_, _02892_);
  and (_02919_, _02662_, WR_DATA_ABSTR_IRAM_1[4]);
  and (_02920_, _02872_, _02919_);
  or (_12648_, _02920_, _02917_);
  and (_02921_, _02651_, WR_DATA_ABSTR_IRAM_0[5]);
  or (_02922_, _02893_, _02921_);
  or (_02923_, _02865_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_02924_, _02923_, _02922_);
  and (_02925_, _02924_, _02892_);
  and (_02926_, _02872_, _02850_);
  or (_12649_, _02926_, _02925_);
  and (_02927_, _02651_, WR_DATA_ABSTR_IRAM_0[6]);
  or (_02928_, _02927_, _02893_);
  or (_02929_, _02865_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_02930_, _02929_, _02928_);
  and (_02931_, _02930_, _02892_);
  and (_02932_, _02662_, WR_DATA_ABSTR_IRAM_1[6]);
  and (_02933_, _02872_, _02932_);
  or (_12650_, _02933_, _02931_);
  or (_02934_, _02893_, _02658_);
  or (_02935_, _02865_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_02936_, _02935_, _02934_);
  and (_02937_, _02936_, _02892_);
  and (_02938_, _02872_, _02670_);
  or (_12651_, _02938_, _02937_);
  not (_02939_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_02940_, WR_ADDR_ABSTR_IRAM_0[0]);
  and (_02941_, _02654_, _02940_);
  and (_02942_, _02941_, _02812_);
  nor (_02943_, _02942_, _02939_);
  and (_02944_, _02942_, _02867_);
  nor (_02945_, _02944_, _02943_);
  not (_02946_, WR_ADDR_ABSTR_IRAM_1[0]);
  and (_02947_, _02663_, _02946_);
  and (_02948_, _02947_, _02806_);
  nor (_02949_, _02948_, _02945_);
  and (_02950_, _02948_, _02874_);
  or (_12652_, _02950_, _02949_);
  or (_02951_, _02890_, _02886_);
  or (_02952_, _02951_, _02883_);
  not (_02953_, _02942_);
  or (_02954_, _02953_, _02824_);
  or (_02955_, _02942_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_02956_, _02955_, _02954_);
  and (_02957_, _02956_, _02952_);
  and (_02958_, _02948_, _02898_);
  or (_12653_, _02958_, _02957_);
  or (_02959_, _02953_, _02831_);
  or (_02960_, _02942_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_02961_, _02960_, _02959_);
  and (_02962_, _02961_, _02952_);
  and (_02963_, _02948_, _02904_);
  or (_12654_, _02963_, _02962_);
  or (_02964_, _02953_, _02906_);
  or (_02965_, _02942_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_02966_, _02965_, _02964_);
  and (_02967_, _02966_, _02952_);
  and (_02968_, _02948_, _02911_);
  or (_12655_, _02968_, _02967_);
  or (_02969_, _02953_, _02913_);
  or (_02970_, _02942_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_02972_, _02970_, _02969_);
  and (_02973_, _02972_, _02952_);
  and (_02974_, _02948_, _02919_);
  or (_12656_, _02974_, _02973_);
  or (_02975_, _02953_, _02921_);
  or (_02976_, _02942_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_02977_, _02976_, _02975_);
  and (_02978_, _02977_, _02952_);
  and (_02979_, _02948_, _02850_);
  or (_12657_, _02979_, _02978_);
  or (_02981_, _02953_, _02927_);
  or (_02982_, _02942_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_02983_, _02982_, _02981_);
  and (_02984_, _02983_, _02952_);
  and (_02985_, _02948_, _02932_);
  or (_12658_, _02985_, _02984_);
  or (_02986_, _02953_, _02658_);
  or (_02987_, _02942_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_02988_, _02987_, _02986_);
  and (_02989_, _02988_, _02952_);
  and (_02990_, _02948_, _02670_);
  or (_12659_, _02990_, _02989_);
  not (_02991_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_02992_, _02812_, _02655_);
  nor (_02993_, _02992_, _02991_);
  and (_02994_, _02992_, _02867_);
  nor (_02995_, _02994_, _02993_);
  and (_02996_, _02806_, _02664_);
  nor (_02997_, _02996_, _02995_);
  and (_02998_, _02996_, _02874_);
  or (_12660_, _02998_, _02997_);
  nand (_03000_, _02889_, _02886_);
  or (_03001_, _02883_, _03000_);
  not (_03002_, _02992_);
  or (_03003_, _03002_, _02824_);
  or (_03004_, _02992_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_03005_, _03004_, _03003_);
  and (_03006_, _03005_, _03001_);
  and (_03007_, _02803_, WR_ADDR_ABSTR_IRAM_1[1]);
  and (_03008_, _02806_, _03007_);
  and (_03009_, _03008_, _02898_);
  or (_12661_, _03009_, _03006_);
  or (_03010_, _03002_, _02831_);
  or (_03011_, _02992_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_03012_, _03011_, _03010_);
  and (_03013_, _03012_, _03001_);
  and (_03014_, _03008_, _02904_);
  or (_12668_[2], _03014_, _03013_);
  or (_03015_, _03002_, _02906_);
  or (_03016_, _02992_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_03018_, _03016_, _03015_);
  and (_03019_, _03018_, _03001_);
  and (_03020_, _03008_, _02911_);
  or (_12668_[3], _03020_, _03019_);
  or (_03021_, _03002_, _02913_);
  or (_03022_, _02992_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_03023_, _03022_, _03021_);
  and (_03024_, _03023_, _03001_);
  and (_03025_, _03008_, _02919_);
  or (_12668_[4], _03025_, _03024_);
  or (_03026_, _03002_, _02921_);
  or (_03027_, _02992_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_03028_, _03027_, _03026_);
  and (_03029_, _03028_, _03001_);
  and (_03030_, _03008_, _02850_);
  or (_12668_[5], _03030_, _03029_);
  or (_03031_, _03002_, _02927_);
  or (_03032_, _02992_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_03033_, _03032_, _03031_);
  and (_03034_, _03033_, _03001_);
  and (_03036_, _03008_, _02932_);
  or (_12668_[6], _03036_, _03034_);
  or (_03037_, _03002_, _02658_);
  or (_03038_, _02992_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_03039_, _03038_, _03037_);
  and (_03040_, _03039_, _03001_);
  and (_03041_, _03008_, _02670_);
  or (_12668_[7], _03041_, _03040_);
  not (_03042_, \oc8051_golden_model_1.IRAM[4] [0]);
  not (_03043_, WR_ADDR_ABSTR_IRAM_0[3]);
  and (_03045_, _02652_, _03043_);
  and (_03046_, _03045_, _02814_);
  nor (_03047_, _03046_, _03042_);
  and (_03048_, _03046_, _02867_);
  nor (_03049_, _03048_, _03047_);
  not (_03050_, WR_ADDR_ABSTR_IRAM_1[3]);
  and (_03051_, _02665_, _03050_);
  and (_03052_, _03051_, _02804_);
  nor (_03053_, _03052_, _03049_);
  and (_03054_, _03052_, _02874_);
  or (_12669_[0], _03054_, _03053_);
  or (_03056_, _02889_, _02886_);
  not (_03057_, _02882_);
  nand (_03058_, _03057_, _02879_);
  or (_03059_, _03058_, _03056_);
  not (_03060_, _03046_);
  or (_03061_, _03060_, _02824_);
  or (_03062_, _03046_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_03063_, _03062_, _03061_);
  and (_03064_, _03063_, _03059_);
  and (_03066_, _03052_, _02898_);
  or (_12669_[1], _03066_, _03064_);
  or (_03067_, _03060_, _02831_);
  or (_03068_, _03046_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_03069_, _03068_, _03067_);
  and (_03070_, _03069_, _03059_);
  and (_03071_, _03052_, _02904_);
  or (_12669_[2], _03071_, _03070_);
  or (_03072_, _03060_, _02906_);
  or (_03073_, _03046_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_03075_, _03073_, _03072_);
  and (_03076_, _03075_, _03059_);
  and (_03077_, _03052_, _02911_);
  or (_12669_[3], _03077_, _03076_);
  or (_03078_, _03060_, _02913_);
  or (_03079_, _03046_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_03080_, _03079_, _03078_);
  and (_03081_, _03080_, _03059_);
  and (_03082_, _03052_, _02919_);
  or (_12669_[4], _03082_, _03081_);
  or (_03084_, _03060_, _02921_);
  or (_03085_, _03046_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_03086_, _03085_, _03084_);
  and (_03087_, _03086_, _03059_);
  and (_03088_, _03052_, _02850_);
  or (_12669_[5], _03088_, _03087_);
  or (_03089_, _03060_, _02927_);
  or (_03090_, _03046_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_03091_, _03090_, _03089_);
  and (_03092_, _03091_, _03059_);
  and (_03094_, _03052_, _02932_);
  or (_12669_[6], _03094_, _03092_);
  or (_03095_, _03060_, _02658_);
  or (_03096_, _03046_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_03097_, _03096_, _03095_);
  and (_03098_, _03097_, _03059_);
  and (_03099_, _03052_, _02670_);
  or (_12669_[7], _03099_, _03098_);
  not (_03100_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_03101_, _03045_, _02864_);
  nor (_03104_, _03101_, _03100_);
  and (_03105_, _03101_, _02867_);
  or (_03106_, _03105_, _03104_);
  and (_03107_, _03051_, _02871_);
  not (_03108_, _03107_);
  and (_03109_, _03108_, _03106_);
  and (_03110_, _03107_, _02874_);
  or (_12670_[0], _03110_, _03109_);
  not (_03111_, _03101_);
  or (_03112_, _03111_, _02824_);
  or (_03114_, _03101_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_03115_, _03114_, _03108_);
  and (_03116_, _03115_, _03112_);
  and (_03117_, _03107_, _02898_);
  or (_12670_[1], _03117_, _03116_);
  or (_03118_, _03111_, _02831_);
  or (_03119_, _03101_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_03120_, _03119_, _03108_);
  and (_03121_, _03120_, _03118_);
  and (_03122_, _03107_, _02904_);
  or (_12670_[2], _03122_, _03121_);
  or (_03123_, _03111_, _02906_);
  or (_03124_, _03101_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_03125_, _03124_, _03108_);
  and (_03126_, _03125_, _03123_);
  and (_03127_, _03107_, _02911_);
  or (_12670_[3], _03127_, _03126_);
  not (_03128_, \oc8051_golden_model_1.IRAM[5] [4]);
  nor (_03129_, _03101_, _03128_);
  and (_03130_, _03101_, _02913_);
  or (_03131_, _03130_, _03129_);
  and (_03132_, _03131_, _03108_);
  and (_03133_, _03107_, _02919_);
  or (_12670_[4], _03133_, _03132_);
  or (_03134_, _03111_, _02921_);
  or (_03135_, _03101_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_03136_, _03135_, _03108_);
  and (_03137_, _03136_, _03134_);
  and (_03138_, _03107_, _02850_);
  or (_12670_[5], _03138_, _03137_);
  or (_03139_, _03111_, _02927_);
  or (_03140_, _03101_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_03141_, _03140_, _03108_);
  and (_03142_, _03141_, _03139_);
  and (_03143_, _03107_, _02932_);
  or (_12670_[6], _03143_, _03142_);
  or (_03144_, _03111_, _02658_);
  or (_03145_, _03101_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_03146_, _03145_, _03108_);
  and (_03147_, _03146_, _03144_);
  and (_03148_, _03107_, _02670_);
  or (_12670_[7], _03148_, _03147_);
  not (_03149_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_03150_, _03045_, _02941_);
  nor (_03151_, _03150_, _03149_);
  and (_03152_, _03150_, _02867_);
  or (_03153_, _03152_, _03151_);
  and (_03154_, _03051_, _02947_);
  not (_03155_, _03154_);
  and (_03156_, _03155_, _03153_);
  and (_03157_, _03154_, _02874_);
  or (_12671_[0], _03157_, _03156_);
  not (_03158_, _03150_);
  or (_03159_, _03158_, _02824_);
  or (_03160_, _03150_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_03161_, _03160_, _03155_);
  and (_03162_, _03161_, _03159_);
  and (_03163_, _03154_, _02898_);
  or (_12671_[1], _03163_, _03162_);
  or (_03164_, _03158_, _02831_);
  or (_03165_, _03150_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_03166_, _03165_, _03155_);
  and (_03167_, _03166_, _03164_);
  and (_03168_, _03154_, _02904_);
  or (_12671_[2], _03168_, _03167_);
  or (_03169_, _03158_, _02906_);
  or (_03170_, _03150_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_03171_, _03170_, _03155_);
  and (_03172_, _03171_, _03169_);
  and (_03173_, _03154_, _02911_);
  or (_12671_[3], _03173_, _03172_);
  or (_03174_, _03158_, _02913_);
  or (_03175_, _03150_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_03176_, _03175_, _03155_);
  and (_03177_, _03176_, _03174_);
  and (_03178_, _03154_, _02919_);
  or (_12671_[4], _03178_, _03177_);
  not (_03179_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor (_03180_, _03150_, _03179_);
  and (_03181_, _03150_, _02921_);
  or (_03182_, _03181_, _03180_);
  and (_03183_, _03182_, _03155_);
  and (_03184_, _03154_, _02850_);
  or (_12671_[5], _03184_, _03183_);
  or (_03185_, _03158_, _02927_);
  or (_03186_, _03150_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_03187_, _03186_, _03155_);
  and (_03188_, _03187_, _03185_);
  and (_03189_, _03154_, _02932_);
  or (_12671_[6], _03189_, _03188_);
  or (_03190_, _03158_, _02658_);
  or (_03191_, _03150_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_03192_, _03191_, _03155_);
  and (_03193_, _03192_, _03190_);
  and (_03194_, _03154_, _02670_);
  or (_12671_[7], _03194_, _03193_);
  not (_03195_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_03196_, _03045_, _02655_);
  nor (_03197_, _03196_, _03195_);
  and (_03198_, _03196_, _02867_);
  nor (_03199_, _03198_, _03197_);
  and (_03200_, _03051_, _02664_);
  nor (_03201_, _03200_, _03199_);
  and (_03202_, _03200_, _02874_);
  or (_12672_[0], _03202_, _03201_);
  or (_03203_, _03058_, _03000_);
  not (_03204_, _03196_);
  or (_03205_, _03204_, _02824_);
  or (_03206_, _03196_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_03207_, _03206_, _03205_);
  and (_03208_, _03207_, _03203_);
  and (_03209_, _03051_, _03007_);
  and (_03210_, _03209_, _02898_);
  or (_12672_[1], _03210_, _03208_);
  or (_03211_, _03204_, _02831_);
  or (_03212_, _03196_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_03213_, _03212_, _03211_);
  and (_03214_, _03213_, _03203_);
  and (_03215_, _03209_, _02904_);
  or (_12672_[2], _03215_, _03214_);
  or (_03216_, _03204_, _02906_);
  or (_03217_, _03196_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_03218_, _03217_, _03216_);
  and (_03219_, _03218_, _03203_);
  and (_03220_, _03209_, _02911_);
  or (_12672_[3], _03220_, _03219_);
  or (_03221_, _03204_, _02913_);
  or (_03222_, _03196_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_03223_, _03222_, _03221_);
  and (_03224_, _03223_, _03203_);
  and (_03225_, _03209_, _02919_);
  or (_12672_[4], _03225_, _03224_);
  or (_03226_, _03204_, _02921_);
  or (_03227_, _03196_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_03228_, _03227_, _03226_);
  and (_03229_, _03228_, _03203_);
  and (_03230_, _03209_, _02850_);
  or (_12672_[5], _03230_, _03229_);
  or (_03231_, _03204_, _02927_);
  or (_03232_, _03196_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_03233_, _03232_, _03231_);
  and (_03234_, _03233_, _03203_);
  and (_03235_, _03209_, _02932_);
  or (_12672_[6], _03235_, _03234_);
  or (_03236_, _03204_, _02658_);
  or (_03237_, _03196_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_03238_, _03237_, _03236_);
  and (_03239_, _03238_, _03203_);
  and (_03240_, _03209_, _02670_);
  or (_12672_[7], _03240_, _03239_);
  not (_03241_, \oc8051_golden_model_1.IRAM[8] [0]);
  not (_03242_, WR_ADDR_ABSTR_IRAM_0[2]);
  and (_03243_, _02811_, _03242_);
  and (_03244_, _03243_, _02814_);
  nor (_03245_, _03244_, _03241_);
  and (_03246_, _03244_, _02867_);
  nor (_03247_, _03246_, _03245_);
  not (_03248_, WR_ADDR_ABSTR_IRAM_1[2]);
  and (_03249_, _02805_, _03248_);
  and (_03250_, _03249_, _02804_);
  nor (_03251_, _03250_, _03247_);
  and (_03252_, _03250_, _02874_);
  or (_12673_[0], _03252_, _03251_);
  or (_03253_, _03057_, _02879_);
  or (_03254_, _03253_, _03056_);
  not (_03255_, _03244_);
  or (_03256_, _03255_, _02824_);
  or (_03257_, _03244_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_03258_, _03257_, _03256_);
  and (_03259_, _03258_, _03254_);
  and (_03260_, _03250_, _02898_);
  or (_12673_[1], _03260_, _03259_);
  or (_03261_, _03255_, _02831_);
  or (_03262_, _03244_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_03263_, _03262_, _03261_);
  and (_03264_, _03263_, _03254_);
  and (_03265_, _03250_, _02904_);
  or (_12673_[2], _03265_, _03264_);
  or (_03266_, _03255_, _02906_);
  or (_03267_, _03244_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_03268_, _03267_, _03266_);
  and (_03269_, _03268_, _03254_);
  and (_03270_, _03250_, _02911_);
  or (_12673_[3], _03270_, _03269_);
  or (_03271_, _03255_, _02913_);
  or (_03272_, _03244_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_03273_, _03272_, _03271_);
  and (_03274_, _03273_, _03254_);
  and (_03275_, _03250_, _02919_);
  or (_12673_[4], _03275_, _03274_);
  or (_03277_, _03255_, _02921_);
  or (_03278_, _03244_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_03279_, _03278_, _03277_);
  and (_03280_, _03279_, _03254_);
  and (_03281_, _03250_, _02850_);
  or (_12673_[5], _03281_, _03280_);
  or (_03282_, _03255_, _02927_);
  or (_03283_, _03244_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_03284_, _03283_, _03282_);
  and (_03285_, _03284_, _03254_);
  and (_03286_, _03250_, _02932_);
  or (_12673_[6], _03286_, _03285_);
  or (_03287_, _03255_, _02658_);
  or (_03288_, _03244_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_03289_, _03288_, _03287_);
  and (_03290_, _03289_, _03254_);
  and (_03291_, _03250_, _02670_);
  or (_12673_[7], _03291_, _03290_);
  not (_03292_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03293_, _03243_, _02864_);
  nor (_03294_, _03293_, _03292_);
  and (_03295_, _03293_, _02867_);
  or (_03296_, _03295_, _03294_);
  and (_03297_, _03249_, _02871_);
  not (_03298_, _03297_);
  and (_03299_, _03298_, _03296_);
  and (_03300_, _03297_, _02874_);
  or (_12674_[0], _03300_, _03299_);
  not (_03301_, _03293_);
  or (_03302_, _03301_, _02824_);
  or (_03303_, _03293_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03304_, _03303_, _03298_);
  and (_03305_, _03304_, _03302_);
  and (_03306_, _03297_, _02898_);
  or (_12674_[1], _03306_, _03305_);
  not (_03307_, \oc8051_golden_model_1.IRAM[9] [2]);
  nor (_03308_, _03293_, _03307_);
  and (_03309_, _03293_, _02831_);
  or (_03310_, _03309_, _03308_);
  and (_03311_, _03310_, _03298_);
  and (_03312_, _03297_, _02904_);
  or (_12674_[2], _03312_, _03311_);
  or (_03313_, _03301_, _02906_);
  or (_03314_, _03293_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_03315_, _03314_, _03298_);
  and (_03316_, _03315_, _03313_);
  and (_03317_, _03297_, _02911_);
  or (_12674_[3], _03317_, _03316_);
  not (_03318_, \oc8051_golden_model_1.IRAM[9] [4]);
  nor (_03319_, _03293_, _03318_);
  and (_03320_, _03293_, _02913_);
  or (_03321_, _03320_, _03319_);
  and (_03322_, _03321_, _03298_);
  and (_03323_, _03297_, _02919_);
  or (_12674_[4], _03323_, _03322_);
  not (_03324_, \oc8051_golden_model_1.IRAM[9] [5]);
  nor (_03325_, _03293_, _03324_);
  and (_03326_, _03293_, _02921_);
  or (_03327_, _03326_, _03325_);
  and (_03328_, _03327_, _03298_);
  and (_03329_, _03297_, _02850_);
  or (_12674_[5], _03329_, _03328_);
  not (_03330_, \oc8051_golden_model_1.IRAM[9] [6]);
  nor (_03331_, _03293_, _03330_);
  and (_03332_, _03293_, _02927_);
  or (_03333_, _03332_, _03331_);
  and (_03334_, _03333_, _03298_);
  and (_03335_, _03297_, _02932_);
  or (_12674_[6], _03335_, _03334_);
  or (_03336_, _03301_, _02658_);
  or (_03337_, _03293_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_03338_, _03337_, _03298_);
  and (_03339_, _03338_, _03336_);
  and (_03340_, _03297_, _02670_);
  or (_12674_[7], _03340_, _03339_);
  not (_03341_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_03342_, _03243_, _02941_);
  nor (_03343_, _03342_, _03341_);
  and (_03344_, _03342_, _02867_);
  nor (_03345_, _03344_, _03343_);
  and (_03346_, _03249_, _02947_);
  nor (_03347_, _03346_, _03345_);
  and (_03348_, _03346_, _02874_);
  or (_12662_[0], _03348_, _03347_);
  or (_03349_, _03253_, _02951_);
  not (_03350_, _03342_);
  or (_03351_, _03350_, _02824_);
  or (_03352_, _03342_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03353_, _03352_, _03351_);
  and (_03354_, _03353_, _03349_);
  and (_03355_, _03346_, _02898_);
  or (_12662_[1], _03355_, _03354_);
  or (_03356_, _03350_, _02831_);
  or (_03357_, _03342_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_03358_, _03357_, _03356_);
  and (_03359_, _03358_, _03349_);
  and (_03360_, _03346_, _02904_);
  or (_12662_[2], _03360_, _03359_);
  or (_03361_, _03350_, _02906_);
  or (_03362_, _03342_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_03363_, _03362_, _03361_);
  and (_03364_, _03363_, _03349_);
  and (_03365_, _03346_, _02911_);
  or (_12662_[3], _03365_, _03364_);
  or (_03366_, _03350_, _02913_);
  or (_03367_, _03342_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_03368_, _03367_, _03366_);
  and (_03369_, _03368_, _03349_);
  and (_03370_, _03346_, _02919_);
  or (_12662_[4], _03370_, _03369_);
  or (_03371_, _03350_, _02921_);
  or (_03372_, _03342_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_03373_, _03372_, _03371_);
  and (_03374_, _03373_, _03349_);
  and (_03375_, _03346_, _02850_);
  or (_12662_[5], _03375_, _03374_);
  or (_03376_, _03350_, _02927_);
  or (_03377_, _03342_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_03378_, _03377_, _03376_);
  and (_03379_, _03378_, _03349_);
  and (_03380_, _03346_, _02932_);
  or (_12662_[6], _03380_, _03379_);
  or (_03381_, _03350_, _02658_);
  or (_03382_, _03342_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_03383_, _03382_, _03381_);
  and (_03384_, _03383_, _03349_);
  and (_03385_, _03346_, _02670_);
  or (_12662_[7], _03385_, _03384_);
  not (_03386_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_03387_, _03243_, _02655_);
  nor (_03388_, _03387_, _03386_);
  and (_03389_, _03387_, _02867_);
  or (_03390_, _03389_, _03388_);
  and (_03391_, _03249_, _02664_);
  not (_03392_, _03391_);
  and (_03393_, _03392_, _03390_);
  and (_03394_, _03391_, _02874_);
  or (_12663_[0], _03394_, _03393_);
  not (_03395_, _03387_);
  or (_03396_, _03395_, _02824_);
  or (_03397_, _03387_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_03398_, _03397_, _03396_);
  or (_03399_, _03398_, _03391_);
  or (_03400_, _03392_, _02898_);
  and (_12663_[1], _03400_, _03399_);
  not (_03401_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor (_03402_, _03387_, _03401_);
  and (_03403_, _03387_, _02831_);
  or (_03404_, _03403_, _03402_);
  and (_03405_, _03404_, _03392_);
  and (_03406_, _03391_, _02904_);
  or (_12663_[2], _03406_, _03405_);
  not (_03407_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor (_03408_, _03387_, _03407_);
  and (_03409_, _03387_, _02906_);
  or (_03410_, _03409_, _03408_);
  and (_03411_, _03410_, _03392_);
  and (_03412_, _03391_, _02911_);
  or (_12663_[3], _03412_, _03411_);
  and (_03413_, _03395_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_03414_, _03387_, _02913_);
  or (_03415_, _03414_, _03413_);
  and (_03416_, _03415_, _03392_);
  and (_03417_, _03391_, _02919_);
  or (_12663_[4], _03417_, _03416_);
  or (_03418_, _03395_, _02921_);
  or (_03419_, _03387_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_03420_, _03419_, _03418_);
  or (_03421_, _03420_, _03391_);
  or (_03422_, _03392_, _02850_);
  and (_12663_[5], _03422_, _03421_);
  and (_03423_, _03395_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_03424_, _03387_, _02927_);
  or (_03425_, _03424_, _03423_);
  and (_03426_, _03425_, _03392_);
  and (_03427_, _03391_, _02932_);
  or (_12663_[6], _03427_, _03426_);
  nor (_03428_, _03387_, _02774_);
  and (_03429_, _03387_, _02658_);
  or (_03430_, _03429_, _03428_);
  and (_03431_, _03430_, _03392_);
  and (_03432_, _03391_, _02670_);
  or (_12663_[7], _03432_, _03431_);
  not (_03433_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_03434_, _02814_, _02653_);
  nor (_03435_, _03434_, _03433_);
  and (_03436_, _03434_, _02867_);
  nor (_03437_, _03436_, _03435_);
  and (_03438_, _02804_, _02666_);
  nor (_03439_, _03438_, _03437_);
  and (_03440_, _03438_, _02874_);
  or (_12664_[0], _03440_, _03439_);
  not (_03441_, _03434_);
  nor (_03442_, _03441_, _02824_);
  and (_03443_, _02805_, WR_ADDR_ABSTR_IRAM_1[2]);
  and (_03444_, _02804_, _03443_);
  nor (_03445_, _03434_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_03446_, _03445_, _03444_);
  nor (_03447_, _03446_, _03442_);
  and (_03448_, _03444_, _02898_);
  or (_12664_[1], _03448_, _03447_);
  or (_03450_, _03441_, _02831_);
  nor (_03451_, _03434_, \oc8051_golden_model_1.IRAM[12] [2]);
  nor (_03452_, _03451_, _03444_);
  and (_03453_, _03452_, _03450_);
  and (_03454_, _03444_, _02904_);
  or (_12664_[2], _03454_, _03453_);
  nor (_03455_, _03441_, _02906_);
  nor (_03456_, _03434_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_03457_, _03456_, _03444_);
  nor (_03458_, _03457_, _03455_);
  and (_03459_, _03444_, _02911_);
  or (_12664_[3], _03459_, _03458_);
  nor (_03460_, _03441_, _02913_);
  nor (_03461_, _03434_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_03462_, _03461_, _03444_);
  nor (_03463_, _03462_, _03460_);
  and (_03464_, _03444_, _02919_);
  or (_12664_[4], _03464_, _03463_);
  or (_03465_, _03441_, _02921_);
  nor (_03466_, _03434_, \oc8051_golden_model_1.IRAM[12] [5]);
  nor (_03467_, _03466_, _03444_);
  and (_03468_, _03467_, _03465_);
  and (_03469_, _03444_, _02850_);
  or (_12664_[5], _03469_, _03468_);
  nor (_03470_, _03441_, _02927_);
  nor (_03471_, _03434_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_03472_, _03471_, _03444_);
  nor (_03473_, _03472_, _03470_);
  and (_03474_, _03444_, _02932_);
  or (_12664_[6], _03474_, _03473_);
  nor (_03475_, _03441_, _02658_);
  nor (_03476_, _03434_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_03477_, _03476_, _03444_);
  nor (_03478_, _03477_, _03475_);
  and (_03479_, _03444_, _02670_);
  or (_12664_[7], _03479_, _03478_);
  and (_03480_, _02864_, _02653_);
  not (_03481_, _03480_);
  or (_03482_, _03481_, _02867_);
  and (_03483_, _02871_, _03443_);
  nor (_03484_, _03480_, \oc8051_golden_model_1.IRAM[13] [0]);
  nor (_03485_, _03484_, _03483_);
  and (_03486_, _03485_, _03482_);
  and (_03487_, _02871_, _02666_);
  and (_03488_, _03487_, _02874_);
  or (_12665_[0], _03488_, _03486_);
  nor (_03489_, _03481_, _02824_);
  nor (_03490_, _03480_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_03491_, _03490_, _03483_);
  nor (_03492_, _03491_, _03489_);
  and (_03493_, _03483_, _02898_);
  or (_12665_[1], _03493_, _03492_);
  nor (_03494_, _03481_, _02831_);
  nor (_03495_, _03480_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_03496_, _03495_, _03483_);
  nor (_03497_, _03496_, _03494_);
  and (_03498_, _03483_, _02904_);
  or (_12665_[2], _03498_, _03497_);
  nor (_03499_, _03481_, _02906_);
  nor (_03500_, _03480_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_03501_, _03500_, _03483_);
  nor (_03502_, _03501_, _03499_);
  and (_03503_, _03483_, _02911_);
  or (_12665_[3], _03503_, _03502_);
  nor (_03504_, _03481_, _02913_);
  nor (_03505_, _03480_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_03506_, _03505_, _03483_);
  nor (_03507_, _03506_, _03504_);
  and (_03508_, _03483_, _02919_);
  or (_12665_[4], _03508_, _03507_);
  not (_03509_, \oc8051_golden_model_1.IRAM[13] [5]);
  nor (_03510_, _03480_, _03509_);
  and (_03511_, _03480_, _02921_);
  nor (_03512_, _03511_, _03510_);
  nor (_03513_, _03512_, _03487_);
  and (_03514_, _03487_, _02850_);
  or (_12665_[5], _03514_, _03513_);
  nor (_03515_, _03481_, _02927_);
  nor (_03516_, _03480_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_03517_, _03516_, _03483_);
  nor (_03518_, _03517_, _03515_);
  and (_03519_, _03483_, _02932_);
  or (_12665_[6], _03519_, _03518_);
  or (_03520_, _03481_, _02658_);
  nor (_03521_, _03480_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor (_03522_, _03521_, _03483_);
  and (_03523_, _03522_, _03520_);
  and (_03524_, _03487_, _02670_);
  or (_12665_[7], _03524_, _03523_);
  not (_03525_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03526_, _02941_, _02653_);
  nor (_03527_, _03526_, _03525_);
  and (_03528_, _03526_, _02867_);
  or (_03529_, _03528_, _03527_);
  and (_03530_, _02947_, _02666_);
  not (_03531_, _03530_);
  and (_03532_, _03531_, _03529_);
  and (_03533_, _03530_, _02874_);
  or (_12666_[0], _03533_, _03532_);
  not (_03534_, _03526_);
  nor (_03535_, _03534_, _02824_);
  and (_03536_, _02947_, _03443_);
  nor (_03537_, _03526_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_03538_, _03537_, _03536_);
  nor (_03539_, _03538_, _03535_);
  and (_03540_, _03536_, _02898_);
  or (_12666_[1], _03540_, _03539_);
  nor (_03541_, _03534_, _02831_);
  nor (_03542_, _03526_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_03543_, _03542_, _03536_);
  nor (_03544_, _03543_, _03541_);
  and (_03545_, _03536_, _02904_);
  or (_12666_[2], _03545_, _03544_);
  nor (_03546_, _03534_, _02906_);
  nor (_03547_, _03526_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_03548_, _03547_, _03536_);
  nor (_03549_, _03548_, _03546_);
  and (_03550_, _03536_, _02911_);
  or (_12666_[3], _03550_, _03549_);
  nor (_03551_, _03534_, _02913_);
  nor (_03552_, _03526_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_03553_, _03552_, _03536_);
  nor (_03554_, _03553_, _03551_);
  and (_03555_, _03536_, _02919_);
  or (_12666_[4], _03555_, _03554_);
  nor (_03556_, _03534_, _02921_);
  nor (_03557_, _03526_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_03558_, _03557_, _03536_);
  nor (_03559_, _03558_, _03556_);
  and (_03560_, _03536_, _02850_);
  or (_12666_[5], _03560_, _03559_);
  nor (_03561_, _03534_, _02927_);
  nor (_03562_, _03526_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_03563_, _03562_, _03536_);
  nor (_03564_, _03563_, _03561_);
  and (_03565_, _03536_, _02932_);
  or (_12666_[6], _03565_, _03564_);
  not (_03566_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_03567_, _03526_, _03566_);
  and (_03568_, _03526_, _02658_);
  or (_03569_, _03568_, _03567_);
  and (_03570_, _03569_, _03531_);
  and (_03571_, _03530_, _02670_);
  or (_12666_[7], _03571_, _03570_);
  nand (_03572_, _02882_, _02879_);
  or (_03573_, _03572_, _03000_);
  not (_03574_, _02656_);
  or (_03575_, _02867_, _03574_);
  or (_03576_, _02656_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_03577_, _03576_, _03575_);
  and (_03578_, _03577_, _03573_);
  and (_03579_, _03443_, _03007_);
  and (_03580_, _02874_, _03579_);
  or (_12667_[0], _03580_, _03578_);
  or (_03581_, _02824_, _03574_);
  or (_03582_, _02656_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_03583_, _03582_, _03581_);
  and (_03584_, _03583_, _03573_);
  and (_03585_, _02898_, _03579_);
  or (_12667_[1], _03585_, _03584_);
  not (_03586_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor (_03587_, _02656_, _03586_);
  and (_03588_, _02831_, _02656_);
  or (_03589_, _03588_, _03587_);
  and (_03590_, _03589_, _02668_);
  and (_03591_, _02904_, _02667_);
  or (_12667_[2], _03591_, _03590_);
  or (_03592_, _02906_, _03574_);
  or (_03593_, _02656_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_03594_, _03593_, _03592_);
  and (_03595_, _03594_, _03573_);
  and (_03596_, _02911_, _03579_);
  or (_12667_[3], _03596_, _03595_);
  or (_03597_, _02913_, _03574_);
  or (_03598_, _02656_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_03599_, _03598_, _03597_);
  and (_03600_, _03599_, _03573_);
  and (_03601_, _02919_, _03579_);
  or (_12667_[4], _03601_, _03600_);
  or (_03602_, _02921_, _03574_);
  or (_03603_, _02656_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_03604_, _03603_, _03602_);
  and (_03605_, _03604_, _03573_);
  and (_03606_, _02850_, _03579_);
  or (_12667_[5], _03606_, _03605_);
  not (_03607_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_03608_, _02656_, _03607_);
  and (_03609_, _02927_, _02656_);
  or (_03610_, _03609_, _03608_);
  and (_03611_, _03610_, _02668_);
  and (_03612_, _02932_, _02667_);
  or (_12667_[6], _03612_, _03611_);
  and (_03613_, _02701_, B_abstr[0]);
  not (_03614_, _02701_);
  and (_03615_, _03614_, \oc8051_golden_model_1.B [0]);
  or (_03616_, _03615_, _03613_);
  and (_12613_[0], _03616_, _12493_);
  and (_03617_, _02701_, B_abstr[1]);
  and (_03618_, _03614_, \oc8051_golden_model_1.B [1]);
  or (_03620_, _03618_, _03617_);
  and (_12613_[1], _03620_, _12493_);
  and (_03621_, _02701_, B_abstr[2]);
  not (_03622_, \oc8051_golden_model_1.B [2]);
  nor (_03623_, _02701_, _03622_);
  or (_03624_, _03623_, _03621_);
  and (_12613_[2], _03624_, _12493_);
  and (_03625_, _02701_, B_abstr[3]);
  and (_03626_, _03614_, \oc8051_golden_model_1.B [3]);
  or (_03627_, _03626_, _03625_);
  and (_12613_[3], _03627_, _12493_);
  and (_03628_, _02701_, B_abstr[4]);
  and (_03629_, _03614_, \oc8051_golden_model_1.B [4]);
  or (_03630_, _03629_, _03628_);
  and (_12613_[4], _03630_, _12493_);
  and (_03631_, _02701_, B_abstr[5]);
  and (_03632_, _03614_, \oc8051_golden_model_1.B [5]);
  or (_03633_, _03632_, _03631_);
  and (_12613_[5], _03633_, _12493_);
  and (_03634_, _02701_, B_abstr[6]);
  and (_03635_, _03614_, \oc8051_golden_model_1.B [6]);
  or (_03636_, _03635_, _03634_);
  and (_12613_[6], _03636_, _12493_);
  and (_03637_, _02738_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_03638_, _02738_, _02862_);
  nor (_03639_, _03638_, _03637_);
  nor (_03640_, _03639_, _02741_);
  and (_03641_, _02738_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor (_03642_, _02738_, _02991_);
  or (_03643_, _03642_, _03641_);
  and (_03644_, _03643_, _02741_);
  nor (_03645_, _03644_, _03640_);
  nor (_03646_, _03645_, _02737_);
  and (_03647_, _02738_, \oc8051_golden_model_1.IRAM[4] [0]);
  nor (_03648_, _02738_, _03100_);
  nor (_03649_, _03648_, _03647_);
  nor (_03650_, _03649_, _02741_);
  and (_03651_, _02738_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor (_03652_, _02738_, _03195_);
  or (_03653_, _03652_, _03651_);
  and (_03654_, _03653_, _02741_);
  nor (_03655_, _03654_, _03650_);
  nor (_03656_, _03655_, _02754_);
  or (_03657_, _03656_, _03646_);
  and (_03658_, _03657_, _02753_);
  and (_03659_, _02738_, \oc8051_golden_model_1.IRAM[8] [0]);
  nor (_03660_, _02738_, _03292_);
  nor (_03661_, _03660_, _03659_);
  nor (_03662_, _03661_, _02741_);
  and (_03663_, _02738_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor (_03664_, _02738_, _03386_);
  or (_03665_, _03664_, _03663_);
  and (_03666_, _03665_, _02741_);
  nor (_03667_, _03666_, _03662_);
  nor (_03668_, _03667_, _02737_);
  not (_03669_, _02741_);
  and (_03670_, _02738_, _03433_);
  nor (_03671_, _02738_, \oc8051_golden_model_1.IRAM[13] [0]);
  nor (_03672_, _03671_, _03670_);
  and (_03673_, _03672_, _03669_);
  and (_03674_, _02738_, \oc8051_golden_model_1.IRAM[14] [0]);
  not (_03675_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor (_03676_, _02738_, _03675_);
  or (_03677_, _03676_, _03674_);
  and (_03678_, _03677_, _02741_);
  nor (_03679_, _03678_, _03673_);
  nor (_03680_, _03679_, _02754_);
  or (_03681_, _03680_, _03668_);
  and (_03682_, _03681_, _02768_);
  or (_03683_, _03682_, _03658_);
  nor (_03684_, _03683_, \oc8051_golden_model_1.ACC [0]);
  not (_03685_, _03684_);
  and (_03686_, _02649_, _11609_);
  and (_03687_, _03686_, _03685_);
  and (_03688_, _11613_, \oc8051_golden_model_1.ACC [0]);
  and (_03689_, _02701_, ACC_abstr[0]);
  or (_03690_, _03689_, _03688_);
  or (_03691_, _03690_, _03687_);
  and (_12612_[0], _03691_, _12493_);
  nand (_03692_, _02738_, _02822_);
  nor (_03693_, _02738_, \oc8051_golden_model_1.IRAM[1] [1]);
  nor (_03694_, _03693_, _02741_);
  and (_03695_, _03694_, _03692_);
  and (_03696_, _02738_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_03697_, _02739_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03698_, _03697_, _03696_);
  and (_03699_, _03698_, _02741_);
  nor (_03700_, _03699_, _03695_);
  nor (_03701_, _03700_, _02737_);
  not (_03702_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand (_03703_, _02738_, _03702_);
  nor (_03704_, _02738_, \oc8051_golden_model_1.IRAM[5] [1]);
  nor (_03705_, _03704_, _02741_);
  and (_03706_, _03705_, _03703_);
  and (_03707_, _02738_, \oc8051_golden_model_1.IRAM[6] [1]);
  not (_03708_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor (_03709_, _02738_, _03708_);
  or (_03710_, _03709_, _03707_);
  and (_03711_, _03710_, _02741_);
  nor (_03712_, _03711_, _03706_);
  nor (_03713_, _03712_, _02754_);
  or (_03714_, _03713_, _03701_);
  and (_03715_, _03714_, _02753_);
  or (_03716_, _02739_, \oc8051_golden_model_1.IRAM[8] [1]);
  nor (_03717_, _02738_, \oc8051_golden_model_1.IRAM[9] [1]);
  nor (_03718_, _03717_, _02741_);
  and (_03719_, _03718_, _03716_);
  and (_03720_, _02738_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03721_, _02739_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_03722_, _03721_, _03720_);
  and (_03723_, _03722_, _02741_);
  nor (_03724_, _03723_, _03719_);
  nor (_03725_, _03724_, _02737_);
  not (_03726_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_03727_, _02738_, _03726_);
  nor (_03728_, _02738_, \oc8051_golden_model_1.IRAM[13] [1]);
  nor (_03729_, _03728_, _03727_);
  and (_03730_, _03729_, _03669_);
  and (_03731_, _02738_, \oc8051_golden_model_1.IRAM[14] [1]);
  not (_03732_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor (_03733_, _02738_, _03732_);
  or (_03734_, _03733_, _03731_);
  and (_03735_, _03734_, _02741_);
  nor (_03736_, _03735_, _03730_);
  nor (_03737_, _03736_, _02754_);
  or (_03738_, _03737_, _03725_);
  and (_03739_, _03738_, _02768_);
  or (_03740_, _03739_, _03715_);
  nor (_03741_, _03740_, \oc8051_golden_model_1.ACC [1]);
  not (_03742_, _03741_);
  and (_03743_, _03742_, _03686_);
  and (_03744_, _11613_, \oc8051_golden_model_1.ACC [1]);
  and (_03745_, _02701_, ACC_abstr[1]);
  or (_03746_, _03745_, _03744_);
  or (_03747_, _03746_, _03743_);
  and (_12612_[1], _03747_, _12493_);
  or (_03748_, _02739_, \oc8051_golden_model_1.IRAM[0] [2]);
  nor (_03749_, _02738_, \oc8051_golden_model_1.IRAM[1] [2]);
  nor (_03750_, _03749_, _02741_);
  and (_03751_, _03750_, _03748_);
  and (_03752_, _02738_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_03753_, _02739_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_03754_, _03753_, _03752_);
  and (_03755_, _03754_, _02741_);
  nor (_03756_, _03755_, _03751_);
  nand (_03757_, _03756_, _02754_);
  or (_03758_, _02739_, \oc8051_golden_model_1.IRAM[4] [2]);
  nor (_03759_, _02738_, \oc8051_golden_model_1.IRAM[5] [2]);
  nor (_03760_, _03759_, _02741_);
  and (_03761_, _03760_, _03758_);
  and (_03762_, _02738_, \oc8051_golden_model_1.IRAM[6] [2]);
  not (_03763_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor (_03764_, _02738_, _03763_);
  or (_03765_, _03764_, _03762_);
  and (_03766_, _03765_, _02741_);
  nor (_03767_, _03766_, _03761_);
  nand (_03768_, _03767_, _02737_);
  and (_03769_, _03768_, _02753_);
  and (_03770_, _03769_, _03757_);
  and (_03771_, _02738_, \oc8051_golden_model_1.IRAM[8] [2]);
  nor (_03772_, _02738_, _03307_);
  nor (_03773_, _03772_, _03771_);
  nor (_03774_, _03773_, _02741_);
  and (_03775_, _02738_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor (_03776_, _02738_, _03401_);
  or (_03777_, _03776_, _03775_);
  and (_03778_, _03777_, _02741_);
  nor (_03779_, _03778_, _03774_);
  nor (_03780_, _03779_, _02737_);
  nor (_03781_, _02739_, \oc8051_golden_model_1.IRAM[12] [2]);
  nor (_03782_, _02738_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_03783_, _03782_, _02741_);
  nor (_03784_, _03783_, _03781_);
  and (_03785_, _02738_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor (_03786_, _02738_, _03586_);
  or (_03787_, _03786_, _03785_);
  and (_03788_, _03787_, _02741_);
  nor (_03789_, _03788_, _03784_);
  nor (_03790_, _03789_, _02754_);
  or (_03791_, _03790_, _03780_);
  and (_03792_, _03791_, _02768_);
  or (_03793_, _03792_, _03770_);
  nor (_03794_, _03793_, \oc8051_golden_model_1.ACC [2]);
  not (_03795_, _03794_);
  and (_03796_, _03795_, _03686_);
  not (_03797_, \oc8051_golden_model_1.ACC [2]);
  nor (_03798_, _11609_, _03797_);
  and (_03799_, _02701_, ACC_abstr[2]);
  or (_03800_, _03799_, _03798_);
  or (_03801_, _03800_, _03796_);
  and (_12612_[2], _03801_, _12493_);
  or (_03802_, _02739_, \oc8051_golden_model_1.IRAM[0] [3]);
  nor (_03803_, _02738_, \oc8051_golden_model_1.IRAM[1] [3]);
  nor (_03804_, _03803_, _02741_);
  and (_03805_, _03804_, _03802_);
  and (_03806_, _02738_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_03807_, _02739_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_03808_, _03807_, _03806_);
  and (_03809_, _03808_, _02741_);
  nor (_03810_, _03809_, _03805_);
  nor (_03812_, _03810_, _02737_);
  and (_03813_, _02738_, \oc8051_golden_model_1.IRAM[4] [3]);
  not (_03814_, \oc8051_golden_model_1.IRAM[5] [3]);
  nor (_03815_, _02738_, _03814_);
  nor (_03816_, _03815_, _03813_);
  nor (_03817_, _03816_, _02741_);
  and (_03818_, _02738_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_03819_, _02739_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_03820_, _03819_, _03818_);
  and (_03821_, _03820_, _02741_);
  nor (_03822_, _03821_, _03817_);
  nor (_03823_, _03822_, _02754_);
  or (_03824_, _03823_, _03812_);
  and (_03825_, _03824_, _02753_);
  not (_03826_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_03827_, _02738_, _03826_);
  nor (_03828_, _02738_, \oc8051_golden_model_1.IRAM[13] [3]);
  nor (_03829_, _03828_, _03827_);
  and (_03830_, _03829_, _03669_);
  and (_03831_, _02738_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_03832_, _02739_, \oc8051_golden_model_1.IRAM[15] [3]);
  or (_03833_, _03832_, _03831_);
  and (_03834_, _03833_, _02741_);
  nor (_03835_, _03834_, _03830_);
  nand (_03836_, _03835_, _02737_);
  or (_03837_, _02739_, \oc8051_golden_model_1.IRAM[8] [3]);
  nor (_03838_, _02738_, \oc8051_golden_model_1.IRAM[9] [3]);
  nor (_03839_, _03838_, _02741_);
  and (_03840_, _03839_, _03837_);
  and (_03841_, _02738_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor (_03842_, _02738_, _03407_);
  or (_03843_, _03842_, _03841_);
  and (_03844_, _03843_, _02741_);
  nor (_03845_, _03844_, _03840_);
  nand (_03846_, _03845_, _02754_);
  and (_03847_, _03846_, _02768_);
  and (_03848_, _03847_, _03836_);
  or (_03849_, _03848_, _03825_);
  nor (_03850_, _03849_, \oc8051_golden_model_1.ACC [3]);
  not (_03851_, _03850_);
  and (_03852_, _03851_, _03686_);
  and (_03853_, _11613_, \oc8051_golden_model_1.ACC [3]);
  and (_03854_, _02701_, ACC_abstr[3]);
  or (_03855_, _03854_, _03853_);
  or (_03856_, _03855_, _03852_);
  and (_12612_[3], _03856_, _12493_);
  and (_03857_, _02738_, \oc8051_golden_model_1.IRAM[0] [4]);
  not (_03858_, \oc8051_golden_model_1.IRAM[1] [4]);
  nor (_03859_, _02738_, _03858_);
  nor (_03860_, _03859_, _03857_);
  nor (_03861_, _03860_, _02741_);
  and (_03862_, _02738_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_03863_, _02739_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_03864_, _03863_, _03862_);
  and (_03865_, _03864_, _02741_);
  nor (_03866_, _03865_, _03861_);
  nor (_03867_, _03866_, _02737_);
  and (_03868_, _02738_, \oc8051_golden_model_1.IRAM[4] [4]);
  nor (_03869_, _02738_, _03128_);
  nor (_03870_, _03869_, _03868_);
  nor (_03871_, _03870_, _02741_);
  and (_03872_, _02738_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_03873_, _02739_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_03874_, _03873_, _03872_);
  and (_03875_, _03874_, _02741_);
  nor (_03876_, _03875_, _03871_);
  nor (_03877_, _03876_, _02754_);
  or (_03878_, _03877_, _03867_);
  and (_03879_, _03878_, _02753_);
  nor (_03880_, _02738_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor (_03881_, RD_IRAM_0_ABSTR_ADDR[0], \oc8051_golden_model_1.IRAM[14] [4]);
  nor (_03882_, _03881_, _03880_);
  or (_03883_, _03882_, _02754_);
  nor (_03884_, _02738_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor (_03885_, RD_IRAM_0_ABSTR_ADDR[0], \oc8051_golden_model_1.IRAM[10] [4]);
  nor (_03886_, _03885_, _03884_);
  or (_03887_, _03886_, _02737_);
  and (_03888_, _03887_, _03883_);
  or (_03889_, _03888_, _03669_);
  and (_03890_, _02738_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_03891_, \oc8051_golden_model_1.IRAM[13] [4]);
  nor (_03892_, _02738_, _03891_);
  or (_03893_, _03892_, _03890_);
  or (_03894_, _03893_, _02754_);
  and (_03895_, _02738_, \oc8051_golden_model_1.IRAM[8] [4]);
  nor (_03896_, _02738_, _03318_);
  or (_03897_, _03896_, _02737_);
  or (_03898_, _03897_, _03895_);
  and (_03899_, _03898_, _03894_);
  or (_03900_, _03899_, _02741_);
  and (_03901_, _03900_, _03889_);
  and (_03902_, _03901_, _02768_);
  or (_03903_, _03902_, _03879_);
  nor (_03904_, _03903_, \oc8051_golden_model_1.ACC [4]);
  not (_03905_, _03904_);
  and (_03906_, _03905_, _03686_);
  and (_03907_, _11613_, \oc8051_golden_model_1.ACC [4]);
  and (_03908_, _02701_, ACC_abstr[4]);
  or (_03909_, _03908_, _03907_);
  or (_03910_, _03909_, _03906_);
  and (_12612_[4], _03910_, _12493_);
  and (_03911_, _02738_, \oc8051_golden_model_1.IRAM[0] [5]);
  not (_03912_, \oc8051_golden_model_1.IRAM[1] [5]);
  nor (_03913_, _02738_, _03912_);
  nor (_03914_, _03913_, _03911_);
  nor (_03915_, _03914_, _02741_);
  and (_03916_, _02738_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_03917_, _02739_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_03918_, _03917_, _03916_);
  and (_03919_, _03918_, _02741_);
  nor (_03920_, _03919_, _03915_);
  nor (_03921_, _03920_, _02737_);
  and (_03922_, _02738_, \oc8051_golden_model_1.IRAM[4] [5]);
  not (_03923_, \oc8051_golden_model_1.IRAM[5] [5]);
  nor (_03924_, _02738_, _03923_);
  nor (_03925_, _03924_, _03922_);
  nor (_03926_, _03925_, _02741_);
  and (_03927_, _02738_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_03928_, _02739_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_03929_, _03928_, _03927_);
  and (_03930_, _03929_, _02741_);
  nor (_03931_, _03930_, _03926_);
  nor (_03932_, _03931_, _02754_);
  or (_03933_, _03932_, _03921_);
  and (_03934_, _03933_, _02753_);
  nor (_03935_, _02738_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor (_03936_, RD_IRAM_0_ABSTR_ADDR[0], \oc8051_golden_model_1.IRAM[14] [5]);
  nor (_03937_, _03936_, _03935_);
  or (_03938_, _03937_, _02754_);
  nor (_03939_, _02738_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor (_03940_, RD_IRAM_0_ABSTR_ADDR[0], \oc8051_golden_model_1.IRAM[10] [5]);
  nor (_03941_, _03940_, _03939_);
  or (_03942_, _03941_, _02737_);
  and (_03943_, _03942_, _03938_);
  or (_03944_, _03943_, _03669_);
  and (_03945_, _02738_, \oc8051_golden_model_1.IRAM[12] [5]);
  nor (_03946_, _02738_, _03509_);
  or (_03947_, _03946_, _03945_);
  or (_03948_, _03947_, _02754_);
  and (_03949_, _02738_, \oc8051_golden_model_1.IRAM[8] [5]);
  nor (_03950_, _02738_, _03324_);
  or (_03951_, _03950_, _02737_);
  or (_03952_, _03951_, _03949_);
  and (_03953_, _03952_, _03948_);
  or (_03954_, _03953_, _02741_);
  and (_03955_, _03954_, _03944_);
  and (_03956_, _03955_, _02768_);
  or (_03957_, _03956_, \oc8051_golden_model_1.ACC [5]);
  nor (_03958_, _03957_, _03934_);
  not (_03959_, _03958_);
  and (_03960_, _03959_, _03686_);
  and (_03961_, _11613_, \oc8051_golden_model_1.ACC [5]);
  and (_03962_, _02701_, ACC_abstr[5]);
  or (_03963_, _03962_, _03961_);
  or (_03964_, _03963_, _03960_);
  and (_12612_[5], _03964_, _12493_);
  or (_03965_, _02739_, \oc8051_golden_model_1.IRAM[0] [6]);
  nor (_03966_, _02738_, \oc8051_golden_model_1.IRAM[1] [6]);
  nor (_03967_, _03966_, _02741_);
  and (_03968_, _03967_, _03965_);
  and (_03969_, _02738_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_03970_, _02739_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_03971_, _03970_, _03969_);
  and (_03972_, _03971_, _02741_);
  nor (_03973_, _03972_, _03968_);
  nor (_03974_, _03973_, _02737_);
  not (_03975_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand (_03976_, _02738_, _03975_);
  nor (_03977_, _02738_, \oc8051_golden_model_1.IRAM[5] [6]);
  nor (_03978_, _03977_, _02741_);
  and (_03979_, _03978_, _03976_);
  and (_03980_, _02738_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_03981_, _02739_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_03982_, _03981_, _03980_);
  and (_03983_, _03982_, _02741_);
  nor (_03984_, _03983_, _03979_);
  nor (_03985_, _03984_, _02754_);
  or (_03986_, _03985_, _03974_);
  and (_03987_, _03986_, _02753_);
  nor (_03988_, _02738_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor (_03989_, RD_IRAM_0_ABSTR_ADDR[0], \oc8051_golden_model_1.IRAM[14] [6]);
  nor (_03990_, _03989_, _03988_);
  or (_03991_, _03990_, _02754_);
  nor (_03992_, _02738_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor (_03993_, RD_IRAM_0_ABSTR_ADDR[0], \oc8051_golden_model_1.IRAM[10] [6]);
  nor (_03994_, _03993_, _03992_);
  or (_03995_, _03994_, _02737_);
  and (_03996_, _03995_, _03991_);
  or (_03997_, _03996_, _03669_);
  not (_03998_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_03999_, _02738_, _03998_);
  nor (_04000_, _02738_, \oc8051_golden_model_1.IRAM[13] [6]);
  nor (_04001_, _04000_, _03999_);
  or (_04002_, _04001_, _02754_);
  and (_04003_, _02738_, \oc8051_golden_model_1.IRAM[8] [6]);
  nor (_04004_, _02738_, _03330_);
  or (_04005_, _04004_, _02737_);
  or (_04006_, _04005_, _04003_);
  and (_04007_, _04006_, _04002_);
  or (_04008_, _04007_, _02741_);
  and (_04010_, _04008_, _03997_);
  and (_04011_, _04010_, _02768_);
  or (_04012_, _04011_, _03987_);
  nor (_04013_, _04012_, \oc8051_golden_model_1.ACC [6]);
  not (_04014_, _04013_);
  and (_04015_, _04014_, _03686_);
  and (_04016_, _11613_, \oc8051_golden_model_1.ACC [6]);
  and (_04017_, _02701_, ACC_abstr[6]);
  or (_04018_, _04017_, _04016_);
  or (_04019_, _04018_, _04015_);
  and (_12612_[6], _04019_, _12493_);
  and (_04020_, _02701_, DPL_abstr[0]);
  and (_04021_, _03614_, \oc8051_golden_model_1.DPL [0]);
  or (_04022_, _04021_, _04020_);
  and (_12615_[0], _04022_, _12493_);
  and (_04023_, _02701_, DPL_abstr[1]);
  and (_04024_, _03614_, \oc8051_golden_model_1.DPL [1]);
  or (_04025_, _04024_, _04023_);
  and (_12615_[1], _04025_, _12493_);
  and (_04026_, _02701_, DPL_abstr[2]);
  not (_04027_, \oc8051_golden_model_1.DPL [2]);
  nor (_04028_, _02701_, _04027_);
  or (_04029_, _04028_, _04026_);
  and (_12615_[2], _04029_, _12493_);
  and (_04030_, _02701_, DPL_abstr[3]);
  and (_04031_, _03614_, \oc8051_golden_model_1.DPL [3]);
  or (_04032_, _04031_, _04030_);
  and (_12615_[3], _04032_, _12493_);
  and (_04033_, _02701_, DPL_abstr[4]);
  and (_04034_, _03614_, \oc8051_golden_model_1.DPL [4]);
  or (_04035_, _04034_, _04033_);
  and (_12615_[4], _04035_, _12493_);
  and (_04036_, _02701_, DPL_abstr[5]);
  and (_04037_, _03614_, \oc8051_golden_model_1.DPL [5]);
  or (_04038_, _04037_, _04036_);
  and (_12615_[5], _04038_, _12493_);
  and (_04039_, _02701_, DPL_abstr[6]);
  and (_04040_, _03614_, \oc8051_golden_model_1.DPL [6]);
  or (_04041_, _04040_, _04039_);
  and (_12615_[6], _04041_, _12493_);
  and (_04042_, _02701_, DPH_abstr[0]);
  and (_04043_, _03614_, \oc8051_golden_model_1.DPH [0]);
  or (_04044_, _04043_, _04042_);
  and (_12614_[0], _04044_, _12493_);
  and (_04045_, _02701_, DPH_abstr[1]);
  and (_04046_, _03614_, \oc8051_golden_model_1.DPH [1]);
  or (_04047_, _04046_, _04045_);
  and (_12614_[1], _04047_, _12493_);
  and (_04048_, _02701_, DPH_abstr[2]);
  not (_04049_, \oc8051_golden_model_1.DPH [2]);
  nor (_04050_, _02701_, _04049_);
  or (_04051_, _04050_, _04048_);
  and (_12614_[2], _04051_, _12493_);
  and (_04052_, _02701_, DPH_abstr[3]);
  and (_04053_, _03614_, \oc8051_golden_model_1.DPH [3]);
  or (_04054_, _04053_, _04052_);
  and (_12614_[3], _04054_, _12493_);
  and (_04055_, _02701_, DPH_abstr[4]);
  and (_04056_, _03614_, \oc8051_golden_model_1.DPH [4]);
  or (_04057_, _04056_, _04055_);
  and (_12614_[4], _04057_, _12493_);
  and (_04058_, _02701_, DPH_abstr[5]);
  and (_04059_, _03614_, \oc8051_golden_model_1.DPH [5]);
  or (_04060_, _04059_, _04058_);
  and (_12614_[5], _04060_, _12493_);
  and (_04061_, _02701_, DPH_abstr[6]);
  and (_04062_, _03614_, \oc8051_golden_model_1.DPH [6]);
  or (_04063_, _04062_, _04061_);
  and (_12614_[6], _04063_, _12493_);
  and (_12616_[0], \oc8051_golden_model_1.IE [0], _12493_);
  and (_12616_[1], \oc8051_golden_model_1.IE [1], _12493_);
  and (_12616_[2], \oc8051_golden_model_1.IE [2], _12493_);
  and (_12616_[3], \oc8051_golden_model_1.IE [3], _12493_);
  and (_12616_[4], \oc8051_golden_model_1.IE [4], _12493_);
  and (_12616_[5], \oc8051_golden_model_1.IE [5], _12493_);
  and (_12616_[6], \oc8051_golden_model_1.IE [6], _12493_);
  and (_12617_[0], \oc8051_golden_model_1.IP [0], _12493_);
  and (_12617_[1], \oc8051_golden_model_1.IP [1], _12493_);
  and (_12617_[2], \oc8051_golden_model_1.IP [2], _12493_);
  and (_12617_[3], \oc8051_golden_model_1.IP [3], _12493_);
  and (_12617_[4], \oc8051_golden_model_1.IP [4], _12493_);
  and (_12617_[5], \oc8051_golden_model_1.IP [5], _12493_);
  and (_12617_[6], \oc8051_golden_model_1.IP [6], _12493_);
  or (_04064_, _02701_, \oc8051_golden_model_1.P0 [0]);
  or (_04065_, _03614_, P0_abstr[0]);
  and (_04066_, _04065_, _04064_);
  or (_12618_[0], _04066_, rst);
  or (_04067_, _02701_, \oc8051_golden_model_1.P0 [1]);
  or (_04068_, _03614_, P0_abstr[1]);
  and (_04069_, _04068_, _04067_);
  or (_12618_[1], _04069_, rst);
  and (_04070_, _02701_, P0_abstr[2]);
  not (_04071_, \oc8051_golden_model_1.P0 [2]);
  nor (_04072_, _02701_, _04071_);
  or (_04073_, _04072_, rst);
  or (_12618_[2], _04073_, _04070_);
  or (_04074_, _02701_, \oc8051_golden_model_1.P0 [3]);
  or (_04075_, _03614_, P0_abstr[3]);
  and (_04076_, _04075_, _04074_);
  or (_12618_[3], _04076_, rst);
  or (_04077_, _02701_, \oc8051_golden_model_1.P0 [4]);
  or (_04078_, _03614_, P0_abstr[4]);
  and (_04079_, _04078_, _04077_);
  or (_12618_[4], _04079_, rst);
  or (_04080_, _02701_, \oc8051_golden_model_1.P0 [5]);
  or (_04081_, _03614_, P0_abstr[5]);
  and (_04082_, _04081_, _04080_);
  or (_12618_[5], _04082_, rst);
  or (_04083_, _02701_, \oc8051_golden_model_1.P0 [6]);
  or (_04084_, _03614_, P0_abstr[6]);
  and (_04085_, _04084_, _04083_);
  or (_12618_[6], _04085_, rst);
  or (_04086_, _02701_, \oc8051_golden_model_1.P1 [0]);
  or (_04087_, _03614_, P1_abstr[0]);
  and (_04088_, _04087_, _04086_);
  or (_12619_[0], _04088_, rst);
  or (_04089_, _02701_, \oc8051_golden_model_1.P1 [1]);
  or (_04090_, _03614_, P1_abstr[1]);
  and (_04091_, _04090_, _04089_);
  or (_12619_[1], _04091_, rst);
  and (_04092_, _02701_, P1_abstr[2]);
  not (_04093_, \oc8051_golden_model_1.P1 [2]);
  nor (_04094_, _02701_, _04093_);
  or (_04095_, _04094_, rst);
  or (_12619_[2], _04095_, _04092_);
  or (_04096_, _02701_, \oc8051_golden_model_1.P1 [3]);
  or (_04097_, _03614_, P1_abstr[3]);
  and (_04098_, _04097_, _04096_);
  or (_12619_[3], _04098_, rst);
  or (_04099_, _02701_, \oc8051_golden_model_1.P1 [4]);
  or (_04100_, _03614_, P1_abstr[4]);
  and (_04101_, _04100_, _04099_);
  or (_12619_[4], _04101_, rst);
  or (_04102_, _02701_, \oc8051_golden_model_1.P1 [5]);
  or (_04103_, _03614_, P1_abstr[5]);
  and (_04104_, _04103_, _04102_);
  or (_12619_[5], _04104_, rst);
  or (_04105_, _02701_, \oc8051_golden_model_1.P1 [6]);
  or (_04106_, _03614_, P1_abstr[6]);
  and (_04107_, _04106_, _04105_);
  or (_12619_[6], _04107_, rst);
  or (_04108_, _02701_, \oc8051_golden_model_1.P2 [0]);
  or (_04109_, _03614_, P2_abstr[0]);
  and (_04110_, _04109_, _04108_);
  or (_12620_[0], _04110_, rst);
  or (_04111_, _02701_, \oc8051_golden_model_1.P2 [1]);
  or (_04112_, _03614_, P2_abstr[1]);
  and (_04113_, _04112_, _04111_);
  or (_12620_[1], _04113_, rst);
  and (_04114_, _02701_, P2_abstr[2]);
  not (_04115_, \oc8051_golden_model_1.P2 [2]);
  nor (_04116_, _02701_, _04115_);
  or (_04117_, _04116_, rst);
  or (_12620_[2], _04117_, _04114_);
  or (_04118_, _02701_, \oc8051_golden_model_1.P2 [3]);
  or (_04119_, _03614_, P2_abstr[3]);
  and (_04120_, _04119_, _04118_);
  or (_12620_[3], _04120_, rst);
  or (_04121_, _02701_, \oc8051_golden_model_1.P2 [4]);
  or (_04122_, _03614_, P2_abstr[4]);
  and (_04123_, _04122_, _04121_);
  or (_12620_[4], _04123_, rst);
  or (_04124_, _02701_, \oc8051_golden_model_1.P2 [5]);
  or (_04125_, _03614_, P2_abstr[5]);
  and (_04126_, _04125_, _04124_);
  or (_12620_[5], _04126_, rst);
  or (_04127_, _02701_, \oc8051_golden_model_1.P2 [6]);
  or (_04128_, _03614_, P2_abstr[6]);
  and (_04129_, _04128_, _04127_);
  or (_12620_[6], _04129_, rst);
  or (_04130_, _02701_, \oc8051_golden_model_1.P3 [0]);
  or (_04131_, _03614_, P3_abstr[0]);
  and (_04132_, _04131_, _04130_);
  or (_12621_[0], _04132_, rst);
  or (_04133_, _02701_, \oc8051_golden_model_1.P3 [1]);
  or (_04134_, _03614_, P3_abstr[1]);
  and (_04135_, _04134_, _04133_);
  or (_12621_[1], _04135_, rst);
  and (_04136_, _02701_, P3_abstr[2]);
  not (_04137_, \oc8051_golden_model_1.P3 [2]);
  nor (_04138_, _02701_, _04137_);
  or (_04139_, _04138_, rst);
  or (_12621_[2], _04139_, _04136_);
  or (_04140_, _02701_, \oc8051_golden_model_1.P3 [3]);
  or (_04141_, _03614_, P3_abstr[3]);
  and (_04142_, _04141_, _04140_);
  or (_12621_[3], _04142_, rst);
  or (_04143_, _02701_, \oc8051_golden_model_1.P3 [4]);
  or (_04144_, _03614_, P3_abstr[4]);
  and (_04145_, _04144_, _04143_);
  or (_12621_[4], _04145_, rst);
  or (_04146_, _02701_, \oc8051_golden_model_1.P3 [5]);
  or (_04147_, _03614_, P3_abstr[5]);
  and (_04148_, _04147_, _04146_);
  or (_12621_[5], _04148_, rst);
  or (_04149_, _02701_, \oc8051_golden_model_1.P3 [6]);
  or (_04150_, _03614_, P3_abstr[6]);
  and (_04151_, _04150_, _04149_);
  or (_12621_[6], _04151_, rst);
  and (_04152_, _02672_, PSW_abstr[0]);
  nor (_04154_, _04152_, _02794_);
  and (_04155_, _03741_, _03684_);
  nor (_04156_, _03741_, _03684_);
  nor (_04157_, _04156_, _04155_);
  nor (_04158_, _04157_, _03959_);
  and (_04159_, _04157_, _03959_);
  nor (_04160_, _04159_, _04158_);
  nor (_04161_, _04013_, _03904_);
  and (_04162_, _04013_, _03904_);
  nor (_04163_, _04162_, _04161_);
  nor (_04164_, _03850_, _03795_);
  and (_04165_, _03850_, _03795_);
  nor (_04166_, _04165_, _04164_);
  nor (_04167_, _04166_, _04163_);
  and (_04168_, _04166_, _04163_);
  nor (_04169_, _04168_, _04167_);
  and (_04170_, _04169_, _04160_);
  nor (_04171_, _04169_, _04160_);
  nor (_04172_, _04171_, _04170_);
  and (_04173_, _04172_, _02649_);
  nor (_04174_, _04173_, _04154_);
  not (_04175_, _02793_);
  and (_04176_, _04173_, _04175_);
  or (_04177_, _04176_, _04174_);
  or (_04178_, _04177_, _11613_);
  or (_04179_, _11609_, \oc8051_golden_model_1.PSW [0]);
  and (_04180_, _04179_, _12493_);
  and (_12624_[0], _04180_, _04178_);
  not (_04181_, \oc8051_golden_model_1.PSW [1]);
  nor (_04182_, _02701_, _04181_);
  and (_04183_, _02701_, PSW_abstr[1]);
  or (_04184_, _04183_, _04182_);
  and (_12624_[1], _04184_, _12493_);
  and (_04185_, _03614_, \oc8051_golden_model_1.PSW [2]);
  and (_04186_, _02701_, PSW_abstr[2]);
  or (_04187_, _04186_, _04185_);
  and (_12624_[2], _04187_, _12493_);
  not (_04188_, \oc8051_golden_model_1.PSW [3]);
  nor (_04189_, _02701_, _04188_);
  and (_04190_, _02701_, PSW_abstr[3]);
  or (_04191_, _04190_, _04189_);
  and (_12624_[3], _04191_, _12493_);
  not (_04192_, \oc8051_golden_model_1.PSW [4]);
  nor (_04193_, _02701_, _04192_);
  and (_04194_, _02701_, PSW_abstr[4]);
  or (_04195_, _04194_, _04193_);
  and (_12624_[4], _04195_, _12493_);
  not (_04196_, \oc8051_golden_model_1.PSW [5]);
  nor (_04197_, _02701_, _04196_);
  and (_04198_, _02701_, PSW_abstr[5]);
  or (_04199_, _04198_, _04197_);
  and (_12624_[5], _04199_, _12493_);
  and (_04200_, _03614_, \oc8051_golden_model_1.PSW [6]);
  and (_04201_, _02701_, PSW_abstr[6]);
  or (_04202_, _04201_, _04200_);
  and (_12624_[6], _04202_, _12493_);
  and (_12622_[0], \oc8051_golden_model_1.PCON [0], _12493_);
  and (_12622_[1], \oc8051_golden_model_1.PCON [1], _12493_);
  and (_12622_[2], \oc8051_golden_model_1.PCON [2], _12493_);
  and (_12622_[3], \oc8051_golden_model_1.PCON [3], _12493_);
  and (_12622_[4], \oc8051_golden_model_1.PCON [4], _12493_);
  and (_12622_[5], \oc8051_golden_model_1.PCON [5], _12493_);
  and (_12622_[6], \oc8051_golden_model_1.PCON [6], _12493_);
  and (_12625_[0], \oc8051_golden_model_1.SBUF [0], _12493_);
  and (_12625_[1], \oc8051_golden_model_1.SBUF [1], _12493_);
  and (_12625_[2], \oc8051_golden_model_1.SBUF [2], _12493_);
  and (_12625_[3], \oc8051_golden_model_1.SBUF [3], _12493_);
  and (_12625_[4], \oc8051_golden_model_1.SBUF [4], _12493_);
  and (_12625_[5], \oc8051_golden_model_1.SBUF [5], _12493_);
  and (_12625_[6], \oc8051_golden_model_1.SBUF [6], _12493_);
  and (_12626_[0], \oc8051_golden_model_1.SCON [0], _12493_);
  and (_12626_[1], \oc8051_golden_model_1.SCON [1], _12493_);
  and (_12626_[2], \oc8051_golden_model_1.SCON [2], _12493_);
  and (_12626_[3], \oc8051_golden_model_1.SCON [3], _12493_);
  and (_12626_[4], \oc8051_golden_model_1.SCON [4], _12493_);
  and (_12626_[5], \oc8051_golden_model_1.SCON [5], _12493_);
  and (_12626_[6], \oc8051_golden_model_1.SCON [6], _12493_);
  and (_04203_, _02701_, SP_abstr[0]);
  not (_04204_, \oc8051_golden_model_1.SP [0]);
  nor (_04205_, _02701_, _04204_);
  or (_04206_, _04205_, rst);
  or (_12627_[0], _04206_, _04203_);
  and (_04207_, _02701_, SP_abstr[1]);
  and (_04208_, _03614_, \oc8051_golden_model_1.SP [1]);
  or (_04209_, _04208_, rst);
  or (_12627_[1], _04209_, _04207_);
  and (_04210_, _02701_, SP_abstr[2]);
  and (_04211_, _03614_, \oc8051_golden_model_1.SP [2]);
  or (_04212_, _04211_, rst);
  or (_12627_[2], _04212_, _04210_);
  and (_04213_, _02701_, SP_abstr[3]);
  and (_04214_, _03614_, \oc8051_golden_model_1.SP [3]);
  or (_04215_, _04214_, _04213_);
  and (_12627_[3], _04215_, _12493_);
  and (_04216_, _02701_, SP_abstr[4]);
  and (_04217_, _03614_, \oc8051_golden_model_1.SP [4]);
  or (_04218_, _04217_, _04216_);
  and (_12627_[4], _04218_, _12493_);
  and (_04219_, _02701_, SP_abstr[5]);
  and (_04220_, _03614_, \oc8051_golden_model_1.SP [5]);
  or (_04222_, _04220_, _04219_);
  and (_12627_[5], _04222_, _12493_);
  and (_04223_, _02701_, SP_abstr[6]);
  and (_04224_, _03614_, \oc8051_golden_model_1.SP [6]);
  or (_04225_, _04224_, _04223_);
  and (_12627_[6], _04225_, _12493_);
  and (_12628_[0], \oc8051_golden_model_1.TCON [0], _12493_);
  and (_12628_[1], \oc8051_golden_model_1.TCON [1], _12493_);
  and (_12628_[2], \oc8051_golden_model_1.TCON [2], _12493_);
  and (_12628_[3], \oc8051_golden_model_1.TCON [3], _12493_);
  and (_12628_[4], \oc8051_golden_model_1.TCON [4], _12493_);
  and (_12628_[5], \oc8051_golden_model_1.TCON [5], _12493_);
  and (_12628_[6], \oc8051_golden_model_1.TCON [6], _12493_);
  and (_12629_[0], \oc8051_golden_model_1.TH0 [0], _12493_);
  and (_12629_[1], \oc8051_golden_model_1.TH0 [1], _12493_);
  and (_12629_[2], \oc8051_golden_model_1.TH0 [2], _12493_);
  and (_12629_[3], \oc8051_golden_model_1.TH0 [3], _12493_);
  and (_12629_[4], \oc8051_golden_model_1.TH0 [4], _12493_);
  and (_12629_[5], \oc8051_golden_model_1.TH0 [5], _12493_);
  and (_12629_[6], \oc8051_golden_model_1.TH0 [6], _12493_);
  and (_12630_[0], \oc8051_golden_model_1.TH1 [0], _12493_);
  and (_12630_[1], \oc8051_golden_model_1.TH1 [1], _12493_);
  and (_12630_[2], \oc8051_golden_model_1.TH1 [2], _12493_);
  and (_12630_[3], \oc8051_golden_model_1.TH1 [3], _12493_);
  and (_12630_[4], \oc8051_golden_model_1.TH1 [4], _12493_);
  and (_12630_[5], \oc8051_golden_model_1.TH1 [5], _12493_);
  and (_12630_[6], \oc8051_golden_model_1.TH1 [6], _12493_);
  and (_12631_[0], \oc8051_golden_model_1.TL0 [0], _12493_);
  and (_12631_[1], \oc8051_golden_model_1.TL0 [1], _12493_);
  and (_12631_[2], \oc8051_golden_model_1.TL0 [2], _12493_);
  and (_12631_[3], \oc8051_golden_model_1.TL0 [3], _12493_);
  and (_12631_[4], \oc8051_golden_model_1.TL0 [4], _12493_);
  and (_12631_[5], \oc8051_golden_model_1.TL0 [5], _12493_);
  and (_12631_[6], \oc8051_golden_model_1.TL0 [6], _12493_);
  and (_12632_[0], \oc8051_golden_model_1.TL1 [0], _12493_);
  and (_12632_[1], \oc8051_golden_model_1.TL1 [1], _12493_);
  and (_12632_[2], \oc8051_golden_model_1.TL1 [2], _12493_);
  and (_12632_[3], \oc8051_golden_model_1.TL1 [3], _12493_);
  and (_12632_[4], \oc8051_golden_model_1.TL1 [4], _12493_);
  and (_12632_[5], \oc8051_golden_model_1.TL1 [5], _12493_);
  and (_12632_[6], \oc8051_golden_model_1.TL1 [6], _12493_);
  and (_12633_[0], \oc8051_golden_model_1.TMOD [0], _12493_);
  and (_12633_[1], \oc8051_golden_model_1.TMOD [1], _12493_);
  and (_12633_[2], \oc8051_golden_model_1.TMOD [2], _12493_);
  and (_12633_[3], \oc8051_golden_model_1.TMOD [3], _12493_);
  and (_12633_[4], \oc8051_golden_model_1.TMOD [4], _12493_);
  and (_12633_[5], \oc8051_golden_model_1.TMOD [5], _12493_);
  and (_12633_[6], \oc8051_golden_model_1.TMOD [6], _12493_);
  and (_04226_, _02672_, XRAM_ADDR_abstr[0]);
  or (_04227_, _04226_, _11613_);
  or (_04228_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [0]);
  and (_04229_, _04228_, _12493_);
  and (_12634_[0], _04229_, _04227_);
  and (_04230_, _02672_, XRAM_ADDR_abstr[1]);
  or (_04231_, _04230_, _11613_);
  or (_04232_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [1]);
  and (_04233_, _04232_, _12493_);
  and (_12634_[1], _04233_, _04231_);
  and (_04234_, _02672_, XRAM_ADDR_abstr[2]);
  or (_04235_, _04234_, _11613_);
  or (_04236_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [2]);
  and (_04237_, _04236_, _12493_);
  and (_12634_[2], _04237_, _04235_);
  and (_04238_, _02672_, XRAM_ADDR_abstr[3]);
  or (_04239_, _04238_, _11613_);
  or (_04240_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [3]);
  and (_04241_, _04240_, _12493_);
  and (_12634_[3], _04241_, _04239_);
  and (_04242_, _02672_, XRAM_ADDR_abstr[4]);
  or (_04243_, _04242_, _11613_);
  or (_04244_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [4]);
  and (_04245_, _04244_, _12493_);
  and (_12634_[4], _04245_, _04243_);
  and (_04246_, _02672_, XRAM_ADDR_abstr[5]);
  or (_04247_, _04246_, _11613_);
  or (_04248_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [5]);
  and (_04249_, _04248_, _12493_);
  and (_12634_[5], _04249_, _04247_);
  and (_04250_, _02672_, XRAM_ADDR_abstr[6]);
  or (_04251_, _04250_, _11613_);
  or (_04252_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [6]);
  and (_04253_, _04252_, _12493_);
  and (_12634_[6], _04253_, _04251_);
  and (_04254_, _02672_, XRAM_ADDR_abstr[7]);
  or (_04255_, _04254_, _11613_);
  or (_04256_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [7]);
  and (_04257_, _04256_, _12493_);
  and (_12634_[7], _04257_, _04255_);
  and (_04258_, _02672_, XRAM_ADDR_abstr[8]);
  or (_04259_, _04258_, _11613_);
  or (_04260_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [8]);
  and (_04261_, _04260_, _12493_);
  and (_12634_[8], _04261_, _04259_);
  and (_04262_, _02672_, XRAM_ADDR_abstr[9]);
  or (_04263_, _04262_, _11613_);
  or (_04264_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [9]);
  and (_04265_, _04264_, _12493_);
  and (_12634_[9], _04265_, _04263_);
  and (_04266_, _02672_, XRAM_ADDR_abstr[10]);
  or (_04267_, _04266_, _11613_);
  or (_04269_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [10]);
  and (_04270_, _04269_, _12493_);
  and (_12634_[10], _04270_, _04267_);
  and (_04271_, _02672_, XRAM_ADDR_abstr[11]);
  or (_04272_, _04271_, _11613_);
  or (_04273_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [11]);
  and (_04274_, _04273_, _12493_);
  and (_12634_[11], _04274_, _04272_);
  and (_04275_, _02672_, XRAM_ADDR_abstr[12]);
  or (_04276_, _04275_, _11613_);
  or (_04277_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [12]);
  and (_04278_, _04277_, _12493_);
  and (_12634_[12], _04278_, _04276_);
  and (_04279_, _02672_, XRAM_ADDR_abstr[13]);
  or (_04280_, _04279_, _11613_);
  or (_04281_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [13]);
  and (_04282_, _04281_, _12493_);
  and (_12634_[13], _04282_, _04280_);
  and (_04283_, _02672_, XRAM_ADDR_abstr[14]);
  or (_04284_, _04283_, _11613_);
  or (_04285_, _11609_, \oc8051_golden_model_1.XRAM_ADDR [14]);
  and (_04286_, _04285_, _12493_);
  and (_12634_[14], _04286_, _04284_);
  and (_04287_, _02649_, \oc8051_golden_model_1.PC [0]);
  nor (_04288_, _02649_, PC_abstr[0]);
  nor (_04289_, _04288_, _04287_);
  or (_04290_, _04289_, _11613_);
  or (_04291_, _11609_, \oc8051_golden_model_1.PC [0]);
  and (_04292_, _04291_, _12493_);
  and (_12623_[0], _04292_, _04290_);
  nor (_04293_, _02386_, _02365_);
  and (_04294_, _04293_, _02649_);
  and (_04295_, _02672_, PC_abstr[1]);
  nor (_04296_, _04295_, _04294_);
  nand (_04297_, _04296_, _11609_);
  or (_04298_, _11609_, \oc8051_golden_model_1.PC [1]);
  and (_04299_, _04298_, _12493_);
  and (_12623_[1], _04299_, _04297_);
  nor (_04300_, _02365_, \oc8051_golden_model_1.PC [2]);
  nor (_04301_, _04300_, _02390_);
  nor (_04302_, _04301_, _02672_);
  nor (_04303_, _02649_, PC_abstr[2]);
  nor (_04304_, _04303_, _04302_);
  or (_04305_, _04304_, _11613_);
  or (_04306_, _11609_, \oc8051_golden_model_1.PC [2]);
  and (_04307_, _04306_, _12493_);
  and (_12623_[2], _04307_, _04305_);
  nor (_04308_, _02649_, PC_abstr[3]);
  nor (_04309_, _02390_, _02371_);
  nor (_04310_, _04309_, _02391_);
  and (_04311_, _02649_, _04310_);
  or (_04312_, _04311_, _04308_);
  nand (_04313_, _04312_, _11609_);
  or (_04314_, _11609_, \oc8051_golden_model_1.PC [3]);
  and (_04315_, _04314_, _12493_);
  and (_12623_[3], _04315_, _04313_);
  nor (_04316_, _02367_, \oc8051_golden_model_1.PC [4]);
  nor (_04317_, _04316_, _02677_);
  nor (_04318_, _04317_, _02672_);
  nor (_04319_, _02649_, PC_abstr[4]);
  nor (_04320_, _04319_, _04318_);
  or (_04321_, _04320_, _11613_);
  or (_04322_, _11609_, \oc8051_golden_model_1.PC [4]);
  and (_04323_, _04322_, _12493_);
  and (_12623_[4], _04323_, _04321_);
  nor (_04324_, _02677_, \oc8051_golden_model_1.PC [5]);
  nor (_04325_, _04324_, _02678_);
  nor (_04326_, _04325_, _02672_);
  nor (_04327_, _02649_, PC_abstr[5]);
  nor (_04328_, _04327_, _04326_);
  or (_04329_, _04328_, _11613_);
  or (_04330_, _11609_, \oc8051_golden_model_1.PC [5]);
  and (_04331_, _04330_, _12493_);
  and (_12623_[5], _04331_, _04329_);
  nor (_04332_, _02678_, \oc8051_golden_model_1.PC [6]);
  nor (_04333_, _04332_, _02679_);
  nor (_04334_, _04333_, _02672_);
  nor (_04335_, _02649_, PC_abstr[6]);
  nor (_04336_, _04335_, _04334_);
  or (_04337_, _04336_, _11613_);
  or (_04338_, _11609_, \oc8051_golden_model_1.PC [6]);
  and (_04339_, _04338_, _12493_);
  and (_12623_[6], _04339_, _04337_);
  nor (_04340_, _02679_, \oc8051_golden_model_1.PC [7]);
  nor (_04341_, _04340_, _02680_);
  nor (_04342_, _04341_, _02672_);
  nor (_04343_, _02649_, PC_abstr[7]);
  nor (_04344_, _04343_, _04342_);
  or (_04345_, _04344_, _11613_);
  or (_04346_, _11609_, \oc8051_golden_model_1.PC [7]);
  and (_04347_, _04346_, _12493_);
  and (_12623_[7], _04347_, _04345_);
  nor (_04348_, _02680_, \oc8051_golden_model_1.PC [8]);
  nor (_04349_, _04348_, _02681_);
  nor (_04350_, _04349_, _02672_);
  nor (_04351_, _02649_, PC_abstr[8]);
  nor (_04352_, _04351_, _04350_);
  or (_04353_, _04352_, _11613_);
  or (_04354_, _11609_, \oc8051_golden_model_1.PC [8]);
  and (_04355_, _04354_, _12493_);
  and (_12623_[8], _04355_, _04353_);
  nor (_04357_, _02681_, \oc8051_golden_model_1.PC [9]);
  nor (_04358_, _04357_, _02682_);
  nor (_04359_, _04358_, _02672_);
  nor (_04360_, _02649_, PC_abstr[9]);
  nor (_04361_, _04360_, _04359_);
  or (_04362_, _04361_, _11613_);
  or (_04363_, _11609_, \oc8051_golden_model_1.PC [9]);
  and (_04364_, _04363_, _12493_);
  and (_12623_[9], _04364_, _04362_);
  nor (_04365_, _02682_, \oc8051_golden_model_1.PC [10]);
  nor (_04366_, _04365_, _02683_);
  nor (_04367_, _04366_, _02672_);
  nor (_04368_, _02649_, PC_abstr[10]);
  nor (_04369_, _04368_, _04367_);
  or (_04370_, _04369_, _11613_);
  or (_04371_, _11609_, \oc8051_golden_model_1.PC [10]);
  and (_04372_, _04371_, _12493_);
  and (_12623_[10], _04372_, _04370_);
  nor (_04373_, _02683_, \oc8051_golden_model_1.PC [11]);
  nor (_04374_, _04373_, _02684_);
  nor (_04375_, _04374_, _02672_);
  nor (_04376_, _02649_, PC_abstr[11]);
  nor (_04377_, _04376_, _04375_);
  or (_04378_, _04377_, _11613_);
  or (_04379_, _11609_, \oc8051_golden_model_1.PC [11]);
  and (_04380_, _04379_, _12493_);
  and (_12623_[11], _04380_, _04378_);
  nor (_04381_, _02684_, \oc8051_golden_model_1.PC [12]);
  nor (_04382_, _04381_, _02685_);
  nor (_04383_, _04382_, _02672_);
  nor (_04384_, _02649_, PC_abstr[12]);
  nor (_04385_, _04384_, _04383_);
  or (_04386_, _04385_, _11613_);
  or (_04387_, _11609_, \oc8051_golden_model_1.PC [12]);
  and (_04388_, _04387_, _12493_);
  and (_12623_[12], _04388_, _04386_);
  nor (_04389_, _02685_, \oc8051_golden_model_1.PC [13]);
  nor (_04390_, _04389_, _02686_);
  nor (_04391_, _04390_, _02672_);
  nor (_04392_, _02649_, PC_abstr[13]);
  nor (_04393_, _04392_, _04391_);
  or (_04394_, _04393_, _11613_);
  or (_04395_, _11609_, \oc8051_golden_model_1.PC [13]);
  and (_04396_, _04395_, _12493_);
  and (_12623_[13], _04396_, _04394_);
  nor (_04397_, _02686_, \oc8051_golden_model_1.PC [14]);
  nor (_04398_, _04397_, _02687_);
  nor (_04399_, _04398_, _02672_);
  nor (_04400_, _02649_, PC_abstr[14]);
  nor (_04401_, _04400_, _04399_);
  or (_04402_, _04401_, _11613_);
  or (_04403_, _11609_, \oc8051_golden_model_1.PC [14]);
  and (_04404_, _04403_, _12493_);
  and (_12623_[14], _04404_, _04402_);
  and (_04405_, _02672_, XRAM_DATA_OUT_abstr[0]);
  or (_04406_, _04405_, _11613_);
  or (_04407_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  and (_04408_, _04407_, _12493_);
  and (_12635_[0], _04408_, _04406_);
  and (_04409_, _02672_, XRAM_DATA_OUT_abstr[1]);
  or (_04410_, _04409_, _11613_);
  or (_04411_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  and (_04412_, _04411_, _12493_);
  and (_12635_[1], _04412_, _04410_);
  and (_04413_, _02672_, XRAM_DATA_OUT_abstr[2]);
  or (_04414_, _04413_, _11613_);
  or (_04415_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  and (_04416_, _04415_, _12493_);
  and (_12635_[2], _04416_, _04414_);
  and (_04417_, _02672_, XRAM_DATA_OUT_abstr[3]);
  or (_04418_, _04417_, _11613_);
  or (_04419_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  and (_04420_, _04419_, _12493_);
  and (_12635_[3], _04420_, _04418_);
  and (_04421_, _02672_, XRAM_DATA_OUT_abstr[4]);
  or (_04422_, _04421_, _11613_);
  or (_04423_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  and (_04424_, _04423_, _12493_);
  and (_12635_[4], _04424_, _04422_);
  and (_04425_, _02672_, XRAM_DATA_OUT_abstr[5]);
  or (_04426_, _04425_, _11613_);
  or (_04427_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  and (_04428_, _04427_, _12493_);
  and (_12635_[5], _04428_, _04426_);
  and (_04429_, _02672_, XRAM_DATA_OUT_abstr[6]);
  or (_04430_, _04429_, _11613_);
  or (_04431_, _11609_, \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  and (_04432_, _04431_, _12493_);
  and (_12635_[6], _04432_, _04430_);
  and (_00007_[6], _00903_, _12493_);
  and (_00007_[5], _00943_, _12493_);
  and (_00007_[4], _00927_, _12493_);
  and (_00007_[3], _00919_, _12493_);
  and (_00007_[2], _00910_, _12493_);
  and (_00007_[1], _00950_, _12493_);
  and (_00007_[0], _00934_, _12493_);
  and (_00006_[6], _00737_, _12493_);
  and (_00006_[5], _00769_, _12493_);
  and (_00006_[4], _00785_, _12493_);
  and (_00006_[3], _00754_, _12493_);
  and (_00006_[2], _00745_, _12493_);
  and (_00006_[1], _00776_, _12493_);
  and (_00006_[0], _00792_, _12493_);
  and (_00005_[6], _00865_, _12493_);
  and (_00005_[5], _00832_, _12493_);
  and (_00005_[4], _00848_, _12493_);
  and (_00005_[3], _00888_, _12493_);
  and (_00005_[2], _00872_, _12493_);
  and (_00005_[1], _00839_, _12493_);
  and (_00005_[0], _00855_, _12493_);
  and (_00004_[6], _01015_, _12493_);
  and (_00004_[5], _01032_, _12493_);
  and (_00004_[4], _00991_, _12493_);
  and (_00004_[3], _01007_, _12493_);
  and (_00004_[2], _01023_, _12493_);
  and (_00004_[1], _01039_, _12493_);
  and (_00004_[0], _00998_, _12493_);
  and (_04434_, _11613_, xram_data_in_reg[6]);
  and (_04435_, _11609_, xram_data_in[6]);
  or (_04436_, _04435_, _04434_);
  and (_00010_[6], _04436_, _12493_);
  and (_04437_, _11613_, xram_data_in_reg[5]);
  and (_04438_, _11609_, xram_data_in[5]);
  or (_04439_, _04438_, _04437_);
  and (_00010_[5], _04439_, _12493_);
  and (_04440_, _11613_, xram_data_in_reg[4]);
  and (_04441_, _11609_, xram_data_in[4]);
  or (_04442_, _04441_, _04440_);
  and (_00010_[4], _04442_, _12493_);
  and (_04443_, _11613_, xram_data_in_reg[3]);
  and (_04444_, _11609_, xram_data_in[3]);
  or (_04445_, _04444_, _04443_);
  and (_00010_[3], _04445_, _12493_);
  and (_04446_, _11613_, xram_data_in_reg[2]);
  and (_04447_, _11609_, xram_data_in[2]);
  or (_04448_, _04447_, _04446_);
  and (_00010_[2], _04448_, _12493_);
  and (_04449_, _11613_, xram_data_in_reg[1]);
  and (_04450_, _11609_, xram_data_in[1]);
  or (_04451_, _04450_, _04449_);
  and (_00010_[1], _04451_, _12493_);
  and (_04452_, _11613_, xram_data_in_reg[0]);
  and (_04453_, _11609_, xram_data_in[0]);
  or (_04454_, _04453_, _04452_);
  and (_00010_[0], _04454_, _12493_);
  nor (_04455_, _04177_, _00691_);
  and (_04456_, _04177_, _00691_);
  or (_04457_, _04456_, _04455_);
  nand (_04458_, _07820_, _02703_);
  or (_04459_, _07820_, _02703_);
  and (_04460_, _04459_, _04458_);
  or (_04461_, _07864_, \oc8051_golden_model_1.SP [6]);
  nand (_04462_, _07864_, \oc8051_golden_model_1.SP [6]);
  and (_04463_, _04462_, _04461_);
  or (_04464_, _07858_, \oc8051_golden_model_1.SP [5]);
  nand (_04465_, _07858_, \oc8051_golden_model_1.SP [5]);
  and (_04466_, _04465_, _04464_);
  or (_04467_, _07852_, \oc8051_golden_model_1.SP [4]);
  nand (_04468_, _07852_, \oc8051_golden_model_1.SP [4]);
  and (_04469_, _04468_, _04467_);
  or (_04470_, _07846_, \oc8051_golden_model_1.SP [3]);
  nand (_04471_, _07846_, \oc8051_golden_model_1.SP [3]);
  and (_04472_, _04471_, _04470_);
  nor (_04473_, _07828_, _04204_);
  and (_04474_, _07828_, _04204_);
  or (_04475_, _04474_, _04473_);
  nor (_04476_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_04477_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_04478_, _04477_, _04476_);
  nor (_04479_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_04480_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_04481_, _04480_, _04479_);
  nor (_04482_, _04481_, _04478_);
  and (_04483_, \oc8051_golden_model_1.IRAM[5] [4], _09567_);
  and (_04484_, _03128_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_04485_, _04484_, _04483_);
  and (_04486_, _03923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_04487_, \oc8051_golden_model_1.IRAM[5] [5], _09570_);
  nor (_04488_, _04487_, _04486_);
  and (_04489_, _04488_, _04485_);
  and (_04490_, _04489_, _04482_);
  nor (_04491_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_04492_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_04493_, _04492_, _04491_);
  nand (_04494_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_04495_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_04496_, _04495_, _04494_);
  nor (_04497_, _04496_, _04493_);
  nor (_04498_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_04499_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_04500_, _04499_, _04498_);
  nand (_04501_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_04502_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_04503_, _04502_, _04501_);
  nor (_04504_, _04503_, _04500_);
  and (_04505_, _04504_, _04497_);
  and (_04506_, _04505_, _04490_);
  and (_04507_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_04508_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_04510_, _04508_, _04507_);
  and (_04511_, _03763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_04512_, \oc8051_golden_model_1.IRAM[7] [2], _09607_);
  nor (_04513_, _04512_, _04511_);
  and (_04514_, _04513_, _04510_);
  and (_04515_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_04516_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_04517_, _04516_, _04515_);
  and (_04518_, \oc8051_golden_model_1.IRAM[7] [7], _09387_);
  nor (_04519_, \oc8051_golden_model_1.IRAM[7] [7], _09387_);
  nor (_04520_, _04519_, _04518_);
  and (_04521_, _04520_, _04517_);
  and (_04522_, _04521_, _04514_);
  nor (_04523_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_04524_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_04525_, _04524_, _04523_);
  nor (_04526_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_04527_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_04528_, _04527_, _04526_);
  nor (_04529_, _04528_, _04525_);
  and (_04530_, \oc8051_golden_model_1.IRAM[6] [4], _09588_);
  nor (_04531_, \oc8051_golden_model_1.IRAM[6] [4], _09588_);
  nor (_04532_, _04531_, _04530_);
  and (_04533_, \oc8051_golden_model_1.IRAM[6] [5], _09591_);
  and (_04534_, _03179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_04535_, _04534_, _04533_);
  and (_04536_, _04535_, _04532_);
  and (_04537_, _04536_, _04529_);
  and (_04538_, _04537_, _04522_);
  and (_04539_, _04538_, _04506_);
  nor (_04540_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_04541_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_04542_, _04541_, _04540_);
  not (_04543_, _04542_);
  and (_04544_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_04545_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_04546_, _04545_, _04544_);
  and (_04547_, _04546_, _04543_);
  nor (_04548_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_04549_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_04550_, _04549_, _04548_);
  not (_04551_, _04550_);
  and (_04552_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_04553_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_04554_, _04553_, _04552_);
  and (_04555_, _04554_, _04551_);
  and (_04556_, _04555_, _04547_);
  and (_04557_, _02810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_04558_, \oc8051_golden_model_1.IRAM[0] [0], _09442_);
  nor (_04559_, _04558_, _04557_);
  and (_04560_, \oc8051_golden_model_1.IRAM[0] [1], _09446_);
  and (_04561_, _02822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_04562_, _04561_, _04560_);
  and (_04563_, _04562_, _04559_);
  nor (_04564_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_04565_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_04566_, _04565_, _04564_);
  nor (_04567_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_04568_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_04569_, _04568_, _04567_);
  nor (_04570_, _04569_, _04566_);
  and (_04571_, _04570_, _04563_);
  and (_04572_, _04571_, _04556_);
  and (_04573_, _02991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_04574_, \oc8051_golden_model_1.IRAM[3] [0], _09512_);
  nor (_04575_, _04574_, _04573_);
  and (_04576_, \oc8051_golden_model_1.IRAM[3] [1], _09515_);
  nor (_04577_, \oc8051_golden_model_1.IRAM[3] [1], _09515_);
  nor (_04578_, _04577_, _04576_);
  and (_04579_, _04578_, _04575_);
  nor (_04580_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_04581_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_04582_, _04581_, _04580_);
  nor (_04583_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_04584_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_04585_, _04584_, _04583_);
  nor (_04586_, _04585_, _04582_);
  and (_04587_, _04586_, _04579_);
  and (_04588_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_04589_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_04590_, _04589_, _04588_);
  nor (_04591_, \oc8051_golden_model_1.IRAM[2] [2], _09495_);
  and (_04592_, \oc8051_golden_model_1.IRAM[2] [2], _09495_);
  nor (_04593_, _04592_, _04591_);
  and (_04594_, _04593_, _04590_);
  and (_04595_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_04596_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_04597_, _04596_, _04595_);
  nor (_04598_, \oc8051_golden_model_1.IRAM[2] [7], _09508_);
  and (_04599_, \oc8051_golden_model_1.IRAM[2] [7], _09508_);
  nor (_04600_, _04599_, _04598_);
  and (_04601_, _04600_, _04597_);
  and (_04602_, _04601_, _04594_);
  and (_04603_, _04602_, _04587_);
  and (_04604_, _04603_, _04572_);
  and (_04605_, _04604_, _04539_);
  nor (_04606_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_04607_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_04608_, _04607_, _04606_);
  nand (_04609_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_04611_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_04612_, _04611_, _04609_);
  nor (_04613_, _04612_, _04608_);
  nor (_04614_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_04615_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_04616_, _04615_, _04614_);
  nand (_04617_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_04618_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_04619_, _04618_, _04617_);
  nor (_04620_, _04619_, _04616_);
  and (_04621_, _04620_, _04613_);
  and (_04622_, _03433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_04623_, \oc8051_golden_model_1.IRAM[12] [0], _09708_);
  nor (_04624_, _04623_, _04622_);
  and (_04625_, _03726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_04626_, \oc8051_golden_model_1.IRAM[12] [1], _09711_);
  nor (_04627_, _04626_, _04625_);
  and (_04628_, _04627_, _04624_);
  nor (_04629_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_04630_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_04631_, _04630_, _04629_);
  nor (_04632_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_04633_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_04634_, _04633_, _04632_);
  nor (_04635_, _04634_, _04631_);
  and (_04636_, _04635_, _04628_);
  and (_04637_, _04636_, _04621_);
  and (_04638_, _03675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_04639_, \oc8051_golden_model_1.IRAM[15] [0], _09774_);
  nor (_04640_, _04639_, _04638_);
  and (_04641_, _03732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_04642_, \oc8051_golden_model_1.IRAM[15] [1], _09777_);
  nor (_04643_, _04642_, _04641_);
  and (_04644_, _04643_, _04640_);
  nor (_04645_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_04646_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_04647_, _04646_, _04645_);
  nor (_04648_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_04649_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_04650_, _04649_, _04648_);
  nor (_04651_, _04650_, _04647_);
  and (_04652_, _04651_, _04644_);
  and (_04653_, \oc8051_golden_model_1.IRAM[14] [2], _09757_);
  nor (_04654_, \oc8051_golden_model_1.IRAM[14] [2], _09757_);
  nor (_04655_, _04654_, _04653_);
  nand (_04656_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_04657_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_04658_, _04657_, _04656_);
  not (_04659_, _04658_);
  and (_04660_, _04659_, _04655_);
  and (_04661_, _03566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_04662_, \oc8051_golden_model_1.IRAM[14] [7], _09412_);
  nor (_04663_, _04662_, _04661_);
  nand (_04664_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_04665_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_04666_, _04665_, _04664_);
  not (_04667_, _04666_);
  and (_04668_, _04667_, _04663_);
  and (_04669_, _04668_, _04660_);
  and (_04670_, _04669_, _04652_);
  and (_04671_, _04670_, _04637_);
  and (_04672_, _03324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_04673_, \oc8051_golden_model_1.IRAM[9] [5], _09655_);
  nor (_04674_, _04673_, _04672_);
  and (_04675_, _03318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_04676_, \oc8051_golden_model_1.IRAM[9] [4], _09652_);
  nor (_04677_, _04676_, _04675_);
  and (_04678_, _04677_, _04674_);
  nor (_04679_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_04680_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_04681_, _04680_, _04679_);
  nor (_04682_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_04683_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_04684_, _04683_, _04682_);
  nor (_04685_, _04684_, _04681_);
  and (_04686_, _04685_, _04678_);
  nor (_04687_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_04688_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_04689_, _04688_, _04687_);
  nor (_04690_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_04691_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_04692_, _04691_, _04690_);
  nor (_04693_, _04692_, _04689_);
  nor (_04694_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_04695_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_04696_, _04695_, _04694_);
  nor (_04697_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_04698_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_04699_, _04698_, _04697_);
  nor (_04700_, _04699_, _04696_);
  and (_04701_, _04700_, _04693_);
  and (_04702_, _04701_, _04686_);
  and (_04703_, \oc8051_golden_model_1.IRAM[11] [2], _09691_);
  and (_04704_, _03401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_04705_, _04704_, _04703_);
  nand (_04706_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_04707_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_04708_, _04707_, _04706_);
  not (_04709_, _04708_);
  and (_04710_, _04709_, _04705_);
  nor (_04712_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_04713_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_04714_, _04713_, _04712_);
  not (_04715_, _04714_);
  and (_04716_, _02774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_04717_, \oc8051_golden_model_1.IRAM[11] [7], _09704_);
  nor (_04718_, _04717_, _04716_);
  and (_04719_, _04718_, _04715_);
  and (_04720_, _04719_, _04710_);
  nor (_04721_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_04722_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_04723_, _04722_, _04721_);
  nor (_04724_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_04725_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_04726_, _04725_, _04724_);
  nor (_04727_, _04726_, _04723_);
  nor (_04728_, \oc8051_golden_model_1.IRAM[10] [5], _09677_);
  and (_04729_, \oc8051_golden_model_1.IRAM[10] [5], _09677_);
  nor (_04730_, _04729_, _04728_);
  nor (_04731_, \oc8051_golden_model_1.IRAM[10] [4], _09674_);
  and (_04732_, \oc8051_golden_model_1.IRAM[10] [4], _09674_);
  nor (_04733_, _04732_, _04731_);
  and (_04734_, _04733_, _04730_);
  and (_04735_, _04734_, _04727_);
  and (_04736_, _04735_, _04720_);
  and (_04737_, _04736_, _04702_);
  and (_04738_, _04737_, _04671_);
  and (_04739_, _04738_, _04605_);
  nor (_04740_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_04741_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_04742_, _04741_, _04740_);
  nand (_04743_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_04744_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_04745_, _04744_, _04743_);
  nor (_04746_, _04745_, _04742_);
  nor (_04747_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_04748_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_04749_, _04748_, _04747_);
  not (_04750_, _04749_);
  and (_04751_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_04752_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_04753_, _04752_, _04751_);
  and (_04754_, _04753_, _04750_);
  and (_04755_, _04754_, _04746_);
  and (_04756_, _03042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_04757_, \oc8051_golden_model_1.IRAM[4] [0], _09535_);
  nor (_04758_, _04757_, _04756_);
  and (_04759_, _03702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_04760_, \oc8051_golden_model_1.IRAM[4] [1], _09538_);
  nor (_04761_, _04760_, _04759_);
  and (_04762_, _04761_, _04758_);
  nor (_04763_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_04764_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_04765_, _04764_, _04763_);
  nor (_04766_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_04767_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_04768_, _04767_, _04766_);
  nor (_04769_, _04768_, _04765_);
  and (_04770_, _04769_, _04762_);
  and (_04771_, _04770_, _04755_);
  and (_04772_, _03708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_04773_, \oc8051_golden_model_1.IRAM[7] [1], _09604_);
  nor (_04774_, _04773_, _04772_);
  and (_04775_, _03195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_04776_, \oc8051_golden_model_1.IRAM[7] [0], _09601_);
  nor (_04777_, _04776_, _04775_);
  and (_04778_, _04777_, _04774_);
  nor (_04779_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_04780_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_04781_, _04780_, _04779_);
  nor (_04782_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_04783_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_04784_, _04783_, _04782_);
  nor (_04785_, _04784_, _04781_);
  and (_04786_, _04785_, _04778_);
  and (_04787_, \oc8051_golden_model_1.IRAM[6] [2], _09583_);
  nor (_04788_, \oc8051_golden_model_1.IRAM[6] [2], _09583_);
  nor (_04789_, _04788_, _04787_);
  and (_04790_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_04791_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_04792_, _04791_, _04790_);
  and (_04793_, _04792_, _04789_);
  nor (_04794_, \oc8051_golden_model_1.IRAM[6] [7], _09597_);
  and (_04795_, \oc8051_golden_model_1.IRAM[6] [7], _09597_);
  nor (_04796_, _04795_, _04794_);
  nand (_04797_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_04798_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_04799_, _04798_, _04797_);
  not (_04800_, _04799_);
  and (_04801_, _04800_, _04796_);
  and (_04802_, _04801_, _04793_);
  and (_04803_, _04802_, _04786_);
  and (_04804_, _04803_, _04771_);
  nor (_04805_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_04806_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_04807_, _04806_, _04805_);
  nor (_04808_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_04809_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_04810_, _04809_, _04808_);
  nor (_04811_, _04810_, _04807_);
  and (_04812_, _03858_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_04813_, \oc8051_golden_model_1.IRAM[1] [4], _09478_);
  nor (_04814_, _04813_, _04812_);
  and (_04815_, _03912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_04816_, \oc8051_golden_model_1.IRAM[1] [5], _09481_);
  nor (_04817_, _04816_, _04815_);
  and (_04818_, _04817_, _04814_);
  and (_04819_, _04818_, _04811_);
  nor (_04820_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_04821_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_04822_, _04821_, _04820_);
  not (_04823_, _04822_);
  and (_04824_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_04825_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_04826_, _04825_, _04824_);
  and (_04827_, _04826_, _04823_);
  nor (_04828_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_04829_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_04830_, _04829_, _04828_);
  not (_04831_, _04830_);
  and (_04832_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_04833_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_04834_, _04833_, _04832_);
  and (_04835_, _04834_, _04831_);
  and (_04836_, _04835_, _04827_);
  and (_04837_, _04836_, _04819_);
  and (_04838_, \oc8051_golden_model_1.IRAM[3] [2], _09518_);
  nor (_04839_, \oc8051_golden_model_1.IRAM[3] [2], _09518_);
  nor (_04840_, _04839_, _04838_);
  nand (_04841_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_04842_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_04843_, _04842_, _04841_);
  not (_04844_, _04843_);
  and (_04845_, _04844_, _04840_);
  and (_04846_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_04847_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_04848_, _04847_, _04846_);
  and (_04849_, _02760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_04850_, \oc8051_golden_model_1.IRAM[3] [7], _09375_);
  nor (_04851_, _04850_, _04849_);
  and (_04852_, _04851_, _04848_);
  and (_04853_, _04852_, _04845_);
  nor (_04854_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_04855_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_04856_, _04855_, _04854_);
  nor (_04857_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_04858_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_04859_, _04858_, _04857_);
  nor (_04860_, _04859_, _04856_);
  nor (_04861_, \oc8051_golden_model_1.IRAM[2] [5], _09503_);
  and (_04862_, \oc8051_golden_model_1.IRAM[2] [5], _09503_);
  nor (_04863_, _04862_, _04861_);
  nor (_04864_, \oc8051_golden_model_1.IRAM[2] [4], _09500_);
  and (_04865_, \oc8051_golden_model_1.IRAM[2] [4], _09500_);
  nor (_04866_, _04865_, _04864_);
  and (_04867_, _04866_, _04863_);
  and (_04868_, _04867_, _04860_);
  and (_04869_, _04868_, _04853_);
  and (_04870_, _04869_, _04837_);
  and (_04871_, _04870_, _04804_);
  nor (_04872_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_04873_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_04874_, _04873_, _04872_);
  nor (_04875_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_04876_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_04877_, _04876_, _04875_);
  nor (_04878_, _04877_, _04874_);
  and (_04879_, _03891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_04880_, \oc8051_golden_model_1.IRAM[13] [4], _09740_);
  nor (_04881_, _04880_, _04879_);
  and (_04882_, \oc8051_golden_model_1.IRAM[13] [5], _09743_);
  and (_04883_, _03509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_04884_, _04883_, _04882_);
  and (_04885_, _04884_, _04881_);
  and (_04886_, _04885_, _04878_);
  nor (_04887_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_04888_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_04889_, _04888_, _04887_);
  nand (_04890_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_04891_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_04892_, _04891_, _04890_);
  nor (_04893_, _04892_, _04889_);
  nor (_04894_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_04895_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_04896_, _04895_, _04894_);
  nand (_04897_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_04898_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_04899_, _04898_, _04897_);
  nor (_04900_, _04899_, _04896_);
  and (_04901_, _04900_, _04893_);
  and (_04902_, _04901_, _04886_);
  and (_04903_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_04904_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_04905_, _04904_, _04903_);
  and (_04906_, _03586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_04907_, \oc8051_golden_model_1.IRAM[15] [2], _09780_);
  nor (_04908_, _04907_, _04906_);
  and (_04909_, _04908_, _04905_);
  and (_04910_, \oc8051_golden_model_1.IRAM[15] [7], _09434_);
  and (_04911_, _02364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_04912_, _04911_, _04910_);
  nand (_04913_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_04914_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_04915_, _04914_, _04913_);
  not (_04916_, _04915_);
  and (_04917_, _04916_, _04912_);
  and (_04918_, _04917_, _04909_);
  nor (_04919_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_04920_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_04921_, _04920_, _04919_);
  nor (_04922_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_04923_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_04924_, _04923_, _04922_);
  nor (_04925_, _04924_, _04921_);
  nor (_04926_, \oc8051_golden_model_1.IRAM[14] [4], _09763_);
  and (_04927_, \oc8051_golden_model_1.IRAM[14] [4], _09763_);
  nor (_04928_, _04927_, _04926_);
  and (_04929_, \oc8051_golden_model_1.IRAM[14] [5], _09766_);
  nor (_04930_, \oc8051_golden_model_1.IRAM[14] [5], _09766_);
  nor (_04931_, _04930_, _04929_);
  and (_04932_, _04931_, _04928_);
  and (_04933_, _04932_, _04925_);
  and (_04934_, _04933_, _04918_);
  and (_04935_, _04934_, _04902_);
  nor (_04936_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_04937_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_04938_, _04937_, _04936_);
  nor (_04939_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_04940_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_04941_, _04940_, _04939_);
  nor (_04942_, _04941_, _04938_);
  nor (_04943_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_04944_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_04945_, _04944_, _04943_);
  nor (_04946_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_04947_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_04948_, _04947_, _04946_);
  nor (_04949_, _04948_, _04945_);
  and (_04950_, _04949_, _04942_);
  and (_04951_, _03241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_04952_, \oc8051_golden_model_1.IRAM[8] [0], _09623_);
  nor (_04953_, _04952_, _04951_);
  and (_04954_, \oc8051_golden_model_1.IRAM[8] [1], _09626_);
  nor (_04955_, \oc8051_golden_model_1.IRAM[8] [1], _09626_);
  nor (_04956_, _04955_, _04954_);
  and (_04957_, _04956_, _04953_);
  nor (_04958_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_04959_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_04960_, _04959_, _04958_);
  nor (_04961_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_04962_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_04963_, _04962_, _04961_);
  nor (_04964_, _04963_, _04960_);
  and (_04965_, _04964_, _04957_);
  and (_04966_, _04965_, _04950_);
  and (_04967_, _03386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_04968_, \oc8051_golden_model_1.IRAM[11] [0], _09685_);
  nor (_04969_, _04968_, _04967_);
  and (_04970_, \oc8051_golden_model_1.IRAM[11] [1], _09688_);
  nor (_04971_, \oc8051_golden_model_1.IRAM[11] [1], _09688_);
  nor (_04972_, _04971_, _04970_);
  and (_04973_, _04972_, _04969_);
  nor (_04974_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_04975_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_04976_, _04975_, _04974_);
  nor (_04977_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_04978_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_04979_, _04978_, _04977_);
  nor (_04980_, _04979_, _04976_);
  and (_04981_, _04980_, _04973_);
  nor (_04982_, \oc8051_golden_model_1.IRAM[10] [2], _09668_);
  and (_04983_, \oc8051_golden_model_1.IRAM[10] [2], _09668_);
  nor (_04984_, _04983_, _04982_);
  nand (_04985_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_04986_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_04987_, _04986_, _04985_);
  not (_04988_, _04987_);
  and (_04989_, _04988_, _04984_);
  nor (_04990_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_04991_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_04992_, _04991_, _04990_);
  not (_04993_, _04992_);
  nor (_04994_, \oc8051_golden_model_1.IRAM[10] [7], _09401_);
  and (_04995_, \oc8051_golden_model_1.IRAM[10] [7], _09401_);
  nor (_04996_, _04995_, _04994_);
  and (_04997_, _04996_, _04993_);
  and (_04998_, _04997_, _04989_);
  and (_04999_, _04998_, _04981_);
  and (_05000_, _04999_, _04966_);
  and (_05001_, _05000_, _04935_);
  and (_05002_, _05001_, _04871_);
  and (_05003_, _05002_, _04739_);
  nor (_05004_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_05005_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_05006_, _05005_, _05004_);
  nor (_05007_, \oc8051_golden_model_1.DPL [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_05008_, \oc8051_golden_model_1.DPL [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_05009_, _05008_, _05007_);
  nor (_05010_, _05009_, _05006_);
  nor (_05011_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_05012_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_05013_, _05012_, _05011_);
  nor (_05014_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_05015_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_05016_, _05015_, _05014_);
  nor (_05017_, _05016_, _05013_);
  and (_05018_, _05017_, _05010_);
  and (_05019_, _04027_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_05020_, \oc8051_golden_model_1.DPL [2], _08190_);
  nor (_05021_, _05020_, _05019_);
  and (_05022_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_05023_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_05024_, _05023_, _05022_);
  and (_05025_, _05024_, _05021_);
  and (_05026_, _02731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_05027_, \oc8051_golden_model_1.DPL [7], _07966_);
  nor (_05028_, _05027_, _05026_);
  and (_05029_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_05030_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_05031_, _05030_, _05029_);
  and (_05032_, _05031_, _05028_);
  and (_05033_, _05032_, _05025_);
  and (_05034_, _05033_, _05018_);
  nor (_05035_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_05036_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_05037_, _05036_, _05035_);
  nor (_05038_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_05039_, \oc8051_golden_model_1.ACC [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_05040_, _05039_, _05038_);
  nor (_05041_, _05040_, _05037_);
  nor (_05042_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_05043_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05044_, _05043_, _05042_);
  nor (_05045_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_05046_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_05047_, _05046_, _05045_);
  nor (_05048_, _05047_, _05044_);
  and (_05049_, _05048_, _05041_);
  and (_05050_, _03797_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_05051_, \oc8051_golden_model_1.ACC [2], _05760_);
  nor (_05052_, _05051_, _05050_);
  and (_05053_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_05054_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_05055_, _05054_, _05053_);
  and (_05056_, _05055_, _05052_);
  and (_05057_, _02735_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_05058_, \oc8051_golden_model_1.ACC [7], _05679_);
  nor (_05059_, _05058_, _05057_);
  and (_05060_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05061_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_05062_, _05061_, _05060_);
  and (_05063_, _05062_, _05059_);
  and (_05064_, _05063_, _05056_);
  and (_05065_, _05064_, _05049_);
  and (_05066_, _05065_, _05034_);
  nor (_05067_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_05068_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_05069_, _05068_, _05067_);
  nor (_05070_, \oc8051_golden_model_1.DPH [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_05071_, \oc8051_golden_model_1.DPH [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor (_05072_, _05071_, _05070_);
  nor (_05073_, _05072_, _05069_);
  nor (_05074_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_05075_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nor (_05076_, _05075_, _05074_);
  nor (_05077_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_05078_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nor (_05079_, _05078_, _05077_);
  nor (_05080_, _05079_, _05076_);
  and (_05081_, _05080_, _05073_);
  and (_05082_, _04049_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_05083_, _04049_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_05084_, _05083_, _05082_);
  and (_05085_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor (_05086_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_05087_, _05086_, _05085_);
  and (_05088_, _05087_, _05084_);
  and (_05089_, _02727_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_05090_, _02727_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_05091_, _05090_, _05089_);
  and (_05092_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nor (_05093_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_05094_, _05093_, _05092_);
  and (_05095_, _05094_, _05091_);
  and (_05096_, _05095_, _05088_);
  and (_05097_, _05096_, _05081_);
  nor (_05098_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_05099_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_05100_, _05099_, _05098_);
  nor (_05101_, \oc8051_golden_model_1.B [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_05102_, \oc8051_golden_model_1.B [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_05103_, _05102_, _05101_);
  nor (_05104_, _05103_, _05100_);
  nor (_05105_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_05106_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_05107_, _05106_, _05105_);
  nor (_05108_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_05109_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_05110_, _05109_, _05108_);
  nor (_05111_, _05110_, _05107_);
  and (_05112_, _05111_, _05104_);
  and (_05113_, _03622_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_05114_, \oc8051_golden_model_1.B [2], _07003_);
  nor (_05115_, _05114_, _05113_);
  and (_05116_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_05117_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_05118_, _05117_, _05116_);
  and (_05119_, _05118_, _05115_);
  and (_05120_, _02800_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_05121_, \oc8051_golden_model_1.B [7], _06778_);
  nor (_05122_, _05121_, _05120_);
  and (_05123_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_05124_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_05125_, _05124_, _05123_);
  and (_05126_, _05125_, _05122_);
  and (_05127_, _05126_, _05119_);
  and (_05128_, _05127_, _05112_);
  and (_05129_, _05128_, _05097_);
  and (_05130_, _05129_, _05066_);
  nor (_05131_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_05132_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_05133_, _05132_, _05131_);
  nor (_05134_, \oc8051_golden_model_1.P2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_05135_, \oc8051_golden_model_1.P2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_05136_, _05135_, _05134_);
  nor (_05137_, _05136_, _05133_);
  nor (_05138_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_05139_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_05140_, _05139_, _05138_);
  nor (_05141_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_05142_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_05143_, _05142_, _05141_);
  nor (_05144_, _05143_, _05140_);
  and (_05145_, _05144_, _05137_);
  and (_05146_, _04115_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_05147_, \oc8051_golden_model_1.P2 [2], _08703_);
  nor (_05148_, _05147_, _05146_);
  and (_05149_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_05150_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_05151_, _05150_, _05149_);
  and (_05152_, _05151_, _05148_);
  and (_05153_, _02715_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_05154_, \oc8051_golden_model_1.P2 [7], _08473_);
  nor (_05155_, _05154_, _05153_);
  and (_05156_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_05157_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_05158_, _05157_, _05156_);
  and (_05159_, _05158_, _05155_);
  and (_05160_, _05159_, _05152_);
  and (_05161_, _05160_, _05145_);
  nor (_05162_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_05163_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_05164_, _05163_, _05162_);
  nor (_05165_, \oc8051_golden_model_1.P0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_05166_, \oc8051_golden_model_1.P0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_05167_, _05166_, _05165_);
  nor (_05168_, _05167_, _05164_);
  nor (_05169_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_05170_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_05171_, _05170_, _05169_);
  nor (_05172_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_05173_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_05174_, _05173_, _05172_);
  nor (_05175_, _05174_, _05171_);
  and (_05176_, _05175_, _05168_);
  and (_05177_, _04071_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_05178_, \oc8051_golden_model_1.P0 [2], _08533_);
  nor (_05179_, _05178_, _05177_);
  and (_05180_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_05181_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_05182_, _05181_, _05180_);
  and (_05183_, _05182_, _05179_);
  and (_05184_, _02723_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_05185_, \oc8051_golden_model_1.P0 [7], _08443_);
  nor (_05186_, _05185_, _05184_);
  and (_05187_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_05188_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_05189_, _05188_, _05187_);
  and (_05190_, _05189_, _05186_);
  and (_05191_, _05190_, _05183_);
  and (_05192_, _05191_, _05176_);
  and (_05193_, _05192_, _05161_);
  nor (_05194_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_05195_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_05196_, _05195_, _05194_);
  nor (_05197_, \oc8051_golden_model_1.P3 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_05198_, \oc8051_golden_model_1.P3 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_05199_, _05198_, _05197_);
  nor (_05200_, _05199_, _05196_);
  nor (_05201_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_05202_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_05203_, _05202_, _05201_);
  nor (_05204_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_05205_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_05206_, _05205_, _05204_);
  nor (_05207_, _05206_, _05203_);
  and (_05208_, _05207_, _05200_);
  and (_05209_, _04137_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_05210_, \oc8051_golden_model_1.P3 [2], _08787_);
  nor (_05211_, _05210_, _05209_);
  and (_05212_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_05213_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_05214_, _05213_, _05212_);
  and (_05215_, _05214_, _05211_);
  and (_05216_, _02711_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_05217_, \oc8051_golden_model_1.P3 [7], _08481_);
  nor (_05218_, _05217_, _05216_);
  and (_05219_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_05220_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_05221_, _05220_, _05219_);
  and (_05222_, _05221_, _05218_);
  and (_05223_, _05222_, _05215_);
  and (_05224_, _05223_, _05208_);
  nor (_05225_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_05226_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_05227_, _05226_, _05225_);
  nor (_05228_, \oc8051_golden_model_1.P1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_05229_, \oc8051_golden_model_1.P1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_05230_, _05229_, _05228_);
  nor (_05231_, _05230_, _05227_);
  nor (_05232_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_05233_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_05234_, _05233_, _05232_);
  nor (_05235_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_05236_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_05237_, _05236_, _05235_);
  nor (_05238_, _05237_, _05234_);
  and (_05239_, _05238_, _05231_);
  and (_05240_, _04093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_05241_, \oc8051_golden_model_1.P1 [2], _08618_);
  nor (_05242_, _05241_, _05240_);
  and (_05243_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_05244_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_05245_, _05244_, _05243_);
  and (_05246_, _05245_, _05242_);
  and (_05247_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_05248_, \oc8051_golden_model_1.P1 [7], _08453_);
  nor (_05249_, _05248_, _05247_);
  and (_05250_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_05251_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_05252_, _05251_, _05250_);
  and (_05253_, _05252_, _05249_);
  and (_05254_, _05253_, _05246_);
  and (_05255_, _05254_, _05239_);
  and (_05256_, _05255_, _05224_);
  and (_05257_, _05256_, _05193_);
  and (_05258_, _05257_, _05130_);
  and (_05259_, _05258_, _05003_);
  and (_05260_, _02672_, PSW_abstr[2]);
  and (_05261_, _02649_, \oc8051_golden_model_1.PSW [2]);
  nor (_05262_, _05261_, _05260_);
  and (_05263_, _05262_, _08262_);
  nor (_05264_, _05262_, _08262_);
  or (_05265_, _05264_, _05263_);
  nor (_05266_, _02649_, PSW_abstr[1]);
  and (_05267_, _02649_, _04181_);
  or (_05268_, _05267_, _05266_);
  and (_05269_, _05268_, _08227_);
  nor (_05270_, _05268_, _08227_);
  or (_05271_, _05270_, _05269_);
  and (_05272_, _02672_, PSW_abstr[6]);
  and (_05273_, _02649_, \oc8051_golden_model_1.PSW [6]);
  nor (_05274_, _05273_, _05272_);
  and (_05275_, _05274_, _07055_);
  nor (_05276_, _05274_, _07055_);
  or (_05277_, _05276_, _05275_);
  and (_05278_, _05277_, _05271_);
  and (_05279_, _05278_, _05265_);
  nor (_05280_, _02649_, PSW_abstr[5]);
  and (_05281_, _02649_, _04196_);
  or (_05282_, _05281_, _05280_);
  or (_05283_, _05282_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_05284_, _05282_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_05285_, _05284_, _05283_);
  nor (_05286_, _02649_, PSW_abstr[4]);
  and (_05287_, _02649_, _04192_);
  or (_05288_, _05287_, _05286_);
  or (_05289_, _05288_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand (_05290_, _05288_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_05291_, _05290_, _05289_);
  and (_05292_, _05291_, _05285_);
  and (_05293_, _02672_, PSW_abstr[3]);
  nor (_05294_, _05293_, _02752_);
  nand (_05295_, _05294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_05296_, _05294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_05297_, _05296_, _05295_);
  nor (_05298_, _02649_, PSW_abstr[7]);
  and (_05299_, _02649_, _02706_);
  or (_05300_, _05299_, _05298_);
  and (_05301_, _05300_, _08218_);
  nor (_05302_, _05300_, _08218_);
  or (_05303_, _05302_, _05301_);
  and (_05304_, _05303_, _05297_);
  and (_05305_, _05304_, _05292_);
  and (_05306_, _05305_, _05279_);
  and (_05307_, _05306_, _05259_);
  and (_05308_, _05307_, _04475_);
  or (_05309_, _07834_, \oc8051_golden_model_1.SP [1]);
  nand (_05310_, _07834_, \oc8051_golden_model_1.SP [1]);
  and (_05311_, _05310_, _05309_);
  and (_05312_, _05311_, _05308_);
  nand (_05313_, _07840_, \oc8051_golden_model_1.SP [2]);
  or (_05314_, _07840_, \oc8051_golden_model_1.SP [2]);
  and (_05315_, _05314_, _05313_);
  and (_05316_, _05315_, _05312_);
  and (_05317_, _05316_, _04472_);
  and (_05318_, _05317_, _04469_);
  and (_05319_, _05318_, _04466_);
  and (_05320_, _05319_, _04463_);
  and (_05321_, _05320_, _04460_);
  nand (_05322_, _05321_, _04457_);
  nand (_05323_, _05322_, inst_finished_r);
  and (_05324_, _05323_, eq_state_2);
  or (_00001_, _05324_, rst);
  and (_05325_, _02693_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_05326_, _02693_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_05327_, _05326_, _05325_);
  nor (_05328_, _04401_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_05329_, _04401_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_05330_, _05329_, _05328_);
  nor (_05331_, _04385_, _07936_);
  and (_05332_, _04385_, _07936_);
  or (_05333_, _05332_, _05331_);
  nor (_05334_, _04320_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_05335_, _04320_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_05336_, _05335_, _05334_);
  nor (_05337_, _04296_, _05879_);
  and (_05338_, _04296_, _05879_);
  nor (_05339_, _05338_, _05337_);
  nor (_05340_, _04312_, _05782_);
  and (_05341_, _04312_, _05782_);
  nor (_05342_, _05341_, _05340_);
  or (_05343_, _05342_, _05339_);
  or (_05344_, _05343_, _05336_);
  and (_05345_, _04289_, _05929_);
  nor (_05346_, _04361_, _07925_);
  or (_05347_, _05346_, _05345_);
  nor (_05348_, _04344_, _05852_);
  and (_05349_, _04361_, _07925_);
  or (_05350_, _05349_, _05348_);
  or (_05351_, _05350_, _05347_);
  nor (_05352_, _04352_, _07919_);
  and (_05353_, _04352_, _07919_);
  nor (_05354_, _05353_, _05352_);
  nor (_05355_, _04289_, _05929_);
  and (_05356_, _04344_, _05852_);
  nor (_05357_, _05356_, _05355_);
  nand (_05358_, _05357_, _05354_);
  or (_05359_, _05358_, _05351_);
  or (_05360_, _05359_, _05344_);
  or (_05361_, _05360_, _05333_);
  nor (_05362_, _04393_, _07911_);
  and (_05363_, _04393_, _07911_);
  or (_05364_, _05363_, _05362_);
  nor (_05365_, _04377_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_05366_, _04377_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_05367_, _05366_, _05365_);
  nor (_05368_, _04304_, _05897_);
  and (_05369_, _04304_, _05897_);
  nor (_05370_, _05369_, _05368_);
  nor (_05371_, _04336_, _05821_);
  and (_05372_, _04336_, _05821_);
  nor (_05373_, _05372_, _05371_);
  nand (_05374_, _05373_, _05370_);
  nor (_05375_, _04328_, _05800_);
  and (_05376_, _04328_, _05800_);
  nor (_05377_, _05376_, _05375_);
  nor (_05378_, _04369_, _07930_);
  and (_05379_, _04369_, _07930_);
  nor (_05380_, _05379_, _05378_);
  nand (_05381_, _05380_, _05377_);
  or (_05382_, _05381_, _05374_);
  or (_05383_, _05382_, _05367_);
  or (_05384_, _05383_, _05364_);
  or (_05385_, _05384_, _05361_);
  or (_05386_, _05385_, _05330_);
  nor (_05387_, _05386_, _05327_);
  nor (_05388_, _05387_, _11613_);
  nor (_05389_, _04409_, _00487_);
  and (_05390_, _04409_, _00487_);
  nor (_05391_, _05390_, _05389_);
  nor (_05392_, _04429_, _00517_);
  and (_05393_, _04429_, _00517_);
  nor (_05394_, _05393_, _05392_);
  and (_05395_, _05394_, _05391_);
  nor (_05396_, _04405_, _00481_);
  and (_05397_, _04405_, _00481_);
  nor (_05398_, _05397_, _05396_);
  nor (_05399_, _02673_, _12174_);
  and (_05400_, _02673_, _12174_);
  nor (_05401_, _05400_, _05399_);
  and (_05402_, _05401_, _05398_);
  and (_05403_, _05402_, _05395_);
  nor (_05404_, _04413_, _00492_);
  and (_05405_, _04413_, _00492_);
  nor (_05406_, _05405_, _05404_);
  nor (_05407_, _04421_, _00503_);
  and (_05408_, _04421_, _00503_);
  nor (_05409_, _05408_, _05407_);
  and (_05410_, _05409_, _05406_);
  nor (_05411_, _04417_, _00497_);
  and (_05412_, _04417_, _00497_);
  nor (_05413_, _05412_, _05411_);
  nor (_05414_, _04425_, _00510_);
  and (_05415_, _04425_, _00510_);
  nor (_05416_, _05415_, _05414_);
  and (_05417_, _05416_, _05413_);
  and (_05418_, _05417_, _05410_);
  and (_05419_, _05418_, _05403_);
  nor (_05420_, _04262_, _00588_);
  and (_05421_, _04262_, _00588_);
  nor (_05422_, _05421_, _05420_);
  nor (_05423_, _04271_, _00598_);
  and (_05424_, _04271_, _00598_);
  or (_05425_, _05424_, _05423_);
  not (_05426_, _05425_);
  and (_05427_, _05426_, _05422_);
  nor (_05428_, _02697_, _12184_);
  and (_05429_, _02697_, _12184_);
  nor (_05430_, _05429_, _05428_);
  nor (_05431_, _04275_, _00603_);
  and (_05432_, _04275_, _00603_);
  nor (_05433_, _05432_, _05431_);
  and (_05434_, _05433_, _05430_);
  and (_05435_, _05434_, _05427_);
  nor (_05436_, _04226_, _00524_);
  and (_05437_, _04226_, _00524_);
  nor (_05438_, _05437_, _05436_);
  nor (_05439_, _04234_, _00540_);
  and (_05440_, _04234_, _00540_);
  nor (_05441_, _05440_, _05439_);
  and (_05442_, _05441_, _05438_);
  nor (_05443_, _04246_, _00562_);
  and (_05444_, _04246_, _00562_);
  nor (_05445_, _05444_, _05443_);
  nor (_05446_, _04254_, _00576_);
  and (_05447_, _04254_, _00576_);
  nor (_05448_, _05447_, _05446_);
  and (_05449_, _05448_, _05445_);
  and (_05450_, _05449_, _05442_);
  and (_05451_, _05450_, _05435_);
  nor (_05452_, _04258_, _00583_);
  and (_05453_, _04258_, _00583_);
  nor (_05454_, _05453_, _05452_);
  and (_05455_, _04266_, _00593_);
  nor (_05456_, _04266_, _00593_);
  nor (_05457_, _05456_, _05455_);
  and (_05458_, _05457_, _05454_);
  nor (_05459_, _04283_, _00613_);
  and (_05460_, _04283_, _00613_);
  nor (_05461_, _05460_, _05459_);
  and (_05462_, _04279_, _00608_);
  nor (_05463_, _04279_, _00608_);
  or (_05464_, _05463_, _05462_);
  not (_05465_, _05464_);
  and (_05466_, _05465_, _05461_);
  and (_05467_, _05466_, _05458_);
  nor (_05468_, _04238_, _00547_);
  and (_05469_, _04238_, _00547_);
  nor (_05470_, _05469_, _05468_);
  nor (_05471_, _04230_, _00533_);
  and (_05472_, _04230_, _00533_);
  or (_05473_, _05472_, _05471_);
  not (_05474_, _05473_);
  and (_05475_, _05474_, _05470_);
  nor (_05476_, _04250_, _00569_);
  and (_05477_, _04250_, _00569_);
  nor (_05478_, _05477_, _05476_);
  nor (_05479_, _04242_, _00555_);
  and (_05480_, _04242_, _00555_);
  nor (_05481_, _05480_, _05479_);
  and (_05482_, _05481_, _05478_);
  and (_05483_, _05482_, _05475_);
  and (_05484_, _05483_, _05467_);
  and (_05485_, _05484_, _05451_);
  and (_05486_, _05485_, _05419_);
  or (_05487_, _05486_, _11613_);
  nand (_05488_, _05487_, eq_state_1);
  nor (_05489_, _05488_, _05388_);
  or (_00000_, _05489_, rst);
  and (_00008_, _05306_, _12493_);
  or (_05490_, _02518_, _02487_);
  not (_05491_, _02615_);
  nand (_05492_, _02454_, _02422_);
  or (_05493_, _05492_, _02583_);
  or (_05494_, _05493_, _02552_);
  or (_05495_, _05494_, _05491_);
  or (_05496_, _02615_, _02584_);
  or (_05497_, _05496_, _05492_);
  and (_05498_, _05497_, _05495_);
  or (_05499_, _05498_, _05490_);
  nand (_05500_, _05491_, _02519_);
  or (_05501_, _05500_, _05494_);
  and (_05502_, _05501_, _05499_);
  or (_05503_, _05502_, _02646_);
  or (_05504_, _05494_, _05490_);
  or (_05505_, _02518_, _02486_);
  or (_05506_, _05505_, _05493_);
  nand (_05507_, _05506_, _05504_);
  nand (_05508_, _05507_, _02647_);
  nand (_05509_, _02646_, _05491_);
  nand (_05510_, _02583_, _02551_);
  not (_05511_, _02454_);
  or (_05512_, _02583_, _05511_);
  and (_05513_, _05512_, _05510_);
  or (_05514_, _05505_, _02423_);
  or (_05515_, _05514_, _05513_);
  and (_05516_, _05515_, _05504_);
  or (_05517_, _05516_, _05509_);
  or (_05518_, _02647_, _02487_);
  or (_05519_, _05510_, _05492_);
  nor (_05520_, _02615_, _02518_);
  or (_05521_, _05520_, _05519_);
  or (_05522_, _05521_, _05518_);
  and (_05523_, _05522_, op0_cnst);
  and (_05524_, _05523_, _05517_);
  and (_05525_, _05524_, _05508_);
  and (_05526_, _05525_, _05503_);
  or (_00003_, _05526_, rst);
  and (_00009_, _02649_, _12493_);
  and (_00007_[7], _00959_, _12493_);
  and (_00006_[7], _00762_, _12493_);
  and (_00005_[7], _00881_, _12493_);
  and (_00004_[7], _01050_, _12493_);
  and (_05527_, _11613_, xram_data_in_reg[7]);
  and (_05528_, _11609_, xram_data_in[7]);
  or (_05529_, _05528_, _05527_);
  and (_00010_[7], _05529_, _12493_);
  not (_05530_, _05419_);
  and (_05531_, _02649_, eq_state_1);
  and (_05532_, _05531_, _05526_);
  and (_05533_, _05532_, _05324_);
  and (_05534_, _05533_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (property_invalid_xram_data_out, _05534_, _05530_);
  not (_05535_, _05485_);
  and (property_invalid_xram_addr, _05534_, _05535_);
  and (_05536_, inst_finished_r, eq_state_2);
  and (_05537_, _05536_, this_op_cnst_r);
  and (_05538_, _05537_, _05526_);
  and (_05539_, _05538_, _05489_);
  nand (_05540_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_05541_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_05542_, _05541_, _05540_);
  and (_05543_, _04181_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_05544_, \oc8051_golden_model_1.PSW [1], _08227_);
  or (_05545_, _05544_, _05543_);
  or (_05546_, _05545_, _05542_);
  and (_05547_, _04192_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_05548_, \oc8051_golden_model_1.PSW [4], _08283_);
  or (_05549_, _05548_, _05547_);
  and (_05550_, _04188_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_05551_, \oc8051_golden_model_1.PSW [3], _08881_);
  or (_05552_, _05551_, _05550_);
  or (_05553_, _05552_, _05549_);
  or (_05554_, _05553_, _05546_);
  and (_05555_, _02706_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_05556_, \oc8051_golden_model_1.PSW [7], _08218_);
  or (_05557_, _05556_, _05555_);
  and (_05558_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_05559_, _04196_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_05560_, _05559_, _05558_);
  nand (_05561_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_05562_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_05563_, _05562_, _05561_);
  or (_05564_, _05563_, _05560_);
  or (_05565_, _05564_, _05557_);
  nor (_05566_, _05565_, _05554_);
  nor (_05567_, _05566_, property_valid_psw_1_r);
  and (property_invalid_psw, _05567_, _05539_);
  not (_05568_, _05224_);
  and (property_invalid_p3, _05539_, _05568_);
  not (_05569_, _05161_);
  and (property_invalid_p2, _05539_, _05569_);
  not (_05570_, _05255_);
  and (property_invalid_p1, _05539_, _05570_);
  not (_05571_, _05192_);
  and (property_invalid_p0, _05539_, _05571_);
  not (_05572_, _05003_);
  and (property_invalid_iram, _05539_, _05572_);
  not (_05573_, _05097_);
  and (property_invalid_dph, _05539_, _05573_);
  not (_05574_, _05034_);
  and (property_invalid_dpl, _05539_, _05574_);
  not (_05575_, _05128_);
  and (property_invalid_b_reg, _05539_, _05575_);
  not (_05576_, _05065_);
  and (property_invalid_acc, _05539_, _05576_);
  and (property_invalid_pc, _05533_, _05388_);
  buf (_12544_, _12493_);
  buf (_12595_, _12493_);
  buf (_00048_, _12493_);
  buf (_00099_, _12493_);
  buf (_00151_, _12493_);
  buf (_00201_, _12493_);
  buf (_00248_, _12493_);
  buf (_00296_, _12493_);
  buf (_00336_, _12493_);
  buf (_00376_, _12493_);
  buf (_00418_, _12493_);
  buf (_00460_, _12493_);
  buf (_00504_, _12493_);
  buf (_00550_, _12493_);
  buf (_12611_, _12493_);
  buf (_12698_[7], _12676_[7]);
  buf (_12699_[7], _12677_[7]);
  buf (_12710_[7], _12676_[7]);
  buf (_12711_[7], _12677_[7]);
  buf (_12698_[0], _12676_[0]);
  buf (_12698_[1], _12676_[1]);
  buf (_12698_[2], _12676_[2]);
  buf (_12698_[3], _12676_[3]);
  buf (_12698_[4], _12676_[4]);
  buf (_12698_[5], _12676_[5]);
  buf (_12698_[6], _12676_[6]);
  buf (_12699_[0], _12677_[0]);
  buf (_12699_[1], _12677_[1]);
  buf (_12699_[2], _12677_[2]);
  buf (_12699_[3], _12677_[3]);
  buf (_12699_[4], _12677_[4]);
  buf (_12699_[5], _12677_[5]);
  buf (_12699_[6], _12677_[6]);
  buf (_12710_[0], _12676_[0]);
  buf (_12710_[1], _12676_[1]);
  buf (_12710_[2], _12676_[2]);
  buf (_12710_[3], _12676_[3]);
  buf (_12710_[4], _12676_[4]);
  buf (_12710_[5], _12676_[5]);
  buf (_12710_[6], _12676_[6]);
  buf (_12711_[0], _12677_[0]);
  buf (_12711_[1], _12677_[1]);
  buf (_12711_[2], _12677_[2]);
  buf (_12711_[3], _12677_[3]);
  buf (_12711_[4], _12677_[4]);
  buf (_12711_[5], _12677_[5]);
  buf (_12711_[6], _12677_[6]);
  buf (_12735_, _12691_);
  buf (_12730_, _12691_);
  dff (xram_data_in_reg[0], _00010_[0]);
  dff (xram_data_in_reg[1], _00010_[1]);
  dff (xram_data_in_reg[2], _00010_[2]);
  dff (xram_data_in_reg[3], _00010_[3]);
  dff (xram_data_in_reg[4], _00010_[4]);
  dff (xram_data_in_reg[5], _00010_[5]);
  dff (xram_data_in_reg[6], _00010_[6]);
  dff (xram_data_in_reg[7], _00010_[7]);
  dff (p0in_reg[0], _00004_[0]);
  dff (p0in_reg[1], _00004_[1]);
  dff (p0in_reg[2], _00004_[2]);
  dff (p0in_reg[3], _00004_[3]);
  dff (p0in_reg[4], _00004_[4]);
  dff (p0in_reg[5], _00004_[5]);
  dff (p0in_reg[6], _00004_[6]);
  dff (p0in_reg[7], _00004_[7]);
  dff (p1in_reg[0], _00005_[0]);
  dff (p1in_reg[1], _00005_[1]);
  dff (p1in_reg[2], _00005_[2]);
  dff (p1in_reg[3], _00005_[3]);
  dff (p1in_reg[4], _00005_[4]);
  dff (p1in_reg[5], _00005_[5]);
  dff (p1in_reg[6], _00005_[6]);
  dff (p1in_reg[7], _00005_[7]);
  dff (p2in_reg[0], _00006_[0]);
  dff (p2in_reg[1], _00006_[1]);
  dff (p2in_reg[2], _00006_[2]);
  dff (p2in_reg[3], _00006_[3]);
  dff (p2in_reg[4], _00006_[4]);
  dff (p2in_reg[5], _00006_[5]);
  dff (p2in_reg[6], _00006_[6]);
  dff (p2in_reg[7], _00006_[7]);
  dff (p3in_reg[0], _00007_[0]);
  dff (p3in_reg[1], _00007_[1]);
  dff (p3in_reg[2], _00007_[2]);
  dff (p3in_reg[3], _00007_[3]);
  dff (p3in_reg[4], _00007_[4]);
  dff (p3in_reg[5], _00007_[5]);
  dff (p3in_reg[6], _00007_[6]);
  dff (p3in_reg[7], _00007_[7]);
  dff (inst_finished_r, _00002_);
  dff (this_op_cnst_r, _00009_);
  dff (op0_cnst, _00003_);
  dff (property_valid_psw_1_r, _00008_);
  dff (eq_state_1, _00000_);
  dff (eq_state_2, _00001_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _12497_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _12501_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _12504_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _12508_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _12512_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _12516_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _12520_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _12490_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _12493_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _12548_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _12551_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _12555_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _12559_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _12563_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _12567_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _12571_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _12541_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _12544_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00379_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00383_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00386_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00389_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00392_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00396_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00399_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00374_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00376_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00421_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00425_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00428_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00431_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00434_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00438_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00441_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00416_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00418_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00463_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00467_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00470_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00473_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00476_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00480_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00483_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00458_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00460_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00508_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00511_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00515_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00518_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00522_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00525_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00529_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00502_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00504_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _12609_[0]);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _12609_[1]);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _12609_[2]);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _12609_[3]);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _12609_[4]);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _12609_[5]);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _12609_[6]);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _12609_[7]);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00550_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _12610_[0]);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _12610_[1]);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _12610_[2]);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _12610_[3]);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _12610_[4]);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _12610_[5]);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _12610_[6]);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _12610_[7]);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _12611_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _12599_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _12602_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _12606_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00012_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00016_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00020_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00024_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _12592_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _12595_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00052_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00056_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00060_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00064_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00067_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00071_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00075_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00045_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00048_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00103_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00107_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00111_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00115_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00119_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00123_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00127_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00096_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00099_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00155_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00158_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00162_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00166_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00170_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00174_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00178_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00148_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00151_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00204_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00208_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00212_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00215_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00219_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00222_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00226_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00198_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00201_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00252_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00256_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00259_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00263_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00266_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00270_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00274_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00245_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00248_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00299_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00303_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00307_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00310_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00314_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00318_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00319_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00293_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00296_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00339_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00342_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00346_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00349_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00352_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00356_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00359_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00333_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00336_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _12652_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _12653_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _12654_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _12655_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _12656_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _12657_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _12658_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _12659_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _12644_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _12645_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _12646_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _12647_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _12648_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _12649_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _12650_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _12651_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _12671_[0]);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _12671_[1]);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _12671_[2]);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _12671_[3]);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _12671_[4]);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _12671_[5]);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _12671_[6]);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _12671_[7]);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _12670_[0]);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _12670_[1]);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _12670_[2]);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _12670_[3]);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _12670_[4]);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _12670_[5]);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _12670_[6]);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _12670_[7]);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _12669_[0]);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _12669_[1]);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _12669_[2]);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _12669_[3]);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _12669_[4]);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _12669_[5]);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _12669_[6]);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _12669_[7]);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _12660_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _12661_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _12668_[2]);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _12668_[3]);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _12668_[4]);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _12668_[5]);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _12668_[6]);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _12668_[7]);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _12636_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _12637_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _12638_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _12639_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _12640_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _12641_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _12642_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _12643_);
  dff (\oc8051_golden_model_1.B [0], _12613_[0]);
  dff (\oc8051_golden_model_1.B [1], _12613_[1]);
  dff (\oc8051_golden_model_1.B [2], _12613_[2]);
  dff (\oc8051_golden_model_1.B [3], _12613_[3]);
  dff (\oc8051_golden_model_1.B [4], _12613_[4]);
  dff (\oc8051_golden_model_1.B [5], _12613_[5]);
  dff (\oc8051_golden_model_1.B [6], _12613_[6]);
  dff (\oc8051_golden_model_1.B [7], _12613_[7]);
  dff (\oc8051_golden_model_1.ACC [0], _12612_[0]);
  dff (\oc8051_golden_model_1.ACC [1], _12612_[1]);
  dff (\oc8051_golden_model_1.ACC [2], _12612_[2]);
  dff (\oc8051_golden_model_1.ACC [3], _12612_[3]);
  dff (\oc8051_golden_model_1.ACC [4], _12612_[4]);
  dff (\oc8051_golden_model_1.ACC [5], _12612_[5]);
  dff (\oc8051_golden_model_1.ACC [6], _12612_[6]);
  dff (\oc8051_golden_model_1.ACC [7], _12612_[7]);
  dff (\oc8051_golden_model_1.DPL [0], _12615_[0]);
  dff (\oc8051_golden_model_1.DPL [1], _12615_[1]);
  dff (\oc8051_golden_model_1.DPL [2], _12615_[2]);
  dff (\oc8051_golden_model_1.DPL [3], _12615_[3]);
  dff (\oc8051_golden_model_1.DPL [4], _12615_[4]);
  dff (\oc8051_golden_model_1.DPL [5], _12615_[5]);
  dff (\oc8051_golden_model_1.DPL [6], _12615_[6]);
  dff (\oc8051_golden_model_1.DPL [7], _12615_[7]);
  dff (\oc8051_golden_model_1.DPH [0], _12614_[0]);
  dff (\oc8051_golden_model_1.DPH [1], _12614_[1]);
  dff (\oc8051_golden_model_1.DPH [2], _12614_[2]);
  dff (\oc8051_golden_model_1.DPH [3], _12614_[3]);
  dff (\oc8051_golden_model_1.DPH [4], _12614_[4]);
  dff (\oc8051_golden_model_1.DPH [5], _12614_[5]);
  dff (\oc8051_golden_model_1.DPH [6], _12614_[6]);
  dff (\oc8051_golden_model_1.DPH [7], _12614_[7]);
  dff (\oc8051_golden_model_1.IE [0], _12616_[0]);
  dff (\oc8051_golden_model_1.IE [1], _12616_[1]);
  dff (\oc8051_golden_model_1.IE [2], _12616_[2]);
  dff (\oc8051_golden_model_1.IE [3], _12616_[3]);
  dff (\oc8051_golden_model_1.IE [4], _12616_[4]);
  dff (\oc8051_golden_model_1.IE [5], _12616_[5]);
  dff (\oc8051_golden_model_1.IE [6], _12616_[6]);
  dff (\oc8051_golden_model_1.IE [7], _12616_[7]);
  dff (\oc8051_golden_model_1.IP [0], _12617_[0]);
  dff (\oc8051_golden_model_1.IP [1], _12617_[1]);
  dff (\oc8051_golden_model_1.IP [2], _12617_[2]);
  dff (\oc8051_golden_model_1.IP [3], _12617_[3]);
  dff (\oc8051_golden_model_1.IP [4], _12617_[4]);
  dff (\oc8051_golden_model_1.IP [5], _12617_[5]);
  dff (\oc8051_golden_model_1.IP [6], _12617_[6]);
  dff (\oc8051_golden_model_1.IP [7], _12617_[7]);
  dff (\oc8051_golden_model_1.P0 [0], _12618_[0]);
  dff (\oc8051_golden_model_1.P0 [1], _12618_[1]);
  dff (\oc8051_golden_model_1.P0 [2], _12618_[2]);
  dff (\oc8051_golden_model_1.P0 [3], _12618_[3]);
  dff (\oc8051_golden_model_1.P0 [4], _12618_[4]);
  dff (\oc8051_golden_model_1.P0 [5], _12618_[5]);
  dff (\oc8051_golden_model_1.P0 [6], _12618_[6]);
  dff (\oc8051_golden_model_1.P0 [7], _12618_[7]);
  dff (\oc8051_golden_model_1.P1 [0], _12619_[0]);
  dff (\oc8051_golden_model_1.P1 [1], _12619_[1]);
  dff (\oc8051_golden_model_1.P1 [2], _12619_[2]);
  dff (\oc8051_golden_model_1.P1 [3], _12619_[3]);
  dff (\oc8051_golden_model_1.P1 [4], _12619_[4]);
  dff (\oc8051_golden_model_1.P1 [5], _12619_[5]);
  dff (\oc8051_golden_model_1.P1 [6], _12619_[6]);
  dff (\oc8051_golden_model_1.P1 [7], _12619_[7]);
  dff (\oc8051_golden_model_1.P2 [0], _12620_[0]);
  dff (\oc8051_golden_model_1.P2 [1], _12620_[1]);
  dff (\oc8051_golden_model_1.P2 [2], _12620_[2]);
  dff (\oc8051_golden_model_1.P2 [3], _12620_[3]);
  dff (\oc8051_golden_model_1.P2 [4], _12620_[4]);
  dff (\oc8051_golden_model_1.P2 [5], _12620_[5]);
  dff (\oc8051_golden_model_1.P2 [6], _12620_[6]);
  dff (\oc8051_golden_model_1.P2 [7], _12620_[7]);
  dff (\oc8051_golden_model_1.P3 [0], _12621_[0]);
  dff (\oc8051_golden_model_1.P3 [1], _12621_[1]);
  dff (\oc8051_golden_model_1.P3 [2], _12621_[2]);
  dff (\oc8051_golden_model_1.P3 [3], _12621_[3]);
  dff (\oc8051_golden_model_1.P3 [4], _12621_[4]);
  dff (\oc8051_golden_model_1.P3 [5], _12621_[5]);
  dff (\oc8051_golden_model_1.P3 [6], _12621_[6]);
  dff (\oc8051_golden_model_1.P3 [7], _12621_[7]);
  dff (\oc8051_golden_model_1.PSW [0], _12624_[0]);
  dff (\oc8051_golden_model_1.PSW [1], _12624_[1]);
  dff (\oc8051_golden_model_1.PSW [2], _12624_[2]);
  dff (\oc8051_golden_model_1.PSW [3], _12624_[3]);
  dff (\oc8051_golden_model_1.PSW [4], _12624_[4]);
  dff (\oc8051_golden_model_1.PSW [5], _12624_[5]);
  dff (\oc8051_golden_model_1.PSW [6], _12624_[6]);
  dff (\oc8051_golden_model_1.PSW [7], _12624_[7]);
  dff (\oc8051_golden_model_1.PCON [0], _12622_[0]);
  dff (\oc8051_golden_model_1.PCON [1], _12622_[1]);
  dff (\oc8051_golden_model_1.PCON [2], _12622_[2]);
  dff (\oc8051_golden_model_1.PCON [3], _12622_[3]);
  dff (\oc8051_golden_model_1.PCON [4], _12622_[4]);
  dff (\oc8051_golden_model_1.PCON [5], _12622_[5]);
  dff (\oc8051_golden_model_1.PCON [6], _12622_[6]);
  dff (\oc8051_golden_model_1.PCON [7], _12622_[7]);
  dff (\oc8051_golden_model_1.SBUF [0], _12625_[0]);
  dff (\oc8051_golden_model_1.SBUF [1], _12625_[1]);
  dff (\oc8051_golden_model_1.SBUF [2], _12625_[2]);
  dff (\oc8051_golden_model_1.SBUF [3], _12625_[3]);
  dff (\oc8051_golden_model_1.SBUF [4], _12625_[4]);
  dff (\oc8051_golden_model_1.SBUF [5], _12625_[5]);
  dff (\oc8051_golden_model_1.SBUF [6], _12625_[6]);
  dff (\oc8051_golden_model_1.SBUF [7], _12625_[7]);
  dff (\oc8051_golden_model_1.SCON [0], _12626_[0]);
  dff (\oc8051_golden_model_1.SCON [1], _12626_[1]);
  dff (\oc8051_golden_model_1.SCON [2], _12626_[2]);
  dff (\oc8051_golden_model_1.SCON [3], _12626_[3]);
  dff (\oc8051_golden_model_1.SCON [4], _12626_[4]);
  dff (\oc8051_golden_model_1.SCON [5], _12626_[5]);
  dff (\oc8051_golden_model_1.SCON [6], _12626_[6]);
  dff (\oc8051_golden_model_1.SCON [7], _12626_[7]);
  dff (\oc8051_golden_model_1.SP [0], _12627_[0]);
  dff (\oc8051_golden_model_1.SP [1], _12627_[1]);
  dff (\oc8051_golden_model_1.SP [2], _12627_[2]);
  dff (\oc8051_golden_model_1.SP [3], _12627_[3]);
  dff (\oc8051_golden_model_1.SP [4], _12627_[4]);
  dff (\oc8051_golden_model_1.SP [5], _12627_[5]);
  dff (\oc8051_golden_model_1.SP [6], _12627_[6]);
  dff (\oc8051_golden_model_1.SP [7], _12627_[7]);
  dff (\oc8051_golden_model_1.TCON [0], _12628_[0]);
  dff (\oc8051_golden_model_1.TCON [1], _12628_[1]);
  dff (\oc8051_golden_model_1.TCON [2], _12628_[2]);
  dff (\oc8051_golden_model_1.TCON [3], _12628_[3]);
  dff (\oc8051_golden_model_1.TCON [4], _12628_[4]);
  dff (\oc8051_golden_model_1.TCON [5], _12628_[5]);
  dff (\oc8051_golden_model_1.TCON [6], _12628_[6]);
  dff (\oc8051_golden_model_1.TCON [7], _12628_[7]);
  dff (\oc8051_golden_model_1.TH0 [0], _12629_[0]);
  dff (\oc8051_golden_model_1.TH0 [1], _12629_[1]);
  dff (\oc8051_golden_model_1.TH0 [2], _12629_[2]);
  dff (\oc8051_golden_model_1.TH0 [3], _12629_[3]);
  dff (\oc8051_golden_model_1.TH0 [4], _12629_[4]);
  dff (\oc8051_golden_model_1.TH0 [5], _12629_[5]);
  dff (\oc8051_golden_model_1.TH0 [6], _12629_[6]);
  dff (\oc8051_golden_model_1.TH0 [7], _12629_[7]);
  dff (\oc8051_golden_model_1.TH1 [0], _12630_[0]);
  dff (\oc8051_golden_model_1.TH1 [1], _12630_[1]);
  dff (\oc8051_golden_model_1.TH1 [2], _12630_[2]);
  dff (\oc8051_golden_model_1.TH1 [3], _12630_[3]);
  dff (\oc8051_golden_model_1.TH1 [4], _12630_[4]);
  dff (\oc8051_golden_model_1.TH1 [5], _12630_[5]);
  dff (\oc8051_golden_model_1.TH1 [6], _12630_[6]);
  dff (\oc8051_golden_model_1.TH1 [7], _12630_[7]);
  dff (\oc8051_golden_model_1.TL0 [0], _12631_[0]);
  dff (\oc8051_golden_model_1.TL0 [1], _12631_[1]);
  dff (\oc8051_golden_model_1.TL0 [2], _12631_[2]);
  dff (\oc8051_golden_model_1.TL0 [3], _12631_[3]);
  dff (\oc8051_golden_model_1.TL0 [4], _12631_[4]);
  dff (\oc8051_golden_model_1.TL0 [5], _12631_[5]);
  dff (\oc8051_golden_model_1.TL0 [6], _12631_[6]);
  dff (\oc8051_golden_model_1.TL0 [7], _12631_[7]);
  dff (\oc8051_golden_model_1.TL1 [0], _12632_[0]);
  dff (\oc8051_golden_model_1.TL1 [1], _12632_[1]);
  dff (\oc8051_golden_model_1.TL1 [2], _12632_[2]);
  dff (\oc8051_golden_model_1.TL1 [3], _12632_[3]);
  dff (\oc8051_golden_model_1.TL1 [4], _12632_[4]);
  dff (\oc8051_golden_model_1.TL1 [5], _12632_[5]);
  dff (\oc8051_golden_model_1.TL1 [6], _12632_[6]);
  dff (\oc8051_golden_model_1.TL1 [7], _12632_[7]);
  dff (\oc8051_golden_model_1.TMOD [0], _12633_[0]);
  dff (\oc8051_golden_model_1.TMOD [1], _12633_[1]);
  dff (\oc8051_golden_model_1.TMOD [2], _12633_[2]);
  dff (\oc8051_golden_model_1.TMOD [3], _12633_[3]);
  dff (\oc8051_golden_model_1.TMOD [4], _12633_[4]);
  dff (\oc8051_golden_model_1.TMOD [5], _12633_[5]);
  dff (\oc8051_golden_model_1.TMOD [6], _12633_[6]);
  dff (\oc8051_golden_model_1.TMOD [7], _12633_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [0], _12634_[0]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [1], _12634_[1]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [2], _12634_[2]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [3], _12634_[3]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [4], _12634_[4]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [5], _12634_[5]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [6], _12634_[6]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [7], _12634_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [8], _12634_[8]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [9], _12634_[9]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [10], _12634_[10]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [11], _12634_[11]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [12], _12634_[12]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [13], _12634_[13]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [14], _12634_[14]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [15], _12634_[15]);
  dff (\oc8051_golden_model_1.PC [0], _12623_[0]);
  dff (\oc8051_golden_model_1.PC [1], _12623_[1]);
  dff (\oc8051_golden_model_1.PC [2], _12623_[2]);
  dff (\oc8051_golden_model_1.PC [3], _12623_[3]);
  dff (\oc8051_golden_model_1.PC [4], _12623_[4]);
  dff (\oc8051_golden_model_1.PC [5], _12623_[5]);
  dff (\oc8051_golden_model_1.PC [6], _12623_[6]);
  dff (\oc8051_golden_model_1.PC [7], _12623_[7]);
  dff (\oc8051_golden_model_1.PC [8], _12623_[8]);
  dff (\oc8051_golden_model_1.PC [9], _12623_[9]);
  dff (\oc8051_golden_model_1.PC [10], _12623_[10]);
  dff (\oc8051_golden_model_1.PC [11], _12623_[11]);
  dff (\oc8051_golden_model_1.PC [12], _12623_[12]);
  dff (\oc8051_golden_model_1.PC [13], _12623_[13]);
  dff (\oc8051_golden_model_1.PC [14], _12623_[14]);
  dff (\oc8051_golden_model_1.PC [15], _12623_[15]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [0], _12635_[0]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [1], _12635_[1]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [2], _12635_[2]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [3], _12635_[3]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [4], _12635_[4]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [5], _12635_[5]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [6], _12635_[6]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [7], _12635_[7]);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _12665_[0]);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _12665_[1]);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _12665_[2]);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _12665_[3]);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _12665_[4]);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _12665_[5]);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _12665_[6]);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _12665_[7]);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _12667_[0]);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _12667_[1]);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _12667_[2]);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _12667_[3]);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _12667_[4]);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _12667_[5]);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _12667_[6]);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _12667_[7]);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _12666_[0]);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _12666_[1]);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _12666_[2]);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _12666_[3]);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _12666_[4]);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _12666_[5]);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _12666_[6]);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _12666_[7]);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _12662_[0]);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _12662_[1]);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _12662_[2]);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _12662_[3]);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _12662_[4]);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _12662_[5]);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _12662_[6]);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _12662_[7]);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _12664_[0]);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _12664_[1]);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _12664_[2]);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _12664_[3]);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _12664_[4]);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _12664_[5]);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _12664_[6]);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _12664_[7]);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _12663_[0]);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _12663_[1]);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _12663_[2]);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _12663_[3]);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _12663_[4]);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _12663_[5]);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _12663_[6]);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _12663_[7]);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _12673_[0]);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _12673_[1]);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _12673_[2]);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _12673_[3]);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _12673_[4]);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _12673_[5]);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _12673_[6]);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _12673_[7]);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _12674_[0]);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _12674_[1]);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _12674_[2]);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _12674_[3]);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _12674_[4]);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _12674_[5]);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _12674_[6]);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _12674_[7]);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _12672_[0]);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _12672_[1]);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _12672_[2]);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _12672_[3]);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _12672_[4]);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _12672_[5]);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _12672_[6]);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _12672_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02971_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02980_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02999_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _03017_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _03035_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _01047_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _03044_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _01016_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03055_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _03065_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _03074_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _03083_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _03093_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _03103_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03113_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _01068_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02732_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _06348_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02918_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _03102_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _03276_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03449_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03619_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03811_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _04009_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _04153_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04221_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04268_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04356_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04433_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04509_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04610_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04711_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _06542_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _12675_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _12675_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _12675_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _12675_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _12675_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _12675_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _12675_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _12675_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _12676_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _12676_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _12676_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _12676_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _12676_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _12676_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _12676_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _12676_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _12677_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _12677_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _12677_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _12677_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _12677_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12677_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _12677_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _12677_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12678_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12678_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _12678_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12679_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _12679_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _12679_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _12680_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _12680_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _12681_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _12681_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _12681_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _12681_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _12681_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _12681_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _12681_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _12681_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _12682_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _12683_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _12683_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _12684_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _12684_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _12685_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _12685_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _12685_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _12686_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _12686_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _12686_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _12687_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _12687_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _12688_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _12688_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _12688_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _12688_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _12689_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _12689_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _12690_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _12691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _12692_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _12692_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _12692_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _12692_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _12692_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _12692_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _12692_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _12692_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _12692_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _12692_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _12692_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _12692_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _12692_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _12692_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _12692_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _12692_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _12693_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _12693_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _12693_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _12693_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _12693_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _12693_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _12693_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _12693_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _12693_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _12693_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _12693_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _12693_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _12693_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _12693_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _12693_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _12693_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _12717_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _12717_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _12717_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _12717_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _12717_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _12717_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _12717_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _12717_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _12717_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _12717_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _12717_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _12717_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _12717_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _12717_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _12717_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _12717_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _12717_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _12717_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _12717_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _12717_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _12717_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _12717_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _12717_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _12717_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _12717_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _12717_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _12717_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _12717_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _12717_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _12717_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _12717_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _12717_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _12694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , _12695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _12696_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _12696_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _12696_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _12696_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _12696_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _12697_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _12697_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _12697_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _12697_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _12697_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _12697_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _12697_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _12697_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _12698_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _12698_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _12698_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _12698_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _12698_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _12698_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _12698_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _12698_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _12699_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _12699_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _12699_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _12699_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _12699_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _12699_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _12699_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _12699_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _12700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _12702_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _12702_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _12702_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _12702_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _12702_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _12702_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _12702_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _12702_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _12703_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _12703_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _12703_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _12703_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _12703_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12703_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _12703_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _12703_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _12703_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _12703_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12703_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _12703_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _12703_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _12703_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _12703_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _12703_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _12704_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _12704_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _12704_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _12704_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _12704_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _12704_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _12704_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _12704_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _12704_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _12704_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _12704_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _12704_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _12704_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _12704_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _12704_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _12704_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _12705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _12707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _12706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12708_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12708_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _12708_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12708_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12708_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _12708_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _12708_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _12708_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _12709_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _12709_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _12709_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _12710_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _12710_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _12710_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _12710_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _12710_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _12710_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _12710_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _12710_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _12711_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _12711_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _12711_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _12711_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _12711_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _12711_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _12711_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _12711_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _12712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _12713_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _12713_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _12713_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _12713_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _12713_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12713_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _12713_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _12713_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _12714_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _12715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _12716_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _12716_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _12716_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _12716_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _12718_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _12718_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _12718_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _12718_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _12718_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _12718_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12718_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _12718_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _12718_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _12718_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12718_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _12718_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _12718_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _12718_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _12718_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _12718_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _12718_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _12718_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _12718_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _12718_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _12718_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _12718_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _12718_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _12718_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _12718_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _12718_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _12718_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _12718_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _12718_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _12718_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _12718_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _12718_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _12719_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _12719_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _12719_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _12719_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _12719_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _12719_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _12719_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _12719_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _12720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _12721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _12722_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _12722_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _12722_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _12722_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _12722_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _12722_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _12722_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _12722_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _12722_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _12722_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _12722_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _12722_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _12722_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _12722_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _12722_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _12722_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _12723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _12724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _12725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _12726_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _12726_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _12726_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _12726_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _12726_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _12726_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _12726_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _12726_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _12726_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _12726_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _12726_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _12726_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _12726_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _12726_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _12726_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _12726_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _12727_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _12728_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _12729_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _12729_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _12729_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _12729_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _12729_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _12729_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _12729_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _12729_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _12730_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _12731_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _12731_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _12731_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _10374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _10380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _10385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _10390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _10395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _10400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _10405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _10408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _10415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _10419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _10422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _10426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _10429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _10433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _10436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _10439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _10589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _10593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _10596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _10600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _10603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _10607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _10610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _10613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _10561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _10565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _10568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _10572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _10575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _10579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _10582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _10585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _10533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _10537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _10540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _10544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _10547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _10551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _10554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _10557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _10505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _10509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _10512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _10516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _10519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _10523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _10526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _10529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _10475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _10478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _10482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _10485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _10489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _10492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _10496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _10498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _10446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _10449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _10453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _10456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _10460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _10463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _10467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _10469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _10620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _10623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _10627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _10630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _10634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _10637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _10641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _10644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _10789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _10793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _10796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _10800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _10803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _10807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _10810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _10813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _10761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _10765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _10768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _10772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _10775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _10779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _10782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _10785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _10733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _10737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _10740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _10744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _10747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _10751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _10754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _10757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _10704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _10708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _10711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _10715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _10718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _10722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _10725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _10728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _10676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _10680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _10683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _10687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _10690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _10694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _10697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _10700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _10648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _10652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _10655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _10659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _10662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _10666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _10669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _10672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _10817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _10821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _10824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _10828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _10831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _10835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _10838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _10127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _12471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _12473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _12475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _12477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _12478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _12480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _12482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _10115_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _12732_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _12733_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _12734_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _12734_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _12734_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _12734_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _12734_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _12734_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _12734_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _12734_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _12735_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _06312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _06314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _06316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _06320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _06136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _05578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _05579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _05580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _05581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _05582_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _05583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _05584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05598_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05600_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05602_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _05594_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _05604_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _05605_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _05606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _05608_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _05609_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _05595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _09974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _09976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _09978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _09980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _09982_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _09984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _09986_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _07330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _09988_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _09990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _09992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _09994_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _09995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _09997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _09999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _07333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _10001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _10003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _10005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _10007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _10009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _10011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _10013_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _07336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _10015_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _10017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _10019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _10021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _10023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _10025_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _10027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _07339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06067_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06069_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _06070_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _06074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _06076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _05620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _05585_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _05587_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _05588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _05589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _05590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _05591_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _05592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _05593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _05586_);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.dack_i , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [0], xram_data_in_reg[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [1], xram_data_in_reg[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [2], xram_data_in_reg[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [3], xram_data_in_reg[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [4], xram_data_in_reg[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [5], xram_data_in_reg[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [6], xram_data_in_reg[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ddat_i [7], xram_data_in_reg[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [0], RD_ROM_1_ABSTR_ADDR[0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [1], RD_ROM_1_ABSTR_ADDR[1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [2], RD_ROM_1_ABSTR_ADDR[2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [3], RD_ROM_1_ABSTR_ADDR[3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [4], RD_ROM_1_ABSTR_ADDR[4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [5], RD_ROM_1_ABSTR_ADDR[5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [6], RD_ROM_1_ABSTR_ADDR[6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [7], RD_ROM_1_ABSTR_ADDR[7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [8], RD_ROM_1_ABSTR_ADDR[8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [9], RD_ROM_1_ABSTR_ADDR[9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [10], RD_ROM_1_ABSTR_ADDR[10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [11], RD_ROM_1_ABSTR_ADDR[11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [12], RD_ROM_1_ABSTR_ADDR[12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [13], RD_ROM_1_ABSTR_ADDR[13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [14], RD_ROM_1_ABSTR_ADDR[14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_1 [15], RD_ROM_1_ABSTR_ADDR[15]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_2 [15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [0], RD_ROM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [1], RD_ROM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [2], RD_ROM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [3], RD_ROM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [4], RD_ROM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [5], RD_ROM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [6], RD_ROM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [7], RD_ROM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [8], RD_ROM_1_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [9], RD_ROM_1_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [10], RD_ROM_1_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [11], RD_ROM_1_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [12], RD_ROM_1_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [13], RD_ROM_1_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [14], RD_ROM_1_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ADDR [15], RD_ROM_1_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ADDR [15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.SBUF_next [0], \oc8051_golden_model_1.SBUF [0]);
  buf(\oc8051_golden_model_1.SBUF_next [1], \oc8051_golden_model_1.SBUF [1]);
  buf(\oc8051_golden_model_1.SBUF_next [2], \oc8051_golden_model_1.SBUF [2]);
  buf(\oc8051_golden_model_1.SBUF_next [3], \oc8051_golden_model_1.SBUF [3]);
  buf(\oc8051_golden_model_1.SBUF_next [4], \oc8051_golden_model_1.SBUF [4]);
  buf(\oc8051_golden_model_1.SBUF_next [5], \oc8051_golden_model_1.SBUF [5]);
  buf(\oc8051_golden_model_1.SBUF_next [6], \oc8051_golden_model_1.SBUF [6]);
  buf(\oc8051_golden_model_1.SBUF_next [7], \oc8051_golden_model_1.SBUF [7]);
  buf(\oc8051_golden_model_1.SCON_next [0], \oc8051_golden_model_1.SCON [0]);
  buf(\oc8051_golden_model_1.SCON_next [1], \oc8051_golden_model_1.SCON [1]);
  buf(\oc8051_golden_model_1.SCON_next [2], \oc8051_golden_model_1.SCON [2]);
  buf(\oc8051_golden_model_1.SCON_next [3], \oc8051_golden_model_1.SCON [3]);
  buf(\oc8051_golden_model_1.SCON_next [4], \oc8051_golden_model_1.SCON [4]);
  buf(\oc8051_golden_model_1.SCON_next [5], \oc8051_golden_model_1.SCON [5]);
  buf(\oc8051_golden_model_1.SCON_next [6], \oc8051_golden_model_1.SCON [6]);
  buf(\oc8051_golden_model_1.SCON_next [7], \oc8051_golden_model_1.SCON [7]);
  buf(\oc8051_golden_model_1.PCON_next [0], \oc8051_golden_model_1.PCON [0]);
  buf(\oc8051_golden_model_1.PCON_next [1], \oc8051_golden_model_1.PCON [1]);
  buf(\oc8051_golden_model_1.PCON_next [2], \oc8051_golden_model_1.PCON [2]);
  buf(\oc8051_golden_model_1.PCON_next [3], \oc8051_golden_model_1.PCON [3]);
  buf(\oc8051_golden_model_1.PCON_next [4], \oc8051_golden_model_1.PCON [4]);
  buf(\oc8051_golden_model_1.PCON_next [5], \oc8051_golden_model_1.PCON [5]);
  buf(\oc8051_golden_model_1.PCON_next [6], \oc8051_golden_model_1.PCON [6]);
  buf(\oc8051_golden_model_1.PCON_next [7], \oc8051_golden_model_1.PCON [7]);
  buf(\oc8051_golden_model_1.TCON_next [0], \oc8051_golden_model_1.TCON [0]);
  buf(\oc8051_golden_model_1.TCON_next [1], \oc8051_golden_model_1.TCON [1]);
  buf(\oc8051_golden_model_1.TCON_next [2], \oc8051_golden_model_1.TCON [2]);
  buf(\oc8051_golden_model_1.TCON_next [3], \oc8051_golden_model_1.TCON [3]);
  buf(\oc8051_golden_model_1.TCON_next [4], \oc8051_golden_model_1.TCON [4]);
  buf(\oc8051_golden_model_1.TCON_next [5], \oc8051_golden_model_1.TCON [5]);
  buf(\oc8051_golden_model_1.TCON_next [6], \oc8051_golden_model_1.TCON [6]);
  buf(\oc8051_golden_model_1.TCON_next [7], \oc8051_golden_model_1.TCON [7]);
  buf(\oc8051_golden_model_1.TL0_next [0], \oc8051_golden_model_1.TL0 [0]);
  buf(\oc8051_golden_model_1.TL0_next [1], \oc8051_golden_model_1.TL0 [1]);
  buf(\oc8051_golden_model_1.TL0_next [2], \oc8051_golden_model_1.TL0 [2]);
  buf(\oc8051_golden_model_1.TL0_next [3], \oc8051_golden_model_1.TL0 [3]);
  buf(\oc8051_golden_model_1.TL0_next [4], \oc8051_golden_model_1.TL0 [4]);
  buf(\oc8051_golden_model_1.TL0_next [5], \oc8051_golden_model_1.TL0 [5]);
  buf(\oc8051_golden_model_1.TL0_next [6], \oc8051_golden_model_1.TL0 [6]);
  buf(\oc8051_golden_model_1.TL0_next [7], \oc8051_golden_model_1.TL0 [7]);
  buf(\oc8051_golden_model_1.TL1_next [0], \oc8051_golden_model_1.TL1 [0]);
  buf(\oc8051_golden_model_1.TL1_next [1], \oc8051_golden_model_1.TL1 [1]);
  buf(\oc8051_golden_model_1.TL1_next [2], \oc8051_golden_model_1.TL1 [2]);
  buf(\oc8051_golden_model_1.TL1_next [3], \oc8051_golden_model_1.TL1 [3]);
  buf(\oc8051_golden_model_1.TL1_next [4], \oc8051_golden_model_1.TL1 [4]);
  buf(\oc8051_golden_model_1.TL1_next [5], \oc8051_golden_model_1.TL1 [5]);
  buf(\oc8051_golden_model_1.TL1_next [6], \oc8051_golden_model_1.TL1 [6]);
  buf(\oc8051_golden_model_1.TL1_next [7], \oc8051_golden_model_1.TL1 [7]);
  buf(\oc8051_golden_model_1.TH0_next [0], \oc8051_golden_model_1.TH0 [0]);
  buf(\oc8051_golden_model_1.TH0_next [1], \oc8051_golden_model_1.TH0 [1]);
  buf(\oc8051_golden_model_1.TH0_next [2], \oc8051_golden_model_1.TH0 [2]);
  buf(\oc8051_golden_model_1.TH0_next [3], \oc8051_golden_model_1.TH0 [3]);
  buf(\oc8051_golden_model_1.TH0_next [4], \oc8051_golden_model_1.TH0 [4]);
  buf(\oc8051_golden_model_1.TH0_next [5], \oc8051_golden_model_1.TH0 [5]);
  buf(\oc8051_golden_model_1.TH0_next [6], \oc8051_golden_model_1.TH0 [6]);
  buf(\oc8051_golden_model_1.TH0_next [7], \oc8051_golden_model_1.TH0 [7]);
  buf(\oc8051_golden_model_1.TH1_next [0], \oc8051_golden_model_1.TH1 [0]);
  buf(\oc8051_golden_model_1.TH1_next [1], \oc8051_golden_model_1.TH1 [1]);
  buf(\oc8051_golden_model_1.TH1_next [2], \oc8051_golden_model_1.TH1 [2]);
  buf(\oc8051_golden_model_1.TH1_next [3], \oc8051_golden_model_1.TH1 [3]);
  buf(\oc8051_golden_model_1.TH1_next [4], \oc8051_golden_model_1.TH1 [4]);
  buf(\oc8051_golden_model_1.TH1_next [5], \oc8051_golden_model_1.TH1 [5]);
  buf(\oc8051_golden_model_1.TH1_next [6], \oc8051_golden_model_1.TH1 [6]);
  buf(\oc8051_golden_model_1.TH1_next [7], \oc8051_golden_model_1.TH1 [7]);
  buf(\oc8051_golden_model_1.TMOD_next [0], \oc8051_golden_model_1.TMOD [0]);
  buf(\oc8051_golden_model_1.TMOD_next [1], \oc8051_golden_model_1.TMOD [1]);
  buf(\oc8051_golden_model_1.TMOD_next [2], \oc8051_golden_model_1.TMOD [2]);
  buf(\oc8051_golden_model_1.TMOD_next [3], \oc8051_golden_model_1.TMOD [3]);
  buf(\oc8051_golden_model_1.TMOD_next [4], \oc8051_golden_model_1.TMOD [4]);
  buf(\oc8051_golden_model_1.TMOD_next [5], \oc8051_golden_model_1.TMOD [5]);
  buf(\oc8051_golden_model_1.TMOD_next [6], \oc8051_golden_model_1.TMOD [6]);
  buf(\oc8051_golden_model_1.TMOD_next [7], \oc8051_golden_model_1.TMOD [7]);
  buf(\oc8051_golden_model_1.IE_next [0], \oc8051_golden_model_1.IE [0]);
  buf(\oc8051_golden_model_1.IE_next [1], \oc8051_golden_model_1.IE [1]);
  buf(\oc8051_golden_model_1.IE_next [2], \oc8051_golden_model_1.IE [2]);
  buf(\oc8051_golden_model_1.IE_next [3], \oc8051_golden_model_1.IE [3]);
  buf(\oc8051_golden_model_1.IE_next [4], \oc8051_golden_model_1.IE [4]);
  buf(\oc8051_golden_model_1.IE_next [5], \oc8051_golden_model_1.IE [5]);
  buf(\oc8051_golden_model_1.IE_next [6], \oc8051_golden_model_1.IE [6]);
  buf(\oc8051_golden_model_1.IE_next [7], \oc8051_golden_model_1.IE [7]);
  buf(\oc8051_golden_model_1.IP_next [0], \oc8051_golden_model_1.IP [0]);
  buf(\oc8051_golden_model_1.IP_next [1], \oc8051_golden_model_1.IP [1]);
  buf(\oc8051_golden_model_1.IP_next [2], \oc8051_golden_model_1.IP [2]);
  buf(\oc8051_golden_model_1.IP_next [3], \oc8051_golden_model_1.IP [3]);
  buf(\oc8051_golden_model_1.IP_next [4], \oc8051_golden_model_1.IP [4]);
  buf(\oc8051_golden_model_1.IP_next [5], \oc8051_golden_model_1.IP [5]);
  buf(\oc8051_golden_model_1.IP_next [6], \oc8051_golden_model_1.IP [6]);
  buf(\oc8051_golden_model_1.IP_next [7], \oc8051_golden_model_1.IP [7]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [0], xram_data_in_reg[0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [1], xram_data_in_reg[1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [2], xram_data_in_reg[2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [3], xram_data_in_reg[3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [4], xram_data_in_reg[4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [5], xram_data_in_reg[5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [6], xram_data_in_reg[6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_IN [7], xram_data_in_reg[7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [0], RD_IRAM_0_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [1], RD_IRAM_0_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [2], RD_IRAM_0_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [3], RD_IRAM_0_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [4], RD_IRAM_0_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [5], RD_IRAM_0_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [6], RD_IRAM_0_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0_ABSTR_ADDR [7], RD_IRAM_0_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [0], RD_IRAM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [1], RD_IRAM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [2], RD_IRAM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [3], RD_IRAM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [4], RD_IRAM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [5], RD_IRAM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [6], RD_IRAM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ABSTR_ADDR [7], RD_IRAM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [0], RD_ROM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [1], RD_ROM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [2], RD_ROM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [3], RD_ROM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [4], RD_ROM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [5], RD_ROM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [6], RD_ROM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [7], RD_ROM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [8], RD_ROM_1_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [9], RD_ROM_1_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [10], RD_ROM_1_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [11], RD_ROM_1_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [12], RD_ROM_1_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [13], RD_ROM_1_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [14], RD_ROM_1_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_1_ABSTR_ADDR [15], RD_ROM_1_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(\oc8051_golden_model_1.RD_ROM_2_ABSTR_ADDR [15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(\oc8051_golden_model_1.ACC_abstr [0], ACC_abstr[0]);
  buf(\oc8051_golden_model_1.ACC_abstr [1], ACC_abstr[1]);
  buf(\oc8051_golden_model_1.ACC_abstr [2], ACC_abstr[2]);
  buf(\oc8051_golden_model_1.ACC_abstr [3], ACC_abstr[3]);
  buf(\oc8051_golden_model_1.ACC_abstr [4], ACC_abstr[4]);
  buf(\oc8051_golden_model_1.ACC_abstr [5], ACC_abstr[5]);
  buf(\oc8051_golden_model_1.ACC_abstr [6], ACC_abstr[6]);
  buf(\oc8051_golden_model_1.ACC_abstr [7], ACC_abstr[7]);
  buf(\oc8051_golden_model_1.P2_abstr [0], P2_abstr[0]);
  buf(\oc8051_golden_model_1.P2_abstr [1], P2_abstr[1]);
  buf(\oc8051_golden_model_1.P2_abstr [2], P2_abstr[2]);
  buf(\oc8051_golden_model_1.P2_abstr [3], P2_abstr[3]);
  buf(\oc8051_golden_model_1.P2_abstr [4], P2_abstr[4]);
  buf(\oc8051_golden_model_1.P2_abstr [5], P2_abstr[5]);
  buf(\oc8051_golden_model_1.P2_abstr [6], P2_abstr[6]);
  buf(\oc8051_golden_model_1.P2_abstr [7], P2_abstr[7]);
  buf(\oc8051_golden_model_1.P0_abstr [0], P0_abstr[0]);
  buf(\oc8051_golden_model_1.P0_abstr [1], P0_abstr[1]);
  buf(\oc8051_golden_model_1.P0_abstr [2], P0_abstr[2]);
  buf(\oc8051_golden_model_1.P0_abstr [3], P0_abstr[3]);
  buf(\oc8051_golden_model_1.P0_abstr [4], P0_abstr[4]);
  buf(\oc8051_golden_model_1.P0_abstr [5], P0_abstr[5]);
  buf(\oc8051_golden_model_1.P0_abstr [6], P0_abstr[6]);
  buf(\oc8051_golden_model_1.P0_abstr [7], P0_abstr[7]);
  buf(\oc8051_golden_model_1.B_abstr [0], B_abstr[0]);
  buf(\oc8051_golden_model_1.B_abstr [1], B_abstr[1]);
  buf(\oc8051_golden_model_1.B_abstr [2], B_abstr[2]);
  buf(\oc8051_golden_model_1.B_abstr [3], B_abstr[3]);
  buf(\oc8051_golden_model_1.B_abstr [4], B_abstr[4]);
  buf(\oc8051_golden_model_1.B_abstr [5], B_abstr[5]);
  buf(\oc8051_golden_model_1.B_abstr [6], B_abstr[6]);
  buf(\oc8051_golden_model_1.B_abstr [7], B_abstr[7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [0], XRAM_ADDR_abstr[0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [1], XRAM_ADDR_abstr[1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [2], XRAM_ADDR_abstr[2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [3], XRAM_ADDR_abstr[3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [4], XRAM_ADDR_abstr[4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [5], XRAM_ADDR_abstr[5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [6], XRAM_ADDR_abstr[6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [7], XRAM_ADDR_abstr[7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [8], XRAM_ADDR_abstr[8]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [9], XRAM_ADDR_abstr[9]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [10], XRAM_ADDR_abstr[10]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [11], XRAM_ADDR_abstr[11]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [12], XRAM_ADDR_abstr[12]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [13], XRAM_ADDR_abstr[13]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [14], XRAM_ADDR_abstr[14]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_abstr [15], XRAM_ADDR_abstr[15]);
  buf(\oc8051_golden_model_1.P3_abstr [0], P3_abstr[0]);
  buf(\oc8051_golden_model_1.P3_abstr [1], P3_abstr[1]);
  buf(\oc8051_golden_model_1.P3_abstr [2], P3_abstr[2]);
  buf(\oc8051_golden_model_1.P3_abstr [3], P3_abstr[3]);
  buf(\oc8051_golden_model_1.P3_abstr [4], P3_abstr[4]);
  buf(\oc8051_golden_model_1.P3_abstr [5], P3_abstr[5]);
  buf(\oc8051_golden_model_1.P3_abstr [6], P3_abstr[6]);
  buf(\oc8051_golden_model_1.P3_abstr [7], P3_abstr[7]);
  buf(\oc8051_golden_model_1.SP_abstr [0], SP_abstr[0]);
  buf(\oc8051_golden_model_1.SP_abstr [1], SP_abstr[1]);
  buf(\oc8051_golden_model_1.SP_abstr [2], SP_abstr[2]);
  buf(\oc8051_golden_model_1.SP_abstr [3], SP_abstr[3]);
  buf(\oc8051_golden_model_1.SP_abstr [4], SP_abstr[4]);
  buf(\oc8051_golden_model_1.SP_abstr [5], SP_abstr[5]);
  buf(\oc8051_golden_model_1.SP_abstr [6], SP_abstr[6]);
  buf(\oc8051_golden_model_1.SP_abstr [7], SP_abstr[7]);
  buf(\oc8051_golden_model_1.PC_abstr [0], PC_abstr[0]);
  buf(\oc8051_golden_model_1.PC_abstr [1], PC_abstr[1]);
  buf(\oc8051_golden_model_1.PC_abstr [2], PC_abstr[2]);
  buf(\oc8051_golden_model_1.PC_abstr [3], PC_abstr[3]);
  buf(\oc8051_golden_model_1.PC_abstr [4], PC_abstr[4]);
  buf(\oc8051_golden_model_1.PC_abstr [5], PC_abstr[5]);
  buf(\oc8051_golden_model_1.PC_abstr [6], PC_abstr[6]);
  buf(\oc8051_golden_model_1.PC_abstr [7], PC_abstr[7]);
  buf(\oc8051_golden_model_1.PC_abstr [8], PC_abstr[8]);
  buf(\oc8051_golden_model_1.PC_abstr [9], PC_abstr[9]);
  buf(\oc8051_golden_model_1.PC_abstr [10], PC_abstr[10]);
  buf(\oc8051_golden_model_1.PC_abstr [11], PC_abstr[11]);
  buf(\oc8051_golden_model_1.PC_abstr [12], PC_abstr[12]);
  buf(\oc8051_golden_model_1.PC_abstr [13], PC_abstr[13]);
  buf(\oc8051_golden_model_1.PC_abstr [14], PC_abstr[14]);
  buf(\oc8051_golden_model_1.PC_abstr [15], PC_abstr[15]);
  buf(\oc8051_golden_model_1.P1_abstr [0], P1_abstr[0]);
  buf(\oc8051_golden_model_1.P1_abstr [1], P1_abstr[1]);
  buf(\oc8051_golden_model_1.P1_abstr [2], P1_abstr[2]);
  buf(\oc8051_golden_model_1.P1_abstr [3], P1_abstr[3]);
  buf(\oc8051_golden_model_1.P1_abstr [4], P1_abstr[4]);
  buf(\oc8051_golden_model_1.P1_abstr [5], P1_abstr[5]);
  buf(\oc8051_golden_model_1.P1_abstr [6], P1_abstr[6]);
  buf(\oc8051_golden_model_1.P1_abstr [7], P1_abstr[7]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [0], XRAM_DATA_OUT_abstr[0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [1], XRAM_DATA_OUT_abstr[1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [2], XRAM_DATA_OUT_abstr[2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [3], XRAM_DATA_OUT_abstr[3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [4], XRAM_DATA_OUT_abstr[4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [5], XRAM_DATA_OUT_abstr[5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [6], XRAM_DATA_OUT_abstr[6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_abstr [7], XRAM_DATA_OUT_abstr[7]);
  buf(\oc8051_golden_model_1.DPL_abstr [0], DPL_abstr[0]);
  buf(\oc8051_golden_model_1.DPL_abstr [1], DPL_abstr[1]);
  buf(\oc8051_golden_model_1.DPL_abstr [2], DPL_abstr[2]);
  buf(\oc8051_golden_model_1.DPL_abstr [3], DPL_abstr[3]);
  buf(\oc8051_golden_model_1.DPL_abstr [4], DPL_abstr[4]);
  buf(\oc8051_golden_model_1.DPL_abstr [5], DPL_abstr[5]);
  buf(\oc8051_golden_model_1.DPL_abstr [6], DPL_abstr[6]);
  buf(\oc8051_golden_model_1.DPL_abstr [7], DPL_abstr[7]);
  buf(\oc8051_golden_model_1.PSW_abstr [0], PSW_abstr[0]);
  buf(\oc8051_golden_model_1.PSW_abstr [1], PSW_abstr[1]);
  buf(\oc8051_golden_model_1.PSW_abstr [2], PSW_abstr[2]);
  buf(\oc8051_golden_model_1.PSW_abstr [3], PSW_abstr[3]);
  buf(\oc8051_golden_model_1.PSW_abstr [4], PSW_abstr[4]);
  buf(\oc8051_golden_model_1.PSW_abstr [5], PSW_abstr[5]);
  buf(\oc8051_golden_model_1.PSW_abstr [6], PSW_abstr[6]);
  buf(\oc8051_golden_model_1.PSW_abstr [7], PSW_abstr[7]);
  buf(\oc8051_golden_model_1.DPH_abstr [0], DPH_abstr[0]);
  buf(\oc8051_golden_model_1.DPH_abstr [1], DPH_abstr[1]);
  buf(\oc8051_golden_model_1.DPH_abstr [2], DPH_abstr[2]);
  buf(\oc8051_golden_model_1.DPH_abstr [3], DPH_abstr[3]);
  buf(\oc8051_golden_model_1.DPH_abstr [4], DPH_abstr[4]);
  buf(\oc8051_golden_model_1.DPH_abstr [5], DPH_abstr[5]);
  buf(\oc8051_golden_model_1.DPH_abstr [6], DPH_abstr[6]);
  buf(\oc8051_golden_model_1.DPH_abstr [7], DPH_abstr[7]);
  buf(\oc8051_golden_model_1.WR_COND_ABSTR_IRAM_0 , WR_COND_ABSTR_IRAM_0);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [0], WR_ADDR_ABSTR_IRAM_0[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [1], WR_ADDR_ABSTR_IRAM_0[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [2], WR_ADDR_ABSTR_IRAM_0[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_0 [3], WR_ADDR_ABSTR_IRAM_0[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [0], WR_DATA_ABSTR_IRAM_0[0]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [1], WR_DATA_ABSTR_IRAM_0[1]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [2], WR_DATA_ABSTR_IRAM_0[2]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [3], WR_DATA_ABSTR_IRAM_0[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [4], WR_DATA_ABSTR_IRAM_0[4]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [5], WR_DATA_ABSTR_IRAM_0[5]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [6], WR_DATA_ABSTR_IRAM_0[6]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_0 [7], WR_DATA_ABSTR_IRAM_0[7]);
  buf(\oc8051_golden_model_1.WR_COND_ABSTR_IRAM_1 , WR_COND_ABSTR_IRAM_1);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [0], WR_ADDR_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [1], WR_ADDR_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [2], WR_ADDR_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_ABSTR_IRAM_1 [3], WR_ADDR_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [0], WR_DATA_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [1], WR_DATA_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [2], WR_DATA_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [3], WR_DATA_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [4], WR_DATA_ABSTR_IRAM_1[4]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [5], WR_DATA_ABSTR_IRAM_1[5]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [6], WR_DATA_ABSTR_IRAM_1[6]);
  buf(\oc8051_golden_model_1.WR_DATA_ABSTR_IRAM_1 [7], WR_DATA_ABSTR_IRAM_1[7]);
  buf(\oc8051_golden_model_1.B_49 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.B_49 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.B_49 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.B_49 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.B_49 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.B_49 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.B_49 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.B_49 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.DPH_49 [0], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.DPH_49 [1], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.DPH_49 [2], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.DPH_49 [3], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.DPH_49 [4], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.DPH_49 [5], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.DPH_49 [6], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.DPH_49 [7], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.DPL_49 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.DPL_49 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.DPL_49 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.DPL_49 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.DPL_49 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.DPL_49 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.DPL_49 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.DPL_49 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.P0_49 [0], \oc8051_golden_model_1.P0 [0]);
  buf(\oc8051_golden_model_1.P0_49 [1], \oc8051_golden_model_1.P0 [1]);
  buf(\oc8051_golden_model_1.P0_49 [2], \oc8051_golden_model_1.P0 [2]);
  buf(\oc8051_golden_model_1.P0_49 [3], \oc8051_golden_model_1.P0 [3]);
  buf(\oc8051_golden_model_1.P0_49 [4], \oc8051_golden_model_1.P0 [4]);
  buf(\oc8051_golden_model_1.P0_49 [5], \oc8051_golden_model_1.P0 [5]);
  buf(\oc8051_golden_model_1.P0_49 [6], \oc8051_golden_model_1.P0 [6]);
  buf(\oc8051_golden_model_1.P0_49 [7], \oc8051_golden_model_1.P0 [7]);
  buf(\oc8051_golden_model_1.P1_49 [0], \oc8051_golden_model_1.P1 [0]);
  buf(\oc8051_golden_model_1.P1_49 [1], \oc8051_golden_model_1.P1 [1]);
  buf(\oc8051_golden_model_1.P1_49 [2], \oc8051_golden_model_1.P1 [2]);
  buf(\oc8051_golden_model_1.P1_49 [3], \oc8051_golden_model_1.P1 [3]);
  buf(\oc8051_golden_model_1.P1_49 [4], \oc8051_golden_model_1.P1 [4]);
  buf(\oc8051_golden_model_1.P1_49 [5], \oc8051_golden_model_1.P1 [5]);
  buf(\oc8051_golden_model_1.P1_49 [6], \oc8051_golden_model_1.P1 [6]);
  buf(\oc8051_golden_model_1.P1_49 [7], \oc8051_golden_model_1.P1 [7]);
  buf(\oc8051_golden_model_1.P2_49 [0], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.P2_49 [1], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.P2_49 [2], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.P2_49 [3], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.P2_49 [4], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.P2_49 [5], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.P2_49 [6], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.P2_49 [7], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.P3_49 [0], \oc8051_golden_model_1.P3 [0]);
  buf(\oc8051_golden_model_1.P3_49 [1], \oc8051_golden_model_1.P3 [1]);
  buf(\oc8051_golden_model_1.P3_49 [2], \oc8051_golden_model_1.P3 [2]);
  buf(\oc8051_golden_model_1.P3_49 [3], \oc8051_golden_model_1.P3 [3]);
  buf(\oc8051_golden_model_1.P3_49 [4], \oc8051_golden_model_1.P3 [4]);
  buf(\oc8051_golden_model_1.P3_49 [5], \oc8051_golden_model_1.P3 [5]);
  buf(\oc8051_golden_model_1.P3_49 [6], \oc8051_golden_model_1.P3 [6]);
  buf(\oc8051_golden_model_1.P3_49 [7], \oc8051_golden_model_1.P3 [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n0185 );
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [0], RD_IRAM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [1], RD_IRAM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [2], RD_IRAM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [3], RD_IRAM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [4], RD_IRAM_1_ABSTR_ADDR[4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [5], RD_IRAM_1_ABSTR_ADDR[5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [6], RD_IRAM_1_ABSTR_ADDR[6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1_ADDR [7], RD_IRAM_1_ABSTR_ADDR[7]);
  buf(\oc8051_golden_model_1.SP_49 [0], \oc8051_golden_model_1.SP [0]);
  buf(\oc8051_golden_model_1.SP_49 [1], \oc8051_golden_model_1.SP [1]);
  buf(\oc8051_golden_model_1.SP_49 [2], \oc8051_golden_model_1.SP [2]);
  buf(\oc8051_golden_model_1.SP_49 [3], \oc8051_golden_model_1.SP [3]);
  buf(\oc8051_golden_model_1.SP_49 [4], \oc8051_golden_model_1.SP [4]);
  buf(\oc8051_golden_model_1.SP_49 [5], \oc8051_golden_model_1.SP [5]);
  buf(\oc8051_golden_model_1.SP_49 [6], \oc8051_golden_model_1.SP [6]);
  buf(\oc8051_golden_model_1.SP_49 [7], \oc8051_golden_model_1.SP [7]);
  buf(\oc8051_golden_model_1.WR_ADDR_0_IRAM [0], WR_ADDR_ABSTR_IRAM_0[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_0_IRAM [1], WR_ADDR_ABSTR_IRAM_0[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_0_IRAM [2], WR_ADDR_ABSTR_IRAM_0[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_0_IRAM [3], WR_ADDR_ABSTR_IRAM_0[3]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [0], WR_ADDR_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [1], WR_ADDR_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [2], WR_ADDR_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_ADDR_1_IRAM [3], WR_ADDR_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [0], WR_DATA_ABSTR_IRAM_0[0]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [1], WR_DATA_ABSTR_IRAM_0[1]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [2], WR_DATA_ABSTR_IRAM_0[2]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [3], WR_DATA_ABSTR_IRAM_0[3]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [4], WR_DATA_ABSTR_IRAM_0[4]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [5], WR_DATA_ABSTR_IRAM_0[5]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [6], WR_DATA_ABSTR_IRAM_0[6]);
  buf(\oc8051_golden_model_1.WR_DATA_0_IRAM [7], WR_DATA_ABSTR_IRAM_0[7]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [0], WR_DATA_ABSTR_IRAM_1[0]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [1], WR_DATA_ABSTR_IRAM_1[1]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [2], WR_DATA_ABSTR_IRAM_1[2]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [3], WR_DATA_ABSTR_IRAM_1[3]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [4], WR_DATA_ABSTR_IRAM_1[4]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [5], WR_DATA_ABSTR_IRAM_1[5]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [6], WR_DATA_ABSTR_IRAM_1[6]);
  buf(\oc8051_golden_model_1.WR_DATA_1_IRAM [7], WR_DATA_ABSTR_IRAM_1[7]);
  buf(\oc8051_golden_model_1.n0004 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0004 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0006 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0006 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0006 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0006 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0006 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0006 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0006 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0010 [0], RD_IRAM_1_ABSTR_ADDR[0]);
  buf(\oc8051_golden_model_1.n0010 [1], RD_IRAM_1_ABSTR_ADDR[1]);
  buf(\oc8051_golden_model_1.n0010 [2], RD_IRAM_1_ABSTR_ADDR[2]);
  buf(\oc8051_golden_model_1.n0010 [3], RD_IRAM_1_ABSTR_ADDR[3]);
  buf(\oc8051_golden_model_1.n0186 [0], \oc8051_golden_model_1.n0185 );
  buf(\oc8051_golden_model_1.n0186 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0186 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0186 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0186 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0186 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0186 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0186 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0237 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0237 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0237 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0237 [3], 1'b0);
  buf(\oc8051_golden_model_1.n0237 [4], 1'b0);
  buf(\oc8051_golden_model_1.n0237 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0237 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0237 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0278 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0278 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0278 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0278 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0279 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0279 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0279 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0279 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0279 [4], \oc8051_golden_model_1.n0277 [0]);
  buf(\oc8051_golden_model_1.n0279 [5], \oc8051_golden_model_1.n0277 [1]);
  buf(\oc8051_golden_model_1.n0279 [6], \oc8051_golden_model_1.n0277 [2]);
  buf(\oc8051_golden_model_1.n0279 [7], \oc8051_golden_model_1.n0277 [3]);
  buf(\oc8051_golden_model_1.n0236 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0170 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n0170 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n0170 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0170 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0170 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n0170 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n0170 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n0085 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0085 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0085 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0085 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0085 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0085 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0085 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0085 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0086 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0086 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0086 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0088 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0088 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0088 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0088 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0090 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0090 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0090 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0090 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0090 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0090 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0090 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0090 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0091 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0091 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0091 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0091 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0093 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0093 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0093 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0093 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0093 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0093 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0093 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0093 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0094 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0094 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0094 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0094 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0096 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0096 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0096 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0096 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0096 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0096 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0096 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0096 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0097 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0097 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0097 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0097 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0099 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0099 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0099 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0099 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0099 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0099 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0099 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0099 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0100 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0100 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0100 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0100 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0102 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0102 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0102 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0102 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0102 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0102 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0102 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0102 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0103 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0103 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0103 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0105 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0105 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0105 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0105 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0105 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0105 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0105 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0105 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0106 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0106 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0106 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0106 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wbd_ack_i , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.wbd_dat_i [0], xram_data_in_reg[0]);
  buf(\oc8051_top_1.wbd_dat_i [1], xram_data_in_reg[1]);
  buf(\oc8051_top_1.wbd_dat_i [2], xram_data_in_reg[2]);
  buf(\oc8051_top_1.wbd_dat_i [3], xram_data_in_reg[3]);
  buf(\oc8051_top_1.wbd_dat_i [4], xram_data_in_reg[4]);
  buf(\oc8051_top_1.wbd_dat_i [5], xram_data_in_reg[5]);
  buf(\oc8051_top_1.wbd_dat_i [6], xram_data_in_reg[6]);
  buf(\oc8051_top_1.wbd_dat_i [7], xram_data_in_reg[7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(xram_data_in_model[0], xram_data_in_reg[0]);
  buf(xram_data_in_model[1], xram_data_in_reg[1]);
  buf(xram_data_in_model[2], xram_data_in_reg[2]);
  buf(xram_data_in_model[3], xram_data_in_reg[3]);
  buf(xram_data_in_model[4], xram_data_in_reg[4]);
  buf(xram_data_in_model[5], xram_data_in_reg[5]);
  buf(xram_data_in_model[6], xram_data_in_reg[6]);
  buf(xram_data_in_model[7], xram_data_in_reg[7]);
  buf(rd_rom_2_addr[0], RD_ROM_2_ABSTR_ADDR[0]);
  buf(rd_rom_2_addr[1], RD_ROM_2_ABSTR_ADDR[1]);
  buf(rd_rom_2_addr[2], RD_ROM_2_ABSTR_ADDR[2]);
  buf(rd_rom_2_addr[3], RD_ROM_2_ABSTR_ADDR[3]);
  buf(rd_rom_2_addr[4], RD_ROM_2_ABSTR_ADDR[4]);
  buf(rd_rom_2_addr[5], RD_ROM_2_ABSTR_ADDR[5]);
  buf(rd_rom_2_addr[6], RD_ROM_2_ABSTR_ADDR[6]);
  buf(rd_rom_2_addr[7], RD_ROM_2_ABSTR_ADDR[7]);
  buf(rd_rom_2_addr[8], RD_ROM_2_ABSTR_ADDR[8]);
  buf(rd_rom_2_addr[9], RD_ROM_2_ABSTR_ADDR[9]);
  buf(rd_rom_2_addr[10], RD_ROM_2_ABSTR_ADDR[10]);
  buf(rd_rom_2_addr[11], RD_ROM_2_ABSTR_ADDR[11]);
  buf(rd_rom_2_addr[12], RD_ROM_2_ABSTR_ADDR[12]);
  buf(rd_rom_2_addr[13], RD_ROM_2_ABSTR_ADDR[13]);
  buf(rd_rom_2_addr[14], RD_ROM_2_ABSTR_ADDR[14]);
  buf(rd_rom_2_addr[15], RD_ROM_2_ABSTR_ADDR[15]);
  buf(rd_rom_1_addr[0], RD_ROM_1_ABSTR_ADDR[0]);
  buf(rd_rom_1_addr[1], RD_ROM_1_ABSTR_ADDR[1]);
  buf(rd_rom_1_addr[2], RD_ROM_1_ABSTR_ADDR[2]);
  buf(rd_rom_1_addr[3], RD_ROM_1_ABSTR_ADDR[3]);
  buf(rd_rom_1_addr[4], RD_ROM_1_ABSTR_ADDR[4]);
  buf(rd_rom_1_addr[5], RD_ROM_1_ABSTR_ADDR[5]);
  buf(rd_rom_1_addr[6], RD_ROM_1_ABSTR_ADDR[6]);
  buf(rd_rom_1_addr[7], RD_ROM_1_ABSTR_ADDR[7]);
  buf(rd_rom_1_addr[8], RD_ROM_1_ABSTR_ADDR[8]);
  buf(rd_rom_1_addr[9], RD_ROM_1_ABSTR_ADDR[9]);
  buf(rd_rom_1_addr[10], RD_ROM_1_ABSTR_ADDR[10]);
  buf(rd_rom_1_addr[11], RD_ROM_1_ABSTR_ADDR[11]);
  buf(rd_rom_1_addr[12], RD_ROM_1_ABSTR_ADDR[12]);
  buf(rd_rom_1_addr[13], RD_ROM_1_ABSTR_ADDR[13]);
  buf(rd_rom_1_addr[14], RD_ROM_1_ABSTR_ADDR[14]);
  buf(rd_rom_1_addr[15], RD_ROM_1_ABSTR_ADDR[15]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm_next[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm_next[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm_next[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm_next[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm_next[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm_next[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm_next[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm_next[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm_next[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm_next[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm_next[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm_next[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm_next[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm_next[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm_next[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm_next[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm_next[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm_next[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm_next[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm_next[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm_next[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm_next[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm_next[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm_next[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm_next[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm_next[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm_next[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm_next[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm_next[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm_next[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm_next[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm_next[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm_next[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm_next[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm_next[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm_next[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm_next[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm_next[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm_next[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm_next[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm_next[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm_next[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm_next[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm_next[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm_next[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm_next[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm_next[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm_next[7], \oc8051_golden_model_1.TCON [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm_next[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm_next[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm_next[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm_next[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm_next[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm_next[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm_next[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm_next[7], \oc8051_golden_model_1.SCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm_next[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm_next[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm_next[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm_next[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm_next[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm_next[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm_next[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm_next[7], \oc8051_golden_model_1.SBUF [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm_next[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm_next[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm_next[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm_next[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm_next[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm_next[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm_next[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm_next[7], \oc8051_golden_model_1.PCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm_next[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm_next[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm_next[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm_next[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm_next[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm_next[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm_next[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm_next[7], \oc8051_golden_model_1.IP [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm_next[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm_next[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm_next[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm_next[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm_next[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm_next[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm_next[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm_next[7], \oc8051_golden_model_1.IE [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(wbd_ack_i, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_i[0], xram_data_in_reg[0]);
  buf(wbd_dat_i[1], xram_data_in_reg[1]);
  buf(wbd_dat_i[2], xram_data_in_reg[2]);
  buf(wbd_dat_i[3], xram_data_in_reg[3]);
  buf(wbd_dat_i[4], xram_data_in_reg[4]);
  buf(wbd_dat_i[5], xram_data_in_reg[5]);
  buf(wbd_dat_i[6], xram_data_in_reg[6]);
  buf(wbd_dat_i[7], xram_data_in_reg[7]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
