
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_inc_dir_iram, property_invalid_inc_acc, property_invalid_pcp1, property_invalid_pcp2, property_invalid_pcp3, property_invalid_sjmp, property_invalid_ljmp, property_invalid_ajmp, property_invalid_jc, property_invalid_jnc);
  wire [7:0] _00000_;
  wire _00001_;
  wire _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire [15:0] _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire [7:0] _36857_;
  wire _36858_;
  wire [1:0] _36859_;
  wire [5:0] _36860_;
  wire [7:0] _36861_;
  wire [1:0] _36862_;
  wire [15:0] _36863_;
  wire [7:0] _36864_;
  wire [7:0] _36865_;
  wire [7:0] _36866_;
  wire [2:0] _36867_;
  wire [2:0] _36868_;
  wire [1:0] _36869_;
  wire [7:0] _36870_;
  wire _36871_;
  wire [1:0] _36872_;
  wire [1:0] _36873_;
  wire [2:0] _36874_;
  wire [2:0] _36875_;
  wire [1:0] _36876_;
  wire [3:0] _36877_;
  wire [1:0] _36878_;
  wire _36879_;
  wire _36880_;
  wire [7:0] _36881_;
  wire [7:0] _36882_;
  wire [7:0] _36883_;
  wire [7:0] _36884_;
  wire [7:0] _36885_;
  wire [7:0] _36886_;
  wire [7:0] _36887_;
  wire [7:0] _36888_;
  wire [15:0] _36889_;
  wire [15:0] _36890_;
  wire _36891_;
  wire [4:0] _36892_;
  wire [7:0] _36893_;
  wire [7:0] _36894_;
  wire [7:0] _36895_;
  wire _36896_;
  wire _36897_;
  wire [7:0] _36898_;
  wire [15:0] _36899_;
  wire [15:0] _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire [7:0] _36904_;
  wire [2:0] _36905_;
  wire [7:0] _36906_;
  wire [7:0] _36907_;
  wire _36908_;
  wire [7:0] _36909_;
  wire _36910_;
  wire _36911_;
  wire [3:0] _36912_;
  wire [31:0] _36913_;
  wire [31:0] _36914_;
  wire [7:0] _36915_;
  wire _36916_;
  wire _36917_;
  wire [15:0] _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire [15:0] _36922_;
  wire _36923_;
  wire _36924_;
  wire [7:0] _36925_;
  wire _36926_;
  wire [2:0] _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire [7:0] _38984_;
  wire _38985_;
  wire [3:0] _38986_;
  wire _38987_;
  wire _38988_;
  wire [7:0] _38989_;
  wire _38990_;
  wire [7:0] _38991_;
  wire [7:0] _38992_;
  wire [7:0] _38993_;
  wire [7:0] _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire [7:0] _38998_;
  wire [1:0] _38999_;
  wire _39000_;
  wire [2:0] _39001_;
  wire [2:0] _39002_;
  wire [1:0] _39003_;
  wire [1:0] _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire [3:0] _39009_;
  wire [7:0] _39010_;
  wire [7:0] _39011_;
  wire [7:0] _39012_;
  wire [7:0] _39013_;
  wire [7:0] _39014_;
  wire [7:0] _39015_;
  wire [6:0] _39016_;
  wire _39017_;
  wire [7:0] _39018_;
  wire _39019_;
  wire _39020_;
  wire [7:0] _39021_;
  wire [7:0] _39022_;
  wire _39023_;
  wire _39024_;
  wire [7:0] _39025_;
  wire [7:0] _39026_;
  wire _39027_;
  wire [7:0] _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire [7:0] _39033_;
  wire [7:0] _39034_;
  wire _39035_;
  wire [7:0] _39036_;
  wire [7:0] _39037_;
  wire _39038_;
  wire [7:0] _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire [1:0] _39046_;
  wire [3:0] _39047_;
  wire [7:0] _39048_;
  wire [11:0] _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire [3:0] _39055_;
  wire [10:0] _39056_;
  wire [7:0] _39057_;
  wire [7:0] _39058_;
  wire [7:0] acc;
  wire [7:0] acc_reg;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] iram_op1;
  wire [7:0] iram_op1_reg;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire [7:0] op1_out_r;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  wire pc_change_r;
  wire pc_inc_acc_r;
  wire pc_inc_dir_r;
  output property_invalid_ajmp;
  output property_invalid_inc_acc;
  output property_invalid_inc_dir_iram;
  output property_invalid_jc;
  output property_invalid_jnc;
  output property_invalid_ljmp;
  output property_invalid_pcp1;
  output property_invalid_pcp2;
  output property_invalid_pcp3;
  output property_invalid_sjmp;
  wire [7:0] psw;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [31:0] word_in;
  and (_33127_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33128_, _33127_);
  not (_33129_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_33130_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_33131_, _33130_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33132_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_33133_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_33134_, _33133_, _33132_);
  and (_33135_, _33130_, _33129_);
  and (_33136_, _33135_, _33134_);
  and (_33137_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_33138_, _33137_);
  not (_33139_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_33140_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_33141_, _33140_);
  not (_33142_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not (_33143_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_33144_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33145_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _33144_);
  nand (_33146_, _33145_, _33143_);
  or (_33147_, _33146_, _33142_);
  not (_33148_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_33149_, _33148_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33150_, _33149_, _33143_);
  nand (_33151_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_33152_, _33151_, _33147_);
  nor (_33153_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_33154_, _33153_, _33143_);
  nand (_33155_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_33156_, _33153_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_33157_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_33158_, _33157_, _33155_);
  and (_33159_, _33153_, _33143_);
  nand (_33160_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_33161_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_33162_, _33161_, _33143_);
  nand (_33163_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_33164_, _33163_, _33160_);
  and (_33165_, _33164_, _33158_);
  nand (_33166_, _33165_, _33152_);
  nand (_33167_, _33166_, _33141_);
  nand (_33168_, _33167_, _33139_);
  nor (_33169_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _33139_);
  nor (_33170_, _33169_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_33171_, _33170_, _33168_);
  and (_33172_, _33171_, _33138_);
  nand (_33173_, _33172_, _33136_);
  not (_33174_, _33134_);
  nor (_33175_, _33135_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_33176_, _33175_, _33174_);
  and (_33177_, _33176_, _33173_);
  and (_33178_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_33179_, _33178_);
  nand (_33180_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_33181_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_33182_, _33181_, _33180_);
  nand (_33183_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  not (_33184_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_33185_, _33146_, _33184_);
  and (_33186_, _33185_, _33183_);
  nand (_33187_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_33188_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_33189_, _33188_, _33187_);
  and (_33190_, _33189_, _33186_);
  and (_33191_, _33190_, _33182_);
  or (_33192_, _33191_, _33140_);
  nand (_33193_, _33192_, _33139_);
  nor (_33194_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _33139_);
  nor (_33195_, _33194_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_33196_, _33195_, _33193_);
  and (_33197_, _33196_, _33179_);
  nand (_33198_, _33197_, _33136_);
  nor (_33199_, _33135_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_33200_, _33199_, _33174_);
  and (_33201_, _33200_, _33198_);
  nor (_33202_, _33201_, _33177_);
  and (_33203_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_33204_, _33203_);
  nand (_33205_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_33206_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_33207_, _33146_, _33206_);
  and (_33208_, _33207_, _33205_);
  nand (_33209_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_33210_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_33211_, _33210_, _33209_);
  nand (_33212_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand (_33213_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_33214_, _33213_, _33212_);
  and (_33215_, _33214_, _33211_);
  nand (_33216_, _33215_, _33208_);
  nand (_33217_, _33216_, _33141_);
  nand (_33218_, _33217_, _33139_);
  nor (_33219_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _33139_);
  nor (_33220_, _33219_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_33221_, _33220_, _33218_);
  and (_33222_, _33221_, _33204_);
  nand (_33223_, _33222_, _33136_);
  nor (_33224_, _33135_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_33225_, _33224_, _33174_);
  and (_33226_, _33225_, _33223_);
  not (_33227_, _33136_);
  and (_33228_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_33229_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_33230_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_33231_, _33230_, _33229_);
  or (_33232_, _33231_, _33228_);
  and (_33233_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_33234_, _33233_, _33140_);
  and (_33235_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_33236_, _33146_);
  and (_33237_, _33236_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_33238_, _33237_, _33235_);
  or (_33239_, _33238_, _33234_);
  or (_33240_, _33239_, _33232_);
  or (_33241_, _33240_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_33242_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _33139_);
  nor (_33243_, _33242_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_33244_, _33243_, _33241_);
  and (_33245_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_33246_, _33245_, _33244_);
  or (_33247_, _33246_, _33227_);
  nor (_33248_, _33135_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_33249_, _33248_, _33174_);
  and (_33250_, _33249_, _33247_);
  nor (_33251_, _33250_, _33226_);
  and (_33252_, _33251_, _33202_);
  nand (_33253_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nand (_33254_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_33255_, _33254_, _33253_);
  not (_33256_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_33257_, _33146_, _33256_);
  and (_33258_, _33141_, _33257_);
  and (_33259_, _33258_, _33255_);
  nand (_33260_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nand (_33261_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand (_33262_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_33263_, _33262_, _33261_);
  and (_33264_, _33263_, _33260_);
  nand (_33265_, _33264_, _33259_);
  or (_33266_, _33265_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_33267_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _33139_);
  nor (_33268_, _33267_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_33269_, _33268_, _33266_);
  and (_33270_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_33271_, _33270_, _33269_);
  or (_33272_, _33271_, _33227_);
  nor (_33273_, _33135_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_33274_, _33273_, _33174_);
  and (_33275_, _33274_, _33272_);
  and (_33276_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_33277_, _33276_);
  nand (_33278_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand (_33279_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_33280_, _33279_, _33278_);
  nand (_33281_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_33282_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_33283_, _33282_, _33281_);
  nand (_33284_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_33285_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_33286_, _33146_, _33285_);
  and (_33287_, _33286_, _33284_);
  and (_33288_, _33287_, _33283_);
  nand (_33289_, _33288_, _33280_);
  and (_33290_, _33289_, _33141_);
  or (_33291_, _33290_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_33292_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _33139_);
  nor (_33293_, _33292_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_33294_, _33293_, _33291_);
  and (_33295_, _33294_, _33277_);
  nand (_33296_, _33295_, _33136_);
  nor (_33297_, _33135_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_33298_, _33297_, _33174_);
  and (_33299_, _33298_, _33296_);
  and (_33300_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  not (_33301_, _33300_);
  nand (_33302_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_33303_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_33304_, _33146_, _33303_);
  and (_33305_, _33304_, _33302_);
  nand (_33306_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_33307_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_33308_, _33307_, _33306_);
  nand (_33309_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_33310_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_33311_, _33310_, _33309_);
  and (_33312_, _33311_, _33308_);
  and (_33313_, _33312_, _33305_);
  or (_33314_, _33313_, _33140_);
  nand (_33315_, _33314_, _33139_);
  nor (_33316_, _33139_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  nor (_33317_, _33316_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_33318_, _33317_, _33315_);
  and (_33319_, _33318_, _33301_);
  nand (_33320_, _33319_, _33136_);
  nor (_33321_, _33135_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_33322_, _33321_, _33174_);
  and (_33323_, _33322_, _33320_);
  not (_33324_, _33323_);
  and (_33325_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_33326_, _33325_);
  nand (_33327_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_33328_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_33329_, _33328_, _33327_);
  nand (_33330_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not (_33331_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_33332_, _33146_, _33331_);
  and (_33333_, _33332_, _33330_);
  nand (_33334_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_33335_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_33336_, _33335_, _33334_);
  and (_33337_, _33336_, _33333_);
  and (_33338_, _33337_, _33329_);
  or (_33339_, _33338_, _33140_);
  nand (_33340_, _33339_, _33139_);
  nor (_33341_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _33139_);
  nor (_33342_, _33341_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nand (_33343_, _33342_, _33340_);
  nand (_33344_, _33343_, _33326_);
  or (_33345_, _33344_, _33227_);
  nor (_33346_, _33135_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_33347_, _33346_, _33174_);
  nand (_33348_, _33347_, _33345_);
  and (_33349_, _33348_, _33324_);
  and (_33350_, _33349_, _33299_);
  and (_33351_, _33350_, _33275_);
  and (_33352_, _33351_, _33252_);
  not (_33353_, _33352_);
  not (_33354_, _33275_);
  and (_33355_, _33350_, _33354_);
  nand (_33356_, _33355_, _33252_);
  not (_33357_, _33299_);
  and (_33358_, _33349_, _33357_);
  and (_33359_, _33358_, _33275_);
  nand (_33360_, _33359_, _33252_);
  and (_33361_, _33360_, _33356_);
  and (_33362_, _33361_, _33353_);
  not (_33363_, _33362_);
  not (_33364_, _33201_);
  and (_33365_, _33364_, _33177_);
  not (_33366_, _33250_);
  and (_33367_, _33366_, _33226_);
  and (_33368_, _33367_, _33365_);
  not (_33369_, _33348_);
  and (_33370_, _33299_, _33369_);
  and (_33371_, _33370_, _33323_);
  and (_33372_, _33371_, _33354_);
  and (_33373_, _33372_, _33368_);
  and (_33374_, _33348_, _33323_);
  and (_33375_, _33374_, _33299_);
  and (_33376_, _33375_, _33275_);
  and (_33377_, _33368_, _33376_);
  or (_33378_, _33377_, _33373_);
  or (_33379_, _33378_, _33363_);
  nor (_33380_, _33299_, _33348_);
  and (_33381_, _33380_, _33324_);
  and (_33382_, _33381_, _33275_);
  or (_33383_, _33350_, _33382_);
  and (_33384_, _33383_, _33368_);
  and (_33385_, _33202_, _33250_);
  and (_33386_, _33382_, _33385_);
  and (_33387_, _33374_, _33357_);
  and (_33388_, _33387_, _33354_);
  nor (_33389_, _33177_, _33366_);
  nor (_33390_, _33201_, _33226_);
  and (_33391_, _33390_, _33389_);
  and (_33392_, _33391_, _33388_);
  or (_33393_, _33392_, _33386_);
  or (_33394_, _33393_, _33384_);
  and (_33395_, _33358_, _33354_);
  and (_33396_, _33395_, _33368_);
  and (_33397_, _33375_, _33354_);
  and (_33398_, _33365_, _33250_);
  and (_33399_, _33398_, _33397_);
  or (_33400_, _33399_, _33396_);
  or (_33401_, _33400_, _33394_);
  or (_33402_, _33401_, _33379_);
  and (_33403_, _33381_, _33354_);
  and (_33404_, _33368_, _33403_);
  and (_33405_, _33397_, _33252_);
  or (_33406_, _33405_, _33404_);
  and (_33407_, _33370_, _33324_);
  and (_33408_, _33407_, _33275_);
  and (_33409_, _33391_, _33408_);
  and (_33410_, _33385_, _33226_);
  and (_33411_, _33403_, _33410_);
  and (_33412_, _33391_, _33403_);
  or (_33413_, _33412_, _33411_);
  or (_33414_, _33413_, _33409_);
  nor (_33415_, _33414_, _33406_);
  and (_33416_, _33252_, _33376_);
  and (_33417_, _33380_, _33323_);
  and (_33418_, _33417_, _33275_);
  and (_33419_, _33418_, _33368_);
  and (_33420_, _33359_, _33368_);
  nor (_33421_, _33420_, _33419_);
  nand (_33422_, _33391_, _33376_);
  and (_33423_, _33417_, _33354_);
  nand (_33424_, _33391_, _33423_);
  and (_33425_, _33424_, _33422_);
  nand (_33426_, _33425_, _33421_);
  nor (_33427_, _33426_, _33416_);
  and (_33428_, _33427_, _33415_);
  and (_33429_, _33407_, _33354_);
  and (_33430_, _33429_, _33385_);
  and (_33431_, _33252_, _33417_);
  or (_33432_, _33431_, _33430_);
  and (_33433_, _33429_, _33368_);
  and (_33434_, _33368_, _33423_);
  or (_33435_, _33434_, _33433_);
  and (_33436_, _33388_, _33368_);
  and (_33437_, _33387_, _33275_);
  and (_33438_, _33437_, _33391_);
  or (_33439_, _33438_, _33436_);
  nor (_33440_, _33439_, _33435_);
  nand (_33441_, _33437_, _33368_);
  nand (_33442_, _33391_, _33350_);
  and (_33443_, _33201_, _33354_);
  nand (_33444_, _33443_, _33375_);
  and (_33445_, _33444_, _33442_);
  and (_33446_, _33445_, _33441_);
  nand (_33447_, _33391_, _33418_);
  nand (_33448_, _33391_, _33397_);
  and (_33449_, _33448_, _33447_);
  and (_33450_, _33449_, _33446_);
  nand (_33451_, _33450_, _33440_);
  nor (_33452_, _33451_, _33432_);
  nand (_33453_, _33452_, _33428_);
  or (_33454_, _33453_, _33402_);
  nand (_33455_, _33454_, _33131_);
  not (_33456_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_33457_, _33129_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_33458_, _33457_, _33456_);
  and (_33459_, _33252_, _33407_);
  and (_33460_, _33459_, _33458_);
  and (_33461_, _33458_, _33252_);
  and (_33462_, _33461_, _33381_);
  nor (_33463_, _33462_, _33460_);
  not (_33464_, _33226_);
  and (_33465_, _33385_, _33464_);
  and (_33466_, _33350_, _33465_);
  and (_33467_, \oc8051_top_1.oc8051_decoder1.state [0], _33129_);
  and (_33468_, _33467_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_33469_, _33468_, _33466_);
  not (_33470_, _33469_);
  and (_33471_, _33470_, _33463_);
  nand (_33472_, _33471_, _33455_);
  nand (_33473_, _33472_, _33129_);
  and (_33474_, _33473_, _33128_);
  not (_33475_, _33474_);
  and (_33476_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33477_, _33131_);
  and (_33478_, _33251_, _33365_);
  and (_33479_, _33478_, _33388_);
  and (_33480_, _33478_, _33397_);
  nor (_33481_, _33480_, _33479_);
  and (_33482_, _33437_, _33410_);
  not (_33483_, _33482_);
  nand (_33484_, _33410_, _33408_);
  nand (_33485_, _33397_, _33410_);
  and (_33486_, _33485_, _33484_);
  and (_33487_, _33486_, _33483_);
  and (_33488_, _33487_, _33481_);
  nor (_33489_, _33488_, _33477_);
  not (_33490_, _33130_);
  and (_33491_, _33480_, _33129_);
  and (_33492_, _33491_, _33490_);
  and (_33493_, _33479_, _33477_);
  nor (_33494_, _33493_, _33492_);
  and (_33495_, _33494_, _33463_);
  not (_33496_, _33495_);
  nor (_33497_, _33496_, _33489_);
  nor (_33498_, _33497_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_33499_, _33498_, _33476_);
  not (_33500_, _33499_);
  and (_33501_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_33502_, _33501_);
  and (_33503_, _33398_, _33383_);
  and (_33504_, _33398_, _33376_);
  nand (_33505_, _33398_, _33358_);
  not (_33506_, _33505_);
  and (_33507_, _33398_, _33388_);
  or (_33508_, _33507_, _33506_);
  nor (_33509_, _33508_, _33504_);
  not (_33510_, _33466_);
  nand (_33511_, _33398_, _33429_);
  and (_33512_, _33511_, _33510_);
  nand (_33513_, _33512_, _33509_);
  nor (_33514_, _33513_, _33503_);
  and (_33515_, _33398_, _33354_);
  nor (_33516_, _33371_, _33381_);
  not (_33517_, _33516_);
  nand (_33518_, _33517_, _33515_);
  nand (_33519_, _33418_, _33252_);
  nand (_33520_, _33398_, _33417_);
  not (_33521_, _33520_);
  and (_33522_, _33398_, _33437_);
  nor (_33523_, _33522_, _33521_);
  and (_33524_, _33523_, _33519_);
  and (_33525_, _33524_, _33518_);
  and (_33526_, _33525_, _33487_);
  nand (_33527_, _33526_, _33514_);
  nand (_33528_, _33527_, _33131_);
  nor (_33529_, _33469_, _33460_);
  nand (_33530_, _33529_, _33528_);
  nand (_33531_, _33530_, _33129_);
  and (_33532_, _33531_, _33502_);
  nor (_33533_, _33532_, _33500_);
  and (_33534_, _33533_, _33475_);
  not (_33535_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_33536_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _33129_);
  and (_33537_, _33536_, _33535_);
  and (_33538_, _33537_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_33539_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_33540_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_33541_, _33537_, _33540_);
  and (_33542_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_33543_, _33542_, _33539_);
  and (_33544_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _33129_);
  nor (_33545_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_33546_, _33545_, _33544_);
  and (_33547_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_33548_, _33547_);
  not (_33549_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_33550_, _33544_, _33540_);
  and (_33551_, _33550_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_33552_, _33551_, _33549_);
  and (_33553_, _33545_, _33535_);
  or (_33554_, _33553_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_33555_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_33556_, _33555_, _33552_);
  and (_33557_, _33556_, _33548_);
  and (_33558_, _33557_, _33543_);
  not (_33559_, _33558_);
  and (_33560_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_33561_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_33562_, _33561_, _33560_);
  and (_33563_, _33562_, _33551_);
  and (_33564_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_33565_, _33564_, _33563_);
  and (_33566_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_33567_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_33568_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_33569_, _33568_, _33567_);
  nor (_33570_, _33569_, _33566_);
  and (_33571_, _33570_, _33565_);
  and (_33572_, _33571_, _33559_);
  and (_33573_, _33560_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_33574_, _33573_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_33575_, _33574_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_33576_, _33575_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_33577_, _33576_);
  not (_33578_, _33551_);
  nor (_33579_, _33575_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_33580_, _33579_, _33578_);
  and (_33581_, _33580_, _33577_);
  not (_33582_, _33581_);
  and (_33583_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_33584_, _33583_, _33544_);
  and (_33585_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_33586_, _33585_, _33584_);
  and (_33587_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_33588_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_33589_, _33588_, _33587_);
  and (_33590_, _33589_, _33586_);
  and (_33591_, _33590_, _33582_);
  and (_33592_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_33593_, _33592_, _33584_);
  not (_33594_, _33575_);
  nor (_33595_, _33574_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_33596_, _33595_, _33578_);
  and (_33597_, _33596_, _33594_);
  and (_33598_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_33599_, _33598_, _33597_);
  and (_33600_, _33599_, _33593_);
  and (_33601_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_33602_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_33603_, _33602_, _33601_);
  and (_33604_, _33603_, _33600_);
  and (_33605_, _33604_, _33591_);
  and (_33606_, _33576_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or (_33607_, _33606_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_33608_, _33606_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_33609_, _33608_, _33551_);
  and (_33610_, _33609_, _33607_);
  not (_33611_, _33610_);
  and (_33612_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_33613_, _33612_, _33584_);
  and (_33614_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  and (_33615_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor (_33616_, _33615_, _33614_);
  and (_33617_, _33616_, _33613_);
  and (_33618_, _33617_, _33611_);
  not (_33619_, _33606_);
  nor (_33620_, _33576_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_33621_, _33620_, _33578_);
  and (_33622_, _33621_, _33619_);
  not (_33623_, _33622_);
  and (_33624_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_33625_, _33624_, _33584_);
  and (_33626_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_33627_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_33628_, _33627_, _33626_);
  and (_33629_, _33628_, _33625_);
  and (_33630_, _33629_, _33623_);
  not (_33631_, _33630_);
  nor (_33632_, _33631_, _33618_);
  and (_33633_, _33632_, _33605_);
  nor (_33634_, _33560_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_33635_, _33634_, _33573_);
  and (_33636_, _33635_, _33551_);
  and (_33637_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_33638_, _33637_, _33636_);
  and (_33639_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_33640_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_33641_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_33642_, _33641_, _33640_);
  nor (_33643_, _33642_, _33639_);
  and (_33644_, _33643_, _33638_);
  and (_33645_, _33538_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_33646_, _33541_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_33647_, _33646_, _33645_);
  not (_33648_, _33574_);
  nor (_33649_, _33573_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_33650_, _33649_, _33578_);
  and (_33651_, _33650_, _33648_);
  not (_33652_, _33651_);
  and (_33653_, _33554_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_33654_, _33546_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_33655_, _33654_, _33653_);
  and (_33656_, _33655_, _33652_);
  and (_33657_, _33656_, _33647_);
  not (_33658_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_33659_, \oc8051_top_1.oc8051_decoder1.wr , _33129_);
  not (_33660_, _33659_);
  nor (_33661_, _33660_, _33550_);
  and (_33662_, _33661_, _33658_);
  and (_33663_, _33662_, _33657_);
  and (_33664_, _33663_, _33644_);
  and (_33665_, _33664_, _33633_);
  and (_33666_, _33665_, _33572_);
  not (_33667_, _33666_);
  and (_33668_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_33669_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_33670_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _33129_);
  and (_33671_, _33670_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_33672_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _33129_);
  and (_33673_, _33672_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_33674_, _33673_, _33671_);
  not (_33675_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  nand (_33676_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _33675_);
  nor (_33677_, _33676_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_33678_, _33677_);
  or (_33679_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  not (_33680_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_33681_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _33680_);
  and (_33682_, _33681_, _33679_);
  not (_33683_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_33684_, _33683_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_33685_, _33684_, _33682_);
  and (_33686_, _33685_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or (_33687_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  or (_33688_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _33680_);
  and (_33689_, _33688_, _33687_);
  nor (_33690_, _33683_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_33691_, _33690_, _33689_);
  or (_33692_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or (_33693_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _33680_);
  and (_33694_, _33693_, _33692_);
  nor (_33695_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_33696_, _33695_, _33694_);
  or (_33697_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or (_33698_, _33680_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_33699_, _33698_, _33697_);
  and (_33700_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_33701_, _33700_, _33699_);
  and (_33702_, _33701_, _33696_);
  and (_33703_, _33702_, _33691_);
  nand (_33704_, _33703_, _33686_);
  not (_33705_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  or (_33706_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  or (_33707_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _33680_);
  and (_33708_, _33707_, _33706_);
  nand (_33709_, _33708_, _33684_);
  and (_33710_, _33709_, _33705_);
  or (_33711_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or (_33712_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _33680_);
  and (_33713_, _33712_, _33711_);
  nand (_33714_, _33713_, _33700_);
  or (_33715_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  or (_33716_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _33680_);
  and (_33717_, _33716_, _33715_);
  nand (_33718_, _33717_, _33695_);
  or (_33719_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or (_33720_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _33680_);
  and (_33721_, _33720_, _33719_);
  nand (_33722_, _33721_, _33690_);
  and (_33723_, _33722_, _33718_);
  and (_33724_, _33723_, _33714_);
  nand (_33725_, _33724_, _33710_);
  nand (_33726_, _33725_, _33704_);
  nand (_33727_, _33726_, _33676_);
  and (_33728_, _33727_, _33678_);
  and (_33729_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_33730_, _33729_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_33731_, _33730_);
  and (_33732_, _33731_, _33728_);
  and (_33733_, _33731_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_33734_, _33733_, _33732_);
  not (_33735_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_33736_, _33735_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_33737_, _33736_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_33738_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_33739_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_33740_, _33739_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_33741_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_33742_, _33741_, _33738_);
  nor (_33743_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_33744_, _33743_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_33745_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_33746_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_33747_, _33736_, _33746_);
  and (_33748_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_33749_, _33748_, _33745_);
  and (_33750_, _33749_, _33742_);
  and (_33751_, _33739_, _33746_);
  not (_33752_, _33751_);
  and (_33753_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _33675_);
  or (_33754_, _33682_, _33753_);
  or (_33755_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_33756_, _33755_, _33754_);
  or (_33757_, _33756_, _33752_);
  and (_33758_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_33759_, _33758_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_33760_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_33761_, _33758_, _33746_);
  and (_33762_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_33763_, _33762_, _33760_);
  and (_33764_, _33763_, _33757_);
  and (_33765_, _33764_, _33750_);
  not (_33766_, _33765_);
  and (_33767_, _33766_, _33734_);
  nor (_33768_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_33769_, _33768_);
  or (_33770_, _33769_, _33756_);
  and (_33771_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_33772_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_33773_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_33774_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_33775_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _33774_);
  nor (_33776_, _33775_, _33773_);
  nor (_33777_, _33776_, _33772_);
  and (_33778_, _33777_, _33770_);
  nor (_33779_, _33778_, _33734_);
  or (_33780_, _33779_, _33767_);
  and (_33781_, _33780_, _33674_);
  nand (_33782_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nand (_33783_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_33784_, _33783_, _33782_);
  nand (_33785_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_33786_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_33787_, _33786_, _33785_);
  and (_33788_, _33787_, _33784_);
  or (_33789_, _33689_, _33753_);
  or (_33790_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_33791_, _33790_, _33789_);
  or (_33792_, _33791_, _33752_);
  nand (_33793_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nand (_33794_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_33795_, _33794_, _33793_);
  and (_33796_, _33795_, _33792_);
  and (_33797_, _33796_, _33788_);
  not (_33798_, _33797_);
  and (_33799_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_33800_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  nor (_33801_, _33800_, _33799_);
  and (_33802_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_33803_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_33804_, _33803_, _33802_);
  and (_33805_, _33804_, _33801_);
  or (_33806_, _33713_, _33753_);
  or (_33807_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_33808_, _33807_, _33806_);
  or (_33809_, _33808_, _33752_);
  and (_33810_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_33811_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_33812_, _33811_, _33810_);
  and (_33813_, _33812_, _33809_);
  and (_33814_, _33813_, _33805_);
  not (_33815_, _33814_);
  nand (_33816_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_33817_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_33818_, _33817_, _33816_);
  nand (_33819_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand (_33820_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_33821_, _33820_, _33819_);
  and (_33822_, _33821_, _33818_);
  or (_33823_, _33721_, _33753_);
  or (_33824_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_33825_, _33824_, _33823_);
  or (_33826_, _33825_, _33752_);
  nand (_33827_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand (_33828_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_33829_, _33828_, _33827_);
  and (_33830_, _33829_, _33826_);
  and (_33831_, _33830_, _33822_);
  and (_33832_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_33833_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_33834_, _33833_, _33832_);
  and (_33835_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_33836_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_33837_, _33836_, _33835_);
  and (_33838_, _33837_, _33834_);
  or (_33839_, _33717_, _33753_);
  or (_33840_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_33841_, _33840_, _33839_);
  and (_33842_, _33841_, _33751_);
  and (_33843_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_33844_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_33845_, _33844_, _33843_);
  not (_33846_, _33845_);
  nor (_33847_, _33846_, _33842_);
  and (_33848_, _33847_, _33838_);
  nor (_33849_, _33848_, _33831_);
  nand (_33850_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand (_33851_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_33852_, _33851_, _33850_);
  nand (_33853_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_33854_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_33855_, _33854_, _33853_);
  and (_33856_, _33855_, _33852_);
  or (_33857_, _33708_, _33753_);
  or (_33858_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_33859_, _33858_, _33857_);
  or (_33860_, _33859_, _33752_);
  nand (_33861_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand (_33862_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_33863_, _33862_, _33861_);
  and (_33864_, _33863_, _33860_);
  nand (_33865_, _33864_, _33856_);
  and (_33866_, _33865_, _33849_);
  and (_33867_, _33866_, _33815_);
  and (_33868_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_33869_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_33870_, _33869_, _33868_);
  and (_33871_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_33872_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_33873_, _33872_, _33871_);
  and (_33874_, _33873_, _33870_);
  or (_33875_, _33694_, _33753_);
  or (_33876_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_33877_, _33876_, _33875_);
  or (_33878_, _33877_, _33752_);
  and (_33879_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_33880_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_33881_, _33880_, _33879_);
  and (_33882_, _33881_, _33878_);
  and (_33883_, _33882_, _33874_);
  not (_33884_, _33883_);
  and (_33885_, _33884_, _33867_);
  and (_33886_, _33885_, _33798_);
  and (_33887_, _33886_, _33734_);
  not (_33888_, _33734_);
  nand (_33889_, _33848_, _33831_);
  nor (_33890_, _33889_, _33865_);
  and (_33891_, _33890_, _33814_);
  and (_33892_, _33891_, _33883_);
  and (_33893_, _33892_, _33797_);
  and (_33894_, _33893_, _33888_);
  or (_33895_, _33894_, _33887_);
  and (_33896_, _33895_, _33766_);
  not (_33897_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_33898_, _33672_, _33897_);
  and (_33899_, _33671_, _33898_);
  or (_33900_, _33895_, _33766_);
  nand (_33901_, _33900_, _33899_);
  nor (_33902_, _33901_, _33896_);
  nor (_33903_, _33902_, _33781_);
  not (_33904_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_33905_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _33129_);
  and (_33906_, _33905_, _33904_);
  not (_33907_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_33908_, _33670_, _33907_);
  and (_33909_, _33908_, _33906_);
  not (_33910_, _33909_);
  and (_33911_, _33778_, _33765_);
  nor (_33912_, _33911_, _33910_);
  nor (_33913_, _33905_, _33672_);
  and (_33914_, _33913_, _33908_);
  nor (_33915_, _33778_, _33765_);
  nor (_33916_, _33915_, _33911_);
  and (_33917_, _33916_, _33914_);
  nor (_33918_, _33917_, _33912_);
  not (_33919_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_33920_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _33129_);
  and (_33921_, _33920_, _33919_);
  and (_33922_, _33921_, _33673_);
  and (_33923_, _33915_, _33922_);
  and (_33924_, _33921_, _33898_);
  and (_33925_, _33924_, _33765_);
  nor (_33926_, _33925_, _33923_);
  and (_33927_, _33908_, _33672_);
  not (_33928_, _33927_);
  nor (_33929_, _33928_, _33765_);
  nor (_33930_, _33670_, _33920_);
  and (_33931_, _33930_, _33905_);
  and (_33932_, _33921_, _33904_);
  nor (_33933_, _33932_, _33931_);
  and (_33934_, _33671_, _33904_);
  and (_33935_, _33930_, _33913_);
  nor (_33936_, _33935_, _33934_);
  and (_33937_, _33936_, _33933_);
  nor (_33938_, _33937_, _33765_);
  nor (_33939_, _33938_, _33929_);
  and (_33940_, _33939_, _33926_);
  and (_33941_, _33940_, _33918_);
  nand (_33942_, _33941_, _33903_);
  and (_33943_, _33942_, _33666_);
  nor (_33944_, _33943_, _33669_);
  and (_33945_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  or (_33946_, _33769_, _33791_);
  nand (_33947_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  not (_33948_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_33949_, _33775_, _33948_);
  and (_33950_, _33949_, _33947_);
  and (_33951_, _33950_, _33946_);
  nor (_33952_, _33951_, _33734_);
  and (_33953_, _33798_, _33734_);
  or (_33954_, _33953_, _33952_);
  and (_33955_, _33954_, _33674_);
  nor (_33956_, _33885_, _33888_);
  nor (_33957_, _33892_, _33734_);
  nor (_33958_, _33957_, _33956_);
  and (_33959_, _33958_, _33798_);
  or (_33960_, _33958_, _33798_);
  nand (_33961_, _33960_, _33899_);
  nor (_33962_, _33961_, _33959_);
  nor (_33963_, _33962_, _33955_);
  and (_33964_, _33951_, _33797_);
  nor (_33965_, _33964_, _33910_);
  nor (_33966_, _33951_, _33797_);
  nor (_33967_, _33966_, _33964_);
  and (_33968_, _33967_, _33914_);
  nor (_33969_, _33968_, _33965_);
  and (_33970_, _33966_, _33922_);
  and (_33971_, _33924_, _33797_);
  nor (_33972_, _33971_, _33970_);
  nor (_33973_, _33928_, _33797_);
  nor (_33974_, _33937_, _33797_);
  nor (_33975_, _33974_, _33973_);
  and (_33976_, _33975_, _33972_);
  and (_33977_, _33976_, _33969_);
  nand (_33978_, _33977_, _33963_);
  and (_33979_, _33978_, _33666_);
  nor (_33980_, _33979_, _33945_);
  and (_33981_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_33982_, _33769_, _33877_);
  nand (_33983_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not (_33984_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_33985_, _33775_, _33984_);
  and (_33986_, _33985_, _33983_);
  and (_33987_, _33986_, _33982_);
  and (_33988_, _33987_, _33883_);
  nor (_33989_, _33988_, _33910_);
  nor (_33990_, _33987_, _33883_);
  nor (_33991_, _33990_, _33988_);
  and (_33992_, _33991_, _33914_);
  nor (_33993_, _33992_, _33989_);
  nor (_33994_, _33928_, _33883_);
  nor (_33995_, _33937_, _33883_);
  nor (_33996_, _33995_, _33994_);
  and (_33997_, _33996_, _33993_);
  nand (_33998_, _33867_, _33734_);
  nand (_33999_, _33891_, _33888_);
  and (_34000_, _33999_, _33998_);
  and (_34001_, _34000_, _33883_);
  or (_34002_, _34000_, _33883_);
  nand (_34003_, _34002_, _33899_);
  or (_34004_, _34003_, _34001_);
  and (_34005_, _33883_, _33734_);
  not (_34006_, _33674_);
  nand (_34007_, _33986_, _33982_);
  nor (_34008_, _34007_, _33734_);
  or (_34009_, _34008_, _34006_);
  nor (_34010_, _34009_, _34005_);
  and (_34011_, _33990_, _33922_);
  and (_34012_, _33924_, _33883_);
  nor (_34013_, _34012_, _34011_);
  not (_34014_, _34013_);
  nor (_34015_, _34014_, _34010_);
  and (_34016_, _34015_, _34004_);
  and (_34017_, _34016_, _33997_);
  nor (_34018_, _34017_, _33667_);
  nor (_34019_, _34018_, _33981_);
  nor (_34020_, _33928_, _33814_);
  nor (_34021_, _33937_, _33814_);
  nor (_34022_, _34021_, _34020_);
  or (_34023_, _33890_, _33734_);
  or (_34024_, _33866_, _33888_);
  and (_34025_, _34024_, _34023_);
  or (_34026_, _34025_, _33814_);
  nand (_34027_, _34025_, _33814_);
  nand (_34028_, _34027_, _34026_);
  nand (_34029_, _34028_, _33899_);
  or (_34030_, _33769_, _33808_);
  nand (_34031_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  not (_34032_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_34033_, _33775_, _34032_);
  and (_34034_, _34033_, _34031_);
  and (_34035_, _34034_, _34030_);
  and (_34036_, _34035_, _33814_);
  nor (_34037_, _34036_, _33910_);
  nor (_34038_, _34035_, _33814_);
  or (_34039_, _34038_, _34036_);
  not (_34040_, _34039_);
  and (_34041_, _34040_, _33914_);
  or (_34042_, _34041_, _34037_);
  and (_34043_, _34038_, _33922_);
  not (_34044_, _34043_);
  nor (_34045_, _34035_, _34006_);
  and (_34046_, _33924_, _33814_);
  nor (_34047_, _34046_, _34045_);
  and (_34048_, _34047_, _34044_);
  not (_34049_, _34048_);
  nor (_34050_, _34049_, _34042_);
  and (_34051_, _34050_, _34029_);
  and (_34052_, _34051_, _34022_);
  nor (_34053_, _34052_, _33667_);
  and (_34054_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_34055_, _34054_, _34053_);
  and (_34056_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or (_34057_, _33769_, _33859_);
  nand (_34058_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_34059_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_34060_, _33775_, _34059_);
  and (_34061_, _34060_, _34058_);
  nand (_34062_, _34061_, _34057_);
  and (_34063_, _34062_, _33674_);
  not (_34064_, _33865_);
  not (_34065_, _33849_);
  and (_34066_, _34065_, _33734_);
  and (_34067_, _33889_, _33888_);
  nor (_34068_, _34067_, _34066_);
  nand (_34069_, _34068_, _34064_);
  or (_34070_, _34068_, _34064_);
  nand (_34071_, _34070_, _34069_);
  and (_34072_, _34071_, _33899_);
  nor (_34073_, _34072_, _34063_);
  nor (_34074_, _34062_, _33865_);
  nor (_34075_, _34074_, _33910_);
  and (_34076_, _34062_, _33865_);
  nor (_34077_, _34076_, _34074_);
  and (_34078_, _34077_, _33914_);
  nor (_34079_, _34078_, _34075_);
  and (_34080_, _34076_, _33922_);
  and (_34081_, _33924_, _34064_);
  nor (_34082_, _34081_, _34080_);
  and (_34083_, _33927_, _33865_);
  not (_34084_, _33937_);
  and (_34085_, _34084_, _33865_);
  nor (_34086_, _34085_, _34083_);
  and (_34087_, _34086_, _34082_);
  and (_34088_, _34087_, _34079_);
  nand (_34089_, _34088_, _34073_);
  and (_34090_, _34089_, _33666_);
  nor (_34091_, _34090_, _34056_);
  and (_34092_, _33667_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or (_34093_, _33769_, _33825_);
  nand (_34094_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  not (_34095_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_34096_, _33775_, _34095_);
  and (_34097_, _34096_, _34094_);
  nand (_34098_, _34097_, _34093_);
  and (_34099_, _34098_, _33674_);
  not (_34100_, _33899_);
  and (_34101_, _33889_, _34065_);
  nand (_34102_, _34101_, _33734_);
  or (_34103_, _34101_, _33734_);
  and (_34104_, _34103_, _34102_);
  nor (_34105_, _34104_, _34100_);
  nor (_34106_, _34105_, _34099_);
  not (_34107_, _34098_);
  and (_34108_, _34107_, _33831_);
  nor (_34109_, _34108_, _33910_);
  nor (_34110_, _34107_, _33831_);
  nor (_34111_, _34110_, _34108_);
  and (_34112_, _34111_, _33914_);
  nor (_34113_, _34112_, _34109_);
  and (_34114_, _34110_, _33922_);
  and (_34115_, _33924_, _33831_);
  nor (_34116_, _34115_, _34114_);
  nor (_34117_, _33928_, _33831_);
  nor (_34118_, _33937_, _33831_);
  nor (_34119_, _34118_, _34117_);
  and (_34120_, _34119_, _34116_);
  and (_34121_, _34120_, _34113_);
  nand (_34122_, _34121_, _34106_);
  and (_34123_, _34122_, _33666_);
  nor (_34124_, _34123_, _34092_);
  or (_34125_, _33666_, _33549_);
  nand (_34126_, _33768_, _33841_);
  nand (_34127_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  not (_34128_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_34129_, _33775_, _34128_);
  and (_34130_, _34129_, _34127_);
  nand (_34131_, _34130_, _34126_);
  not (_34132_, _34131_);
  and (_34133_, _34132_, _33848_);
  nor (_34134_, _34132_, _33848_);
  nor (_34135_, _34134_, _34133_);
  nand (_34136_, _34135_, _33914_);
  nand (_34137_, _34134_, _33922_);
  nor (_34138_, _34133_, _33910_);
  and (_34139_, _34131_, _33674_);
  and (_34140_, _33920_, _33898_);
  and (_34141_, _34140_, _33848_);
  or (_34142_, _34141_, _34139_);
  nor (_34143_, _34142_, _34138_);
  and (_34144_, _34143_, _34137_);
  and (_34145_, _34144_, _34136_);
  and (_34146_, _33937_, _33928_);
  or (_34147_, _34146_, _33848_);
  and (_34148_, _34147_, _34145_);
  not (_34149_, _34148_);
  nand (_34150_, _34149_, _33666_);
  and (_34151_, _34150_, _34125_);
  and (_34152_, _34151_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_34153_, _34152_, _34124_);
  and (_34154_, _34153_, _34091_);
  and (_34155_, _34154_, _34055_);
  and (_34156_, _34155_, _34019_);
  and (_34157_, _34156_, _33980_);
  and (_34158_, _34157_, _33944_);
  nand (_34159_, _34158_, _33668_);
  or (_34160_, _34158_, _33668_);
  and (_34161_, _34160_, _33578_);
  nand (_34162_, _34161_, _34159_);
  nor (_34163_, _33666_, _33610_);
  and (_34164_, _34163_, _34162_);
  and (_34165_, _33737_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_34166_, _33740_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_34167_, _34166_, _34165_);
  and (_34168_, _33744_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_34169_, _33747_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_34170_, _34169_, _34168_);
  and (_34171_, _34170_, _34167_);
  or (_34172_, _33699_, _33753_);
  or (_34173_, _33676_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_34174_, _34173_, _34172_);
  or (_34175_, _34174_, _33752_);
  and (_34176_, _33761_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_34177_, _33759_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_34178_, _34177_, _34176_);
  and (_34179_, _34178_, _34175_);
  and (_34180_, _34179_, _34171_);
  and (_34181_, _33886_, _33766_);
  nor (_34182_, _34181_, _33888_);
  and (_34183_, _33797_, _33765_);
  and (_34184_, _34183_, _33892_);
  nor (_34185_, _34184_, _33734_);
  or (_34186_, _34185_, _34182_);
  and (_34187_, _34186_, _34180_);
  nor (_34188_, _34186_, _34180_);
  nor (_34189_, _34188_, _34187_);
  and (_34190_, _34189_, _33899_);
  or (_34191_, _33769_, _34174_);
  and (_34192_, _33771_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_34193_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_34194_, _33775_, _34193_);
  nor (_34195_, _34194_, _34192_);
  and (_34196_, _34195_, _34191_);
  not (_34197_, _34196_);
  nor (_34198_, _34197_, _33734_);
  not (_34199_, _34198_);
  and (_34200_, _33734_, _34180_);
  nor (_34201_, _34200_, _34006_);
  and (_34202_, _34201_, _34199_);
  nor (_34203_, _34202_, _34190_);
  and (_34204_, _34196_, _34180_);
  nor (_34205_, _34204_, _33910_);
  nor (_34206_, _34196_, _34180_);
  nor (_34207_, _34206_, _34204_);
  and (_34208_, _34207_, _33914_);
  nor (_34209_, _34208_, _34205_);
  and (_34210_, _33922_, _34206_);
  and (_34211_, _33924_, _34180_);
  nor (_34212_, _34211_, _34210_);
  not (_34213_, _33934_);
  nor (_34214_, _34213_, _34180_);
  nor (_34215_, _33927_, _33935_);
  and (_34216_, _34215_, _33933_);
  nor (_34217_, _34216_, _34180_);
  nor (_34218_, _34217_, _34214_);
  and (_34219_, _34218_, _34212_);
  and (_34220_, _34219_, _34209_);
  and (_34221_, _34220_, _34203_);
  and (_34222_, _34221_, _33666_);
  nor (_34223_, _34222_, _34164_);
  nand (_34224_, _34223_, _33534_);
  not (_34225_, _33532_);
  and (_34226_, _34225_, _33474_);
  not (_34227_, _33604_);
  and (_34228_, _33571_, _33558_);
  and (_34229_, _34228_, _33644_);
  and (_34230_, _34229_, _33663_);
  nor (_34231_, _33630_, _33618_);
  not (_34232_, _33591_);
  nor (_34233_, _33604_, _34232_);
  and (_34234_, _34233_, _34231_);
  and (_34235_, _34234_, _34230_);
  not (_34236_, _34235_);
  and (_34237_, _34236_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_34238_, _34236_, _34017_);
  nor (_34239_, _34238_, _34237_);
  nor (_34240_, _34239_, _34227_);
  and (_34241_, _34239_, _34227_);
  nor (_34242_, _34241_, _34240_);
  nand (_34243_, _33559_, _33226_);
  or (_34244_, _33559_, _33226_);
  and (_34245_, _34244_, _34243_);
  not (_34246_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_34247_, _33659_, _34246_);
  not (_34248_, _34247_);
  and (_34249_, _33630_, _33618_);
  and (_34250_, _34249_, _33605_);
  not (_34251_, _33657_);
  and (_34252_, _33644_, _33571_);
  and (_34253_, _34252_, _33559_);
  and (_34254_, _34253_, _34251_);
  and (_34255_, _34254_, _34250_);
  not (_34256_, _34255_);
  and (_34257_, _34229_, _33657_);
  and (_34258_, _34250_, _34257_);
  and (_34259_, _34253_, _33657_);
  and (_34260_, _34250_, _34259_);
  nor (_34261_, _34260_, _34258_);
  and (_34262_, _34229_, _34251_);
  and (_34263_, _34262_, _34250_);
  not (_34264_, _34263_);
  and (_34265_, _34264_, _34261_);
  and (_34266_, _34265_, _34256_);
  and (_34267_, _34249_, _34233_);
  and (_34268_, _34267_, _34257_);
  and (_34269_, _34267_, _34259_);
  nor (_34270_, _34269_, _34268_);
  and (_34271_, _34267_, _34262_);
  not (_34272_, _34271_);
  and (_34273_, _34272_, _34270_);
  and (_34274_, _34273_, _34266_);
  or (_34275_, _34274_, _34248_);
  and (_34276_, _34254_, _34247_);
  and (_34277_, _34276_, _34267_);
  not (_34278_, _34277_);
  and (_34279_, _34278_, _34275_);
  nor (_34280_, _34279_, _34245_);
  and (_34281_, _34236_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_34282_, _34236_, _34052_);
  nor (_34283_, _34282_, _34281_);
  and (_34284_, _34283_, _34251_);
  nor (_34285_, _34283_, _34251_);
  nor (_34286_, _34285_, _34284_);
  and (_34287_, _34286_, _34280_);
  and (_34288_, _34287_, _34242_);
  and (_34289_, _34283_, _33226_);
  and (_34290_, _34289_, _34239_);
  nand (_34291_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_34292_, _34283_, _33464_);
  and (_34293_, _34292_, _34239_);
  nand (_34294_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_34295_, _34294_, _34291_);
  nor (_34296_, _34283_, _33464_);
  and (_34297_, _34296_, _34239_);
  nand (_34298_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_34299_, _34283_, _33226_);
  and (_34300_, _34299_, _34239_);
  nand (_34301_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_34302_, _34301_, _34298_);
  and (_34303_, _34302_, _34295_);
  not (_34304_, _34239_);
  and (_34305_, _34299_, _34304_);
  nand (_34306_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_34307_, _34296_, _34304_);
  nand (_34308_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_34309_, _34308_, _34306_);
  and (_34310_, _34289_, _34304_);
  nand (_34311_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_34312_, _34292_, _34304_);
  nand (_34313_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_34314_, _34313_, _34311_);
  and (_34315_, _34314_, _34309_);
  and (_34316_, _34315_, _34303_);
  nor (_34317_, _34316_, _34288_);
  not (_34318_, _34221_);
  and (_34319_, _34288_, _34318_);
  or (_34320_, _34319_, _34317_);
  nand (_34321_, _34320_, _34226_);
  and (_34322_, _33532_, _33499_);
  not (_34323_, _34322_);
  or (_34324_, _34323_, _33474_);
  not (_34325_, _33135_);
  and (_34326_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_34327_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_34328_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_34329_, _34328_, _34327_);
  and (_34330_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_34331_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34332_, _34331_, _34330_);
  and (_34333_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_34334_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_34335_, _33146_, _34334_);
  nor (_34336_, _34335_, _34333_);
  and (_34337_, _34336_, _34332_);
  and (_34338_, _34337_, _34329_);
  and (_34339_, _33141_, _33135_);
  not (_34340_, _34339_);
  nor (_34341_, _34340_, _34338_);
  nor (_34342_, _34341_, _34326_);
  or (_34343_, _34342_, _34324_);
  and (_34344_, _34343_, _33499_);
  and (_34345_, _34344_, _34321_);
  nand (_34346_, _34345_, _34224_);
  and (_34347_, _33376_, _33385_);
  and (_34348_, _34347_, _33464_);
  and (_34349_, _33423_, _33465_);
  or (_34350_, _34349_, _34348_);
  and (_34351_, _33437_, _33465_);
  nor (_34352_, _34351_, _34350_);
  and (_34353_, _34352_, _33362_);
  and (_34354_, _33418_, _33385_);
  and (_34355_, _34354_, _33464_);
  and (_34356_, _33397_, _33465_);
  or (_34357_, _34356_, _34355_);
  and (_34358_, _33388_, _33465_);
  and (_34359_, _33465_, _33408_);
  or (_34360_, _33416_, _33405_);
  or (_34361_, _34360_, _34359_);
  or (_34362_, _34361_, _34358_);
  nor (_34363_, _34362_, _34357_);
  and (_34364_, _34363_, _34353_);
  nor (_34365_, _34364_, _33477_);
  and (_34366_, _33360_, _33353_);
  not (_34367_, _33458_);
  nor (_34368_, _34367_, _34366_);
  nor (_34369_, _34368_, _34365_);
  or (_34370_, _34369_, _34346_);
  and (_34371_, _34226_, _33499_);
  not (_34372_, _34371_);
  and (_34373_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_34374_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_34375_, _34374_, _34373_);
  and (_34376_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_34377_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_34378_, _34377_, _34376_);
  and (_34379_, _34378_, _34375_);
  and (_34380_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_34381_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_34382_, _34381_, _34380_);
  and (_34383_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_34384_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_34385_, _34384_, _34383_);
  and (_34386_, _34385_, _34382_);
  and (_34387_, _34386_, _34379_);
  nor (_34388_, _34387_, _34288_);
  not (_34389_, _34052_);
  and (_34390_, _34288_, _34389_);
  nor (_34391_, _34390_, _34388_);
  or (_34392_, _34391_, _34372_);
  not (_34393_, _34283_);
  and (_34394_, _34322_, _33474_);
  and (_34395_, _34394_, _34393_);
  nor (_34396_, _34154_, _34055_);
  or (_34397_, _34396_, _34155_);
  nand (_34398_, _34397_, _33578_);
  nand (_34399_, _34398_, _33652_);
  and (_34400_, _34399_, _33667_);
  or (_34401_, _34400_, _34053_);
  nand (_34402_, _34401_, _33534_);
  and (_34403_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_34404_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  not (_34405_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_34406_, _33146_, _34405_);
  nor (_34407_, _34406_, _34404_);
  and (_34408_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_34409_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_34410_, _34409_, _34408_);
  and (_34411_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_34412_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_34413_, _34412_, _34411_);
  and (_34414_, _34413_, _34410_);
  and (_34415_, _34414_, _34407_);
  nor (_34416_, _34415_, _34340_);
  nor (_34417_, _34416_, _34403_);
  or (_34418_, _34417_, _34324_);
  nand (_34419_, _34418_, _34402_);
  nor (_34420_, _34419_, _34395_);
  and (_34421_, _34420_, _34392_);
  or (_34422_, _34421_, _34370_);
  not (_34423_, _34369_);
  and (_34424_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_34425_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_34426_, _34425_, _34424_);
  and (_34427_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_34428_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_34429_, _34428_, _34427_);
  and (_34430_, _34429_, _34426_);
  and (_34431_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_34432_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_34433_, _34432_, _34431_);
  and (_34434_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_34435_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_34436_, _34435_, _34434_);
  and (_34437_, _34436_, _34433_);
  and (_34438_, _34437_, _34430_);
  nor (_34439_, _34438_, _34288_);
  and (_34440_, _34288_, _34149_);
  nor (_34441_, _34440_, _34439_);
  or (_34442_, _34441_, _34372_);
  and (_34443_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_34444_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  not (_34445_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_34446_, _33146_, _34445_);
  nor (_34447_, _34446_, _34444_);
  and (_34448_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_34449_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_34450_, _34449_, _34448_);
  and (_34451_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_34452_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_34453_, _34452_, _34451_);
  and (_34454_, _34453_, _34450_);
  and (_34455_, _34454_, _34447_);
  nor (_34456_, _34455_, _34340_);
  nor (_34457_, _34456_, _34443_);
  nor (_34458_, _34457_, _34324_);
  not (_34459_, _33534_);
  nor (_34460_, _34151_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_34461_, _34460_, _34152_);
  nor (_34462_, _34461_, _33551_);
  nor (_34463_, _34462_, _33552_);
  nor (_34464_, _34463_, _33666_);
  not (_34465_, _34464_);
  and (_34466_, _34465_, _34150_);
  or (_34467_, _34466_, _34459_);
  nand (_34468_, _34394_, _33226_);
  nand (_34469_, _34468_, _34467_);
  nor (_34470_, _34469_, _34458_);
  and (_34471_, _34470_, _34442_);
  or (_34472_, _34471_, _34423_);
  nand (_34473_, _34472_, _34422_);
  and (_34474_, _33618_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_34475_, _34474_, _34251_);
  nor (_34476_, _33558_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_34477_, _34476_, _34475_);
  nor (_34478_, _34477_, _34473_);
  and (_34479_, _34477_, _34473_);
  nor (_34480_, _34479_, _34478_);
  and (_34481_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_34482_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  not (_34483_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_34484_, _33146_, _34483_);
  nor (_34485_, _34484_, _34482_);
  and (_34486_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_34487_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_34488_, _34487_, _34486_);
  and (_34489_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_34490_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_34491_, _34490_, _34489_);
  and (_34492_, _34491_, _34488_);
  and (_34493_, _34492_, _34485_);
  nor (_34494_, _34493_, _34340_);
  nor (_34495_, _34494_, _34481_);
  nor (_34496_, _34495_, _34324_);
  and (_34497_, _34394_, _34304_);
  nor (_34498_, _34497_, _34496_);
  and (_34499_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_34500_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_34501_, _34500_, _34499_);
  and (_34502_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_34503_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_34504_, _34503_, _34502_);
  and (_34505_, _34504_, _34501_);
  and (_34506_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_34507_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_34508_, _34507_, _34506_);
  and (_34509_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_34510_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_34511_, _34510_, _34509_);
  and (_34512_, _34511_, _34508_);
  and (_34513_, _34512_, _34505_);
  nor (_34514_, _34513_, _34288_);
  not (_34515_, _34017_);
  and (_34516_, _34288_, _34515_);
  nor (_34517_, _34516_, _34514_);
  or (_34518_, _34517_, _34372_);
  and (_34519_, _33532_, _33500_);
  nor (_34520_, _34155_, _34019_);
  or (_34521_, _34520_, _34156_);
  and (_34522_, _34521_, _33578_);
  or (_34523_, _34522_, _33597_);
  and (_34524_, _34523_, _33667_);
  or (_34525_, _34524_, _34018_);
  and (_34526_, _34525_, _33534_);
  nor (_34527_, _34526_, _34519_);
  and (_34528_, _34527_, _34518_);
  and (_34529_, _34528_, _34498_);
  or (_34530_, _34529_, _34370_);
  and (_34531_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_34532_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_34533_, _34532_, _34531_);
  and (_34534_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_34535_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_34536_, _34535_, _34534_);
  and (_34537_, _34536_, _34533_);
  and (_34538_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_34539_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_34540_, _34539_, _34538_);
  and (_34541_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_34542_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_34543_, _34542_, _34541_);
  and (_34544_, _34543_, _34540_);
  and (_34545_, _34544_, _34537_);
  nor (_34546_, _34545_, _34288_);
  and (_34547_, _34288_, _34122_);
  nor (_34548_, _34547_, _34546_);
  nor (_34549_, _34548_, _34372_);
  not (_34550_, _34549_);
  and (_34551_, _34226_, _33500_);
  nor (_34552_, _34152_, _34124_);
  nor (_34553_, _34552_, _34153_);
  nor (_34554_, _34553_, _33551_);
  nor (_34555_, _34554_, _33563_);
  nor (_34556_, _34555_, _33666_);
  nor (_34557_, _34556_, _34123_);
  not (_34558_, _34557_);
  and (_34559_, _34558_, _33534_);
  nor (_34560_, _34559_, _34551_);
  and (_34561_, _34394_, _33250_);
  and (_34562_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_34563_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_34564_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_34565_, _34564_, _34563_);
  and (_34566_, _33236_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_34567_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_34568_, _34567_, _34566_);
  and (_34569_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_34570_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_34571_, _34570_, _34569_);
  and (_34572_, _34571_, _34568_);
  and (_34573_, _34572_, _34565_);
  nor (_34574_, _34573_, _34340_);
  nor (_34575_, _34574_, _34562_);
  nor (_34576_, _34575_, _34324_);
  nor (_34577_, _34576_, _34561_);
  and (_34578_, _34577_, _34560_);
  and (_34579_, _34578_, _34550_);
  or (_34580_, _34579_, _34423_);
  and (_34581_, _34580_, _34530_);
  and (_34582_, _34474_, _34227_);
  nor (_34583_, _33571_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_34584_, _34583_, _34582_);
  and (_34585_, _34584_, _34581_);
  nor (_34586_, _34584_, _34581_);
  or (_34587_, _34586_, _34585_);
  and (_34588_, _34587_, _34480_);
  and (_34589_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_34590_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not (_34591_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34592_, _33146_, _34591_);
  nor (_34593_, _34592_, _34590_);
  and (_34594_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_34595_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_34596_, _34595_, _34594_);
  and (_34597_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34598_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_34599_, _34598_, _34597_);
  and (_34600_, _34599_, _34596_);
  and (_34601_, _34600_, _34593_);
  nor (_34602_, _34601_, _34340_);
  nor (_34603_, _34602_, _34589_);
  nor (_34604_, _34603_, _34324_);
  nor (_34605_, _34225_, _33474_);
  not (_34606_, _34605_);
  nor (_34607_, _34226_, _33499_);
  and (_34608_, _34607_, _34606_);
  or (_34609_, _34608_, _34604_);
  nor (_34610_, _34156_, _33980_);
  nor (_34611_, _34610_, _34157_);
  nor (_34612_, _34611_, _33551_);
  nor (_34613_, _34612_, _33581_);
  nor (_34614_, _34613_, _33666_);
  nor (_34615_, _34614_, _33979_);
  nor (_34616_, _34615_, _34459_);
  and (_34617_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_34618_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_34619_, _34618_, _34617_);
  and (_34620_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_34621_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_34622_, _34621_, _34620_);
  and (_34623_, _34622_, _34619_);
  and (_34624_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_34625_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_34626_, _34625_, _34624_);
  and (_34627_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_34628_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_34629_, _34628_, _34627_);
  and (_34630_, _34629_, _34626_);
  and (_34631_, _34630_, _34623_);
  nor (_34632_, _34631_, _34288_);
  and (_34633_, _34288_, _33978_);
  nor (_34634_, _34633_, _34632_);
  nor (_34635_, _34634_, _34372_);
  or (_34636_, _34635_, _34616_);
  nor (_34637_, _34636_, _34609_);
  and (_34638_, _34637_, _34370_);
  nor (_34639_, _34474_, _34232_);
  not (_34640_, _34639_);
  nor (_34641_, _34640_, _34638_);
  not (_34642_, _34641_);
  not (_34643_, _34370_);
  nor (_34644_, _34157_, _33944_);
  nor (_34645_, _34644_, _34158_);
  nor (_34646_, _34645_, _33551_);
  nor (_34647_, _34646_, _33622_);
  nor (_34648_, _34647_, _33666_);
  nor (_34649_, _34648_, _33943_);
  nor (_34650_, _34649_, _34459_);
  not (_34651_, _34650_);
  and (_34652_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_34653_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_34654_, _34653_, _34652_);
  and (_34655_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_34656_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_34657_, _34656_, _34655_);
  and (_34658_, _34657_, _34654_);
  and (_34659_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_34660_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_34661_, _34660_, _34659_);
  and (_34662_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_34663_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_34664_, _34663_, _34662_);
  and (_34665_, _34664_, _34661_);
  and (_34666_, _34665_, _34658_);
  nor (_34667_, _34666_, _34288_);
  and (_34668_, _34288_, _33942_);
  nor (_34669_, _34668_, _34667_);
  nor (_34670_, _34669_, _34372_);
  and (_34671_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_34672_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not (_34673_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_34674_, _33146_, _34673_);
  nor (_34675_, _34674_, _34672_);
  and (_34676_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_34677_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_34678_, _34677_, _34676_);
  and (_34679_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34680_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34681_, _34680_, _34679_);
  and (_34682_, _34681_, _34678_);
  and (_34683_, _34682_, _34675_);
  nor (_34684_, _34683_, _34340_);
  nor (_34685_, _34684_, _34671_);
  not (_34686_, _34685_);
  and (_34687_, _34686_, _34605_);
  nor (_34688_, _34607_, _34687_);
  not (_34689_, _34688_);
  nor (_34690_, _34689_, _34670_);
  and (_34691_, _34690_, _34651_);
  nor (_34692_, _34691_, _34643_);
  nor (_34693_, _34474_, _33630_);
  not (_34694_, _34693_);
  and (_34695_, _34694_, _34692_);
  nor (_34696_, _34694_, _34692_);
  nor (_34697_, _34696_, _34695_);
  and (_34698_, _34697_, _34642_);
  not (_34699_, _34529_);
  and (_34700_, _34699_, _34370_);
  nor (_34701_, _34474_, _33604_);
  not (_34702_, _34701_);
  and (_34703_, _34702_, _34700_);
  and (_34704_, _34640_, _34638_);
  nor (_34705_, _34704_, _34703_);
  not (_34706_, _33618_);
  and (_34707_, _34346_, _34706_);
  nor (_34708_, _34346_, _34706_);
  nor (_34709_, _34708_, _34707_);
  not (_34710_, _34709_);
  and (_34711_, _34710_, _34705_);
  and (_34712_, _34711_, _34698_);
  and (_34713_, _34712_, _34588_);
  and (_34714_, _34474_, _33631_);
  nor (_34715_, _34474_, _33657_);
  nor (_34716_, _34715_, _34714_);
  and (_34717_, _34691_, _34643_);
  and (_34718_, _34421_, _34370_);
  nor (_34719_, _34718_, _34717_);
  and (_34720_, _34719_, _34716_);
  nor (_34721_, _34719_, _34716_);
  or (_34722_, _34721_, _34720_);
  nor (_34723_, _34637_, _34370_);
  and (_34724_, _34300_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_34725_, _34297_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_34726_, _34725_, _34724_);
  and (_34727_, _34290_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_34728_, _34293_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_34729_, _34728_, _34727_);
  and (_34730_, _34729_, _34726_);
  and (_34731_, _34305_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_34732_, _34312_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_34733_, _34732_, _34731_);
  and (_34734_, _34310_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_34735_, _34307_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_34736_, _34735_, _34734_);
  and (_34737_, _34736_, _34733_);
  and (_34738_, _34737_, _34730_);
  nor (_34739_, _34738_, _34288_);
  and (_34740_, _34288_, _34089_);
  nor (_34741_, _34740_, _34739_);
  nor (_34742_, _34741_, _34372_);
  and (_34743_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_34744_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_34745_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_34746_, _34745_, _34744_);
  not (_34747_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_34748_, _33146_, _34747_);
  and (_34749_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_34750_, _34749_, _34748_);
  and (_34751_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_34752_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_34753_, _34752_, _34751_);
  and (_34754_, _34753_, _34750_);
  and (_34755_, _34754_, _34746_);
  nor (_34756_, _34755_, _34340_);
  nor (_34757_, _34756_, _34743_);
  nor (_34758_, _34757_, _34324_);
  nor (_34759_, _34758_, _34742_);
  and (_34760_, _34394_, _33177_);
  nor (_34761_, _34153_, _34091_);
  nor (_34762_, _34761_, _34154_);
  nor (_34763_, _34762_, _33551_);
  nor (_34764_, _34763_, _33636_);
  nor (_34765_, _34764_, _33666_);
  nor (_34766_, _34765_, _34090_);
  not (_34767_, _34766_);
  and (_34768_, _34767_, _33534_);
  nor (_34769_, _34768_, _34760_);
  and (_34770_, _34769_, _34759_);
  nor (_34771_, _34770_, _34423_);
  nor (_34772_, _34771_, _34723_);
  and (_34773_, _34474_, _34232_);
  nor (_34774_, _33644_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_34775_, _34774_, _34773_);
  not (_34776_, _34775_);
  and (_34777_, _34776_, _34772_);
  nor (_34778_, _34776_, _34772_);
  nor (_34779_, _34778_, _34777_);
  not (_34780_, _34779_);
  nor (_34781_, _34780_, _34722_);
  nor (_34782_, _34702_, _34700_);
  nor (_34783_, _33618_, _33550_);
  nor (_34784_, _34783_, _33660_);
  not (_34785_, _34784_);
  nor (_34786_, _34785_, _34782_);
  and (_34787_, _34786_, _34781_);
  and (_34788_, _34787_, _34713_);
  not (_34789_, _34700_);
  not (_34790_, _34772_);
  and (_34791_, _34472_, _34422_);
  and (_34792_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_34793_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_34794_, _34793_, _34792_);
  and (_34795_, _34794_, _34581_);
  not (_34796_, _34581_);
  and (_34797_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_34798_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_34799_, _34798_, _34797_);
  and (_34800_, _34799_, _34796_);
  or (_34801_, _34800_, _34795_);
  or (_34802_, _34801_, _34790_);
  not (_34803_, _34719_);
  and (_34804_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_34805_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_34806_, _34805_, _34804_);
  and (_34807_, _34806_, _34581_);
  and (_34808_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_34809_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_34810_, _34809_, _34808_);
  and (_34811_, _34810_, _34796_);
  or (_34812_, _34811_, _34807_);
  or (_34813_, _34812_, _34772_);
  and (_34814_, _34813_, _34803_);
  and (_34815_, _34814_, _34802_);
  or (_34816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_34817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_34818_, _34817_, _34816_);
  and (_34819_, _34818_, _34581_);
  or (_34820_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_34821_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_34822_, _34821_, _34820_);
  and (_34823_, _34822_, _34796_);
  or (_34824_, _34823_, _34819_);
  or (_34825_, _34824_, _34790_);
  or (_34826_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_34827_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_34828_, _34827_, _34826_);
  and (_34829_, _34828_, _34581_);
  or (_34830_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_34831_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_34832_, _34831_, _34830_);
  and (_34833_, _34832_, _34796_);
  or (_34834_, _34833_, _34829_);
  or (_34835_, _34834_, _34772_);
  and (_34836_, _34835_, _34719_);
  and (_34837_, _34836_, _34825_);
  or (_34838_, _34837_, _34815_);
  or (_34839_, _34838_, _34789_);
  not (_34840_, _34638_);
  and (_34841_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_34842_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_34843_, _34842_, _34841_);
  and (_34844_, _34843_, _34581_);
  and (_34845_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_34846_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_34847_, _34846_, _34845_);
  and (_34848_, _34847_, _34796_);
  or (_34849_, _34848_, _34844_);
  or (_34850_, _34849_, _34790_);
  and (_34851_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_34852_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_34853_, _34852_, _34851_);
  and (_34854_, _34853_, _34581_);
  and (_34855_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_34856_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_34857_, _34856_, _34855_);
  and (_34858_, _34857_, _34796_);
  or (_34859_, _34858_, _34854_);
  or (_34860_, _34859_, _34772_);
  and (_34861_, _34860_, _34803_);
  and (_34862_, _34861_, _34850_);
  or (_34863_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_34864_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_34865_, _34864_, _34796_);
  and (_34866_, _34865_, _34863_);
  or (_34867_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_34868_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_34869_, _34868_, _34581_);
  and (_34870_, _34869_, _34867_);
  or (_34871_, _34870_, _34866_);
  or (_34872_, _34871_, _34790_);
  or (_34873_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_34874_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_34875_, _34874_, _34796_);
  and (_34876_, _34875_, _34873_);
  or (_34877_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_34878_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_34879_, _34878_, _34581_);
  and (_34880_, _34879_, _34877_);
  or (_34881_, _34880_, _34876_);
  or (_34882_, _34881_, _34772_);
  and (_34883_, _34882_, _34719_);
  and (_34884_, _34883_, _34872_);
  or (_34885_, _34884_, _34862_);
  or (_34886_, _34885_, _34700_);
  and (_34887_, _34886_, _34840_);
  and (_34888_, _34887_, _34839_);
  and (_34889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_34890_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_34891_, _34890_, _34889_);
  and (_34892_, _34891_, _34581_);
  and (_34893_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_34894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_34895_, _34894_, _34893_);
  and (_34896_, _34895_, _34796_);
  or (_34897_, _34896_, _34892_);
  and (_34898_, _34897_, _34772_);
  and (_34899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_34900_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_34901_, _34900_, _34899_);
  and (_34902_, _34901_, _34581_);
  and (_34903_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_34904_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_34905_, _34904_, _34903_);
  and (_34906_, _34905_, _34796_);
  or (_34907_, _34906_, _34902_);
  and (_34908_, _34907_, _34790_);
  or (_34909_, _34908_, _34719_);
  or (_34910_, _34909_, _34898_);
  or (_34911_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_34912_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_34913_, _34912_, _34796_);
  and (_34914_, _34913_, _34911_);
  or (_34915_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_34916_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_34917_, _34916_, _34581_);
  and (_34918_, _34917_, _34915_);
  or (_34919_, _34918_, _34914_);
  and (_34920_, _34919_, _34772_);
  or (_34921_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_34922_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_34923_, _34922_, _34796_);
  and (_34924_, _34923_, _34921_);
  or (_34925_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_34926_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_34927_, _34926_, _34581_);
  and (_34928_, _34927_, _34925_);
  or (_34929_, _34928_, _34924_);
  and (_34930_, _34929_, _34790_);
  or (_34931_, _34930_, _34803_);
  or (_34932_, _34931_, _34920_);
  and (_34933_, _34932_, _34910_);
  or (_34934_, _34933_, _34700_);
  and (_34935_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_34936_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_34937_, _34936_, _34935_);
  and (_34938_, _34937_, _34581_);
  and (_34939_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_34940_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_34941_, _34940_, _34939_);
  and (_34942_, _34941_, _34796_);
  or (_34943_, _34942_, _34938_);
  and (_34944_, _34943_, _34772_);
  and (_34945_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_34946_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_34947_, _34946_, _34945_);
  and (_34948_, _34947_, _34581_);
  and (_34949_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_34950_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_34951_, _34950_, _34949_);
  and (_34952_, _34951_, _34796_);
  or (_34953_, _34952_, _34948_);
  and (_34954_, _34953_, _34790_);
  or (_34955_, _34954_, _34719_);
  or (_34956_, _34955_, _34944_);
  or (_34957_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_34958_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_34959_, _34958_, _34957_);
  and (_34960_, _34959_, _34581_);
  or (_34961_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_34962_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_34963_, _34962_, _34961_);
  and (_34964_, _34963_, _34796_);
  or (_34965_, _34964_, _34960_);
  and (_34966_, _34965_, _34772_);
  or (_34967_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_34968_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_34969_, _34968_, _34967_);
  and (_34970_, _34969_, _34581_);
  or (_34971_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_34972_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_34973_, _34972_, _34971_);
  and (_34974_, _34973_, _34796_);
  or (_34975_, _34974_, _34970_);
  and (_34976_, _34975_, _34790_);
  or (_34977_, _34976_, _34803_);
  or (_34978_, _34977_, _34966_);
  and (_34979_, _34978_, _34956_);
  or (_34980_, _34979_, _34789_);
  and (_34981_, _34980_, _34638_);
  and (_34982_, _34981_, _34934_);
  or (_34983_, _34982_, _34888_);
  or (_34984_, _34983_, _34692_);
  not (_34985_, _34692_);
  and (_34986_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and (_34987_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_34988_, _34987_, _34986_);
  and (_34989_, _34988_, _34581_);
  and (_34990_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  and (_34991_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or (_34992_, _34991_, _34990_);
  and (_34993_, _34992_, _34796_);
  or (_34994_, _34993_, _34989_);
  and (_34995_, _34994_, _34772_);
  and (_34996_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  and (_34997_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_34998_, _34997_, _34996_);
  and (_34999_, _34998_, _34581_);
  and (_35000_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  and (_35001_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or (_35002_, _35001_, _35000_);
  and (_35003_, _35002_, _34796_);
  or (_35004_, _35003_, _34999_);
  and (_35005_, _35004_, _34790_);
  or (_35006_, _35005_, _34719_);
  or (_35007_, _35006_, _34995_);
  or (_35008_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or (_35009_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and (_35010_, _35009_, _35008_);
  and (_35011_, _35010_, _34581_);
  or (_35012_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_35013_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  and (_35014_, _35013_, _35012_);
  and (_35015_, _35014_, _34796_);
  or (_35016_, _35015_, _35011_);
  and (_35017_, _35016_, _34772_);
  or (_35018_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or (_35019_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and (_35020_, _35019_, _35018_);
  and (_35021_, _35020_, _34581_);
  or (_35022_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or (_35023_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  and (_35024_, _35023_, _35022_);
  and (_35025_, _35024_, _34796_);
  or (_35026_, _35025_, _35021_);
  and (_35027_, _35026_, _34790_);
  or (_35028_, _35027_, _34803_);
  or (_35029_, _35028_, _35017_);
  and (_35030_, _35029_, _35007_);
  or (_35031_, _35030_, _34700_);
  and (_35032_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_35033_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_35034_, _35033_, _35032_);
  and (_35035_, _35034_, _34581_);
  and (_35036_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_35037_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_35038_, _35037_, _35036_);
  and (_35039_, _35038_, _34796_);
  or (_35040_, _35039_, _35035_);
  and (_35041_, _35040_, _34772_);
  and (_35042_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_35043_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_35044_, _35043_, _35042_);
  and (_35045_, _35044_, _34581_);
  and (_35046_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_35047_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_35048_, _35047_, _35046_);
  and (_35049_, _35048_, _34796_);
  or (_35050_, _35049_, _35045_);
  and (_35051_, _35050_, _34790_);
  or (_35052_, _35051_, _34719_);
  or (_35053_, _35052_, _35041_);
  or (_35054_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_35055_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_35056_, _35055_, _35054_);
  and (_35057_, _35056_, _34581_);
  or (_35058_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_35059_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_35060_, _35059_, _35058_);
  and (_35061_, _35060_, _34796_);
  or (_35062_, _35061_, _35057_);
  and (_35063_, _35062_, _34772_);
  or (_35064_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_35065_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_35066_, _35065_, _35064_);
  and (_35067_, _35066_, _34581_);
  or (_35068_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_35069_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_35070_, _35069_, _35068_);
  and (_35071_, _35070_, _34796_);
  or (_35072_, _35071_, _35067_);
  and (_35073_, _35072_, _34790_);
  or (_35074_, _35073_, _34803_);
  or (_35075_, _35074_, _35063_);
  and (_35076_, _35075_, _35053_);
  or (_35077_, _35076_, _34789_);
  and (_35078_, _35077_, _34638_);
  and (_35079_, _35078_, _35031_);
  and (_35080_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_35081_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_35082_, _35081_, _35080_);
  and (_35083_, _35082_, _34796_);
  and (_35084_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_35085_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_35086_, _35085_, _35084_);
  and (_35087_, _35086_, _34581_);
  or (_35088_, _35087_, _35083_);
  or (_35089_, _35088_, _34790_);
  and (_35090_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_35091_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_35092_, _35091_, _35090_);
  and (_35093_, _35092_, _34796_);
  and (_35094_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_35095_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_35096_, _35095_, _35094_);
  and (_35097_, _35096_, _34581_);
  or (_35098_, _35097_, _35093_);
  or (_35099_, _35098_, _34772_);
  and (_35100_, _35099_, _34803_);
  and (_35101_, _35100_, _35089_);
  or (_35102_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_35103_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_35104_, _35103_, _34581_);
  and (_35105_, _35104_, _35102_);
  or (_35106_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_35107_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_35108_, _35107_, _34796_);
  and (_35109_, _35108_, _35106_);
  or (_35110_, _35109_, _35105_);
  or (_35111_, _35110_, _34790_);
  or (_35112_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_35113_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_35114_, _35113_, _34581_);
  and (_35115_, _35114_, _35112_);
  or (_35116_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_35117_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_35118_, _35117_, _34796_);
  and (_35119_, _35118_, _35116_);
  or (_35120_, _35119_, _35115_);
  or (_35121_, _35120_, _34772_);
  and (_35122_, _35121_, _34719_);
  and (_35123_, _35122_, _35111_);
  or (_35124_, _35123_, _35101_);
  and (_35125_, _35124_, _34789_);
  and (_35126_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_35127_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_35128_, _35127_, _34581_);
  or (_35129_, _35128_, _35126_);
  and (_35130_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_35131_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_35132_, _35131_, _34796_);
  or (_35133_, _35132_, _35130_);
  and (_35134_, _35133_, _35129_);
  or (_35135_, _35134_, _34790_);
  and (_35136_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_35137_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_35138_, _35137_, _34581_);
  or (_35139_, _35138_, _35136_);
  and (_35140_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_35141_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_35142_, _35141_, _34796_);
  or (_35143_, _35142_, _35140_);
  and (_35144_, _35143_, _35139_);
  or (_35145_, _35144_, _34772_);
  and (_35146_, _35145_, _34803_);
  and (_35147_, _35146_, _35135_);
  or (_35148_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_35149_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_35150_, _35149_, _35148_);
  or (_35151_, _35150_, _34796_);
  or (_35152_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_35153_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_35154_, _35153_, _35152_);
  or (_35155_, _35154_, _34581_);
  and (_35156_, _35155_, _35151_);
  or (_35157_, _35156_, _34790_);
  or (_35158_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_35159_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_35160_, _35159_, _35158_);
  or (_35161_, _35160_, _34796_);
  or (_35162_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_35163_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_35164_, _35163_, _35162_);
  or (_35165_, _35164_, _34581_);
  and (_35166_, _35165_, _35161_);
  or (_35167_, _35166_, _34772_);
  and (_35168_, _35167_, _34719_);
  and (_35169_, _35168_, _35157_);
  or (_35170_, _35169_, _35147_);
  and (_35171_, _35170_, _34700_);
  or (_35172_, _35171_, _35125_);
  and (_35173_, _35172_, _34840_);
  or (_35174_, _35173_, _35079_);
  or (_35175_, _35174_, _34985_);
  and (_35176_, _35175_, _34984_);
  or (_35177_, _35176_, _34346_);
  not (_35178_, _34346_);
  and (_35179_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_35180_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_35181_, _35180_, _35179_);
  and (_35182_, _35181_, _34796_);
  and (_35183_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_35184_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_35185_, _35184_, _35183_);
  and (_35186_, _35185_, _34581_);
  or (_35187_, _35186_, _35182_);
  or (_35188_, _35187_, _34790_);
  and (_35189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_35190_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_35191_, _35190_, _35189_);
  and (_35192_, _35191_, _34796_);
  and (_35193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_35194_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_35195_, _35194_, _35193_);
  and (_35196_, _35195_, _34581_);
  or (_35197_, _35196_, _35192_);
  or (_35198_, _35197_, _34772_);
  and (_35199_, _35198_, _34803_);
  and (_35200_, _35199_, _35188_);
  or (_35201_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_35202_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_35203_, _35202_, _34581_);
  and (_35204_, _35203_, _35201_);
  or (_35205_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_35206_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_35207_, _35206_, _34796_);
  and (_35208_, _35207_, _35205_);
  or (_35209_, _35208_, _35204_);
  or (_35210_, _35209_, _34790_);
  or (_35211_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_35212_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_35213_, _35212_, _34581_);
  and (_35214_, _35213_, _35211_);
  or (_35215_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_35216_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_35217_, _35216_, _34796_);
  and (_35218_, _35217_, _35215_);
  or (_35219_, _35218_, _35214_);
  or (_35220_, _35219_, _34772_);
  and (_35221_, _35220_, _34719_);
  and (_35222_, _35221_, _35210_);
  or (_35223_, _35222_, _35200_);
  and (_35224_, _35223_, _34789_);
  and (_35225_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_35226_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_35227_, _35226_, _34581_);
  or (_35228_, _35227_, _35225_);
  and (_35229_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_35230_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_35231_, _35230_, _34796_);
  or (_35232_, _35231_, _35229_);
  and (_35233_, _35232_, _35228_);
  or (_35234_, _35233_, _34790_);
  and (_35235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_35236_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_35237_, _35236_, _34581_);
  or (_35238_, _35237_, _35235_);
  and (_35239_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_35240_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_35241_, _35240_, _34796_);
  or (_35242_, _35241_, _35239_);
  and (_35243_, _35242_, _35238_);
  or (_35244_, _35243_, _34772_);
  and (_35245_, _35244_, _34803_);
  and (_35246_, _35245_, _35234_);
  or (_35247_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_35248_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_35249_, _35248_, _35247_);
  or (_35250_, _35249_, _34796_);
  or (_35251_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_35252_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_35253_, _35252_, _35251_);
  or (_35254_, _35253_, _34581_);
  and (_35255_, _35254_, _35250_);
  or (_35256_, _35255_, _34790_);
  or (_35257_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_35258_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_35259_, _35258_, _35257_);
  or (_35260_, _35259_, _34796_);
  or (_35261_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_35262_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_35263_, _35262_, _35261_);
  or (_35264_, _35263_, _34581_);
  and (_35265_, _35264_, _35260_);
  or (_35266_, _35265_, _34772_);
  and (_35267_, _35266_, _34719_);
  and (_35268_, _35267_, _35256_);
  or (_35269_, _35268_, _35246_);
  and (_35270_, _35269_, _34700_);
  or (_35271_, _35270_, _35224_);
  and (_35272_, _35271_, _34840_);
  and (_35273_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  and (_35274_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_35275_, _35274_, _35273_);
  and (_35276_, _35275_, _34581_);
  and (_35277_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  and (_35278_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_35279_, _35278_, _35277_);
  and (_35280_, _35279_, _34796_);
  or (_35281_, _35280_, _35276_);
  and (_35282_, _35281_, _34772_);
  and (_35283_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and (_35284_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_35285_, _35284_, _35283_);
  and (_35286_, _35285_, _34581_);
  and (_35287_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and (_35288_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or (_35289_, _35288_, _35287_);
  and (_35290_, _35289_, _34796_);
  or (_35291_, _35290_, _35286_);
  and (_35292_, _35291_, _34790_);
  or (_35293_, _35292_, _35282_);
  and (_35294_, _35293_, _34803_);
  or (_35295_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_35296_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and (_35297_, _35296_, _35295_);
  and (_35298_, _35297_, _34581_);
  or (_35299_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or (_35300_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and (_35301_, _35300_, _35299_);
  and (_35302_, _35301_, _34796_);
  or (_35303_, _35302_, _35298_);
  and (_35304_, _35303_, _34772_);
  or (_35305_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_35306_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and (_35307_, _35306_, _35305_);
  and (_35308_, _35307_, _34581_);
  or (_35309_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_35310_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and (_35311_, _35310_, _35309_);
  and (_35312_, _35311_, _34796_);
  or (_35313_, _35312_, _35308_);
  and (_35314_, _35313_, _34790_);
  or (_35315_, _35314_, _35304_);
  and (_35316_, _35315_, _34719_);
  or (_35317_, _35316_, _35294_);
  and (_35318_, _35317_, _34789_);
  and (_35319_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_35320_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_35321_, _35320_, _35319_);
  and (_35322_, _35321_, _34581_);
  and (_35323_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_35324_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_35325_, _35324_, _35323_);
  and (_35326_, _35325_, _34796_);
  or (_35327_, _35326_, _35322_);
  and (_35328_, _35327_, _34772_);
  and (_35329_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_35330_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_35331_, _35330_, _35329_);
  and (_35332_, _35331_, _34581_);
  and (_35333_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_35334_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_35335_, _35334_, _35333_);
  and (_35336_, _35335_, _34796_);
  or (_35337_, _35336_, _35332_);
  and (_35338_, _35337_, _34790_);
  or (_35339_, _35338_, _35328_);
  and (_35340_, _35339_, _34803_);
  or (_35341_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_35342_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_35343_, _35342_, _35341_);
  and (_35344_, _35343_, _34581_);
  or (_35345_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_35346_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_35347_, _35346_, _35345_);
  and (_35348_, _35347_, _34796_);
  or (_35349_, _35348_, _35344_);
  and (_35350_, _35349_, _34772_);
  or (_35351_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_35352_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_35353_, _35352_, _35351_);
  and (_35354_, _35353_, _34581_);
  or (_35355_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_35356_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_35357_, _35356_, _35355_);
  and (_35358_, _35357_, _34796_);
  or (_35359_, _35358_, _35354_);
  and (_35360_, _35359_, _34790_);
  or (_35361_, _35360_, _35350_);
  and (_35362_, _35361_, _34719_);
  or (_35363_, _35362_, _35340_);
  and (_35364_, _35363_, _34700_);
  or (_35365_, _35364_, _35318_);
  and (_35366_, _35365_, _34638_);
  or (_35367_, _35366_, _35272_);
  or (_35368_, _35367_, _34692_);
  and (_35369_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_35370_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_35371_, _35370_, _35369_);
  and (_35372_, _35371_, _34581_);
  and (_35373_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_35374_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_35375_, _35374_, _35373_);
  and (_35376_, _35375_, _34796_);
  or (_35377_, _35376_, _35372_);
  or (_35378_, _35377_, _34790_);
  and (_35379_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_35380_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_35381_, _35380_, _35379_);
  and (_35382_, _35381_, _34581_);
  and (_35383_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_35384_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_35385_, _35384_, _35383_);
  and (_35386_, _35385_, _34796_);
  or (_35387_, _35386_, _35382_);
  or (_35388_, _35387_, _34772_);
  and (_35389_, _35388_, _34803_);
  and (_35390_, _35389_, _35378_);
  or (_35391_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_35392_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_35393_, _35392_, _34796_);
  and (_35394_, _35393_, _35391_);
  or (_35395_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_35396_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_35397_, _35396_, _34581_);
  and (_35398_, _35397_, _35395_);
  or (_35399_, _35398_, _35394_);
  or (_35400_, _35399_, _34790_);
  or (_35401_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_35402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_35403_, _35402_, _34796_);
  and (_35404_, _35403_, _35401_);
  or (_35405_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_35406_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_35407_, _35406_, _34581_);
  and (_35408_, _35407_, _35405_);
  or (_35409_, _35408_, _35404_);
  or (_35410_, _35409_, _34772_);
  and (_35411_, _35410_, _34719_);
  and (_35412_, _35411_, _35400_);
  or (_35413_, _35412_, _35390_);
  and (_35414_, _35413_, _34789_);
  and (_35415_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_35416_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_35417_, _35416_, _35415_);
  and (_35418_, _35417_, _34581_);
  and (_35419_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_35420_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_35421_, _35420_, _35419_);
  and (_35422_, _35421_, _34796_);
  or (_35423_, _35422_, _35418_);
  or (_35424_, _35423_, _34790_);
  and (_35425_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_35426_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_35427_, _35426_, _35425_);
  and (_35428_, _35427_, _34581_);
  and (_35429_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_35430_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_35431_, _35430_, _35429_);
  and (_35432_, _35431_, _34796_);
  or (_35433_, _35432_, _35428_);
  or (_35434_, _35433_, _34772_);
  and (_35435_, _35434_, _34803_);
  and (_35436_, _35435_, _35424_);
  or (_35437_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_35438_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_35439_, _35438_, _35437_);
  and (_35440_, _35439_, _34581_);
  or (_35441_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_35442_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_35443_, _35442_, _35441_);
  and (_35444_, _35443_, _34796_);
  or (_35445_, _35444_, _35440_);
  or (_35446_, _35445_, _34790_);
  or (_35447_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_35448_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_35449_, _35448_, _35447_);
  and (_35450_, _35449_, _34581_);
  or (_35451_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_35452_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_35453_, _35452_, _35451_);
  and (_35454_, _35453_, _34796_);
  or (_35455_, _35454_, _35450_);
  or (_35456_, _35455_, _34772_);
  and (_35457_, _35456_, _34719_);
  and (_35458_, _35457_, _35446_);
  or (_35459_, _35458_, _35436_);
  and (_35460_, _35459_, _34700_);
  or (_35461_, _35460_, _35414_);
  and (_35462_, _35461_, _34840_);
  or (_35463_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_35464_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_35465_, _35464_, _35463_);
  and (_35466_, _35465_, _34581_);
  or (_35467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_35468_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_35469_, _35468_, _35467_);
  and (_35470_, _35469_, _34796_);
  or (_35471_, _35470_, _35466_);
  and (_35472_, _35471_, _34790_);
  or (_35473_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_35474_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_35475_, _35474_, _35473_);
  and (_35476_, _35475_, _34581_);
  or (_35477_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_35478_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_35479_, _35478_, _35477_);
  and (_35480_, _35479_, _34796_);
  or (_35481_, _35480_, _35476_);
  and (_35482_, _35481_, _34772_);
  or (_35483_, _35482_, _35472_);
  and (_35484_, _35483_, _34719_);
  and (_35485_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_35486_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_35487_, _35486_, _35485_);
  and (_35488_, _35487_, _34581_);
  and (_35489_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_35490_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_35491_, _35490_, _35489_);
  and (_35492_, _35491_, _34796_);
  or (_35493_, _35492_, _35488_);
  and (_35494_, _35493_, _34790_);
  and (_35495_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_35496_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_35497_, _35496_, _35495_);
  and (_35498_, _35497_, _34581_);
  and (_35499_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_35500_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_35501_, _35500_, _35499_);
  and (_35502_, _35501_, _34796_);
  or (_35503_, _35502_, _35498_);
  and (_35504_, _35503_, _34772_);
  or (_35505_, _35504_, _35494_);
  and (_35506_, _35505_, _34803_);
  or (_35507_, _35506_, _35484_);
  and (_35508_, _35507_, _34700_);
  or (_35509_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_35510_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_35511_, _35510_, _34796_);
  and (_35512_, _35511_, _35509_);
  or (_35513_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_35514_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_35515_, _35514_, _34581_);
  and (_35516_, _35515_, _35513_);
  or (_35517_, _35516_, _35512_);
  and (_35518_, _35517_, _34790_);
  or (_35519_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_35520_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_35521_, _35520_, _34796_);
  and (_35522_, _35521_, _35519_);
  or (_35523_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_35524_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_35525_, _35524_, _34581_);
  and (_35526_, _35525_, _35523_);
  or (_35527_, _35526_, _35522_);
  and (_35528_, _35527_, _34772_);
  or (_35529_, _35528_, _35518_);
  and (_35530_, _35529_, _34719_);
  and (_35531_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_35532_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_35533_, _35532_, _35531_);
  and (_35534_, _35533_, _34581_);
  and (_35535_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_35536_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_35537_, _35536_, _35535_);
  and (_35538_, _35537_, _34796_);
  or (_35539_, _35538_, _35534_);
  and (_35540_, _35539_, _34790_);
  and (_35541_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_35542_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_35543_, _35542_, _35541_);
  and (_35544_, _35543_, _34581_);
  and (_35545_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_35546_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_35547_, _35546_, _35545_);
  and (_35548_, _35547_, _34796_);
  or (_35549_, _35548_, _35544_);
  and (_35550_, _35549_, _34772_);
  or (_35551_, _35550_, _35540_);
  and (_35552_, _35551_, _34803_);
  or (_35553_, _35552_, _35530_);
  and (_35554_, _35553_, _34789_);
  or (_35555_, _35554_, _35508_);
  and (_35556_, _35555_, _34638_);
  or (_35557_, _35556_, _35462_);
  or (_35558_, _35557_, _34985_);
  and (_35559_, _35558_, _35368_);
  or (_35560_, _35559_, _35178_);
  and (_35561_, _35560_, _35177_);
  or (_35562_, _35561_, _34788_);
  not (_38997_, rst);
  not (_35563_, _34788_);
  or (_35564_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_35565_, _35564_, _38997_);
  and (_38984_[7], _35565_, _35562_);
  nor (_35566_, _34785_, _34477_);
  nor (_35567_, _34785_, _34584_);
  nor (_35568_, _35567_, _35566_);
  nor (_35569_, _34785_, _34775_);
  nor (_35570_, _34785_, _34716_);
  nor (_35571_, _35570_, _35569_);
  and (_35572_, _35571_, _35568_);
  and (_35573_, _34784_, _34701_);
  and (_35574_, _34784_, _34640_);
  nor (_35575_, _35574_, _35573_);
  nor (_35576_, _34474_, _34249_);
  and (_35577_, _35576_, _34784_);
  not (_35578_, _35577_);
  and (_35579_, _35578_, _35575_);
  and (_35580_, _35579_, _34784_);
  and (_35581_, _35580_, _35572_);
  and (_35582_, _33930_, _33898_);
  not (_35583_, _35582_);
  and (_35584_, _34197_, _34180_);
  not (_35585_, _33778_);
  nor (_35586_, _35585_, _33765_);
  not (_35587_, _33951_);
  nor (_35588_, _35587_, _33797_);
  and (_35589_, _34007_, _33883_);
  nor (_35590_, _35589_, _33967_);
  nor (_35591_, _35590_, _35588_);
  nor (_35592_, _35591_, _33916_);
  nor (_35593_, _35592_, _35586_);
  and (_35594_, _35591_, _33916_);
  nor (_35595_, _35594_, _35592_);
  not (_35596_, _35595_);
  and (_35597_, _35589_, _33967_);
  nor (_35598_, _35597_, _35590_);
  not (_35599_, _35598_);
  not (_35600_, _33991_);
  and (_35601_, _34061_, _34057_);
  and (_35602_, _35601_, _33865_);
  nor (_35603_, _34098_, _33831_);
  and (_35604_, _34131_, _33848_);
  nor (_35605_, _35604_, _34111_);
  nor (_35606_, _35605_, _35603_);
  nor (_35607_, _35606_, _34077_);
  nor (_35608_, _35607_, _35602_);
  nor (_35609_, _35608_, _34040_);
  and (_35610_, _35608_, _34040_);
  nor (_35611_, _35610_, _35609_);
  not (_35612_, _35611_);
  and (_35613_, _35606_, _34077_);
  nor (_35614_, _35613_, _35607_);
  not (_35615_, _35614_);
  and (_35616_, _35604_, _34111_);
  nor (_35617_, _35616_, _35605_);
  not (_35618_, _35617_);
  nor (_35619_, _34135_, _33734_);
  and (_35620_, _35619_, _35618_);
  and (_35621_, _35620_, _35615_);
  and (_35622_, _35621_, _35612_);
  not (_35623_, _34035_);
  or (_35624_, _35623_, _33814_);
  and (_35625_, _35623_, _33814_);
  or (_35626_, _35608_, _35625_);
  and (_35627_, _35626_, _35624_);
  or (_35628_, _35627_, _35622_);
  and (_35629_, _35628_, _35600_);
  and (_35630_, _35629_, _35599_);
  and (_35631_, _35630_, _35596_);
  nor (_35632_, _35631_, _35593_);
  nor (_35633_, _35632_, _34207_);
  nor (_35634_, _35633_, _35584_);
  nor (_35635_, _35634_, _35583_);
  not (_35636_, _35635_);
  and (_35637_, _33930_, _33906_);
  not (_35638_, _35637_);
  not (_35639_, _34207_);
  not (_35640_, _34077_);
  and (_35641_, _34134_, _34111_);
  nor (_35642_, _35641_, _34110_);
  nor (_35643_, _35642_, _35640_);
  nor (_35644_, _35643_, _34076_);
  nor (_35645_, _35644_, _34040_);
  and (_35646_, _35644_, _34040_);
  nor (_35647_, _35646_, _35645_);
  not (_35648_, _34135_);
  nor (_35649_, _35648_, _33734_);
  and (_35650_, _35649_, _34111_);
  and (_35651_, _35642_, _35640_);
  nor (_35652_, _35651_, _35643_);
  and (_35653_, _35652_, _35650_);
  not (_35654_, _35653_);
  nor (_35655_, _35654_, _35647_);
  nor (_35656_, _35644_, _34036_);
  or (_35657_, _35656_, _34038_);
  or (_35658_, _35657_, _35655_);
  and (_35659_, _35658_, _33991_);
  and (_35660_, _35659_, _33967_);
  not (_35661_, _33916_);
  and (_35662_, _33990_, _33967_);
  nor (_35663_, _35662_, _33966_);
  nor (_35664_, _35663_, _35661_);
  and (_35665_, _35663_, _35661_);
  nor (_35666_, _35665_, _35664_);
  and (_35667_, _35666_, _35660_);
  not (_35668_, _35667_);
  nor (_35669_, _35664_, _33915_);
  and (_35670_, _35669_, _35668_);
  nor (_35671_, _35670_, _35639_);
  nor (_35672_, _35671_, _34206_);
  nor (_35673_, _35672_, _35638_);
  and (_35674_, _33730_, _33728_);
  and (_35675_, _33908_, _33898_);
  and (_35676_, _33922_, _33728_);
  nor (_35677_, _35676_, _35675_);
  nor (_35678_, _35677_, _35674_);
  nor (_35679_, _33924_, _33888_);
  not (_35680_, _33733_);
  and (_35681_, _33913_, _33671_);
  nor (_35682_, _35681_, _35680_);
  nor (_35683_, _35682_, _33732_);
  not (_35684_, _35683_);
  nor (_35685_, _35684_, _35679_);
  nor (_35686_, _35685_, _35678_);
  not (_35687_, _34183_);
  and (_35688_, _33921_, _33906_);
  and (_35689_, _34064_, _33831_);
  nor (_35690_, _35689_, _33814_);
  and (_35691_, _35690_, _35688_);
  and (_35692_, _35691_, _33884_);
  nor (_35693_, _35692_, _35687_);
  and (_35694_, _35693_, _33734_);
  nor (_35695_, _35694_, _34200_);
  not (_35696_, _35688_);
  nor (_35697_, _33734_, _34180_);
  not (_35698_, _35697_);
  nor (_35699_, _35698_, _35693_);
  nor (_35700_, _35699_, _35696_);
  and (_35701_, _35700_, _35695_);
  nor (_35702_, _33733_, _33728_);
  not (_35703_, _33914_);
  nor (_35704_, _35703_, _33732_);
  nor (_35705_, _35704_, _33909_);
  nor (_35706_, _35705_, _35702_);
  not (_35707_, _34180_);
  and (_35708_, _33908_, _33673_);
  and (_35709_, _35708_, _35707_);
  and (_35710_, _33935_, _33888_);
  not (_35711_, _33848_);
  and (_35712_, _33906_, _33671_);
  and (_35713_, _35712_, _35711_);
  or (_35714_, _35691_, _35713_);
  or (_35715_, _35714_, _35710_);
  or (_35716_, _35715_, _35709_);
  or (_35717_, _35716_, _35706_);
  nor (_35718_, _35717_, _35701_);
  and (_35719_, _35718_, _35686_);
  not (_35720_, _35719_);
  nor (_35721_, _35720_, _35673_);
  and (_35722_, _35721_, _35636_);
  not (_35723_, _35722_);
  and (_35724_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _33705_);
  and (_35725_, _35724_, _33695_);
  and (_35726_, _35725_, _35723_);
  nor (_35727_, _34148_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_35728_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_35729_, _35725_, _35728_);
  and (_35730_, _35729_, _33717_);
  or (_35731_, _35730_, _35727_);
  or (_35732_, _35731_, _35726_);
  and (_35733_, _35732_, _35581_);
  not (_35734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_35735_, _35581_, _35734_);
  or (_36928_, _35735_, _35733_);
  not (_35736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_35737_, _35581_, _35736_);
  nand (_35738_, _35724_, _33690_);
  nor (_35739_, _35738_, _35722_);
  and (_35740_, _34122_, _35728_);
  and (_35741_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_35742_, _35724_, _33700_);
  or (_35743_, _35742_, _35741_);
  and (_35744_, _35724_, _33683_);
  or (_35745_, _35744_, _35743_);
  and (_35746_, _35745_, _33721_);
  or (_35747_, _35746_, _35740_);
  or (_35748_, _35747_, _35739_);
  and (_35749_, _35748_, _35581_);
  or (_36929_, _35749_, _35737_);
  nand (_35750_, _35724_, _33684_);
  nor (_35751_, _35750_, _35722_);
  and (_35752_, _34089_, _35728_);
  nand (_35753_, _33684_, _33705_);
  and (_35754_, _33708_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_35755_, _35754_, _35753_);
  or (_35756_, _35755_, _35752_);
  or (_35757_, _35756_, _35751_);
  and (_35758_, _35757_, _35581_);
  not (_35759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_35760_, _35581_, _35759_);
  or (_36930_, _35760_, _35758_);
  and (_35761_, _35742_, _35723_);
  nor (_35762_, _34052_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_35763_, _33700_, _33705_);
  and (_35764_, _33713_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_35765_, _35764_, _35763_);
  or (_35766_, _35765_, _35762_);
  or (_35767_, _35766_, _35761_);
  and (_35768_, _35767_, _35581_);
  not (_35769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_35770_, _35581_, _35769_);
  or (_36931_, _35770_, _35768_);
  nand (_35771_, _35741_, _33695_);
  nor (_35772_, _35771_, _35722_);
  nor (_35773_, _34017_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_35774_, _33695_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_35775_, _33694_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_35776_, _35775_, _35774_);
  or (_35777_, _35776_, _35773_);
  or (_35778_, _35777_, _35772_);
  and (_35779_, _35778_, _35581_);
  not (_35780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_35781_, _35581_, _35780_);
  or (_36932_, _35781_, _35779_);
  not (_35782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_35783_, _35581_, _35782_);
  nand (_35784_, _35741_, _33690_);
  nor (_35785_, _35784_, _35722_);
  and (_35786_, _33978_, _35728_);
  nand (_35787_, _33690_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_35788_, _33689_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_35789_, _35788_, _35787_);
  or (_35790_, _35789_, _35786_);
  or (_35791_, _35790_, _35785_);
  and (_35792_, _35791_, _35581_);
  or (_36933_, _35792_, _35783_);
  not (_35793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_35794_, _35581_, _35793_);
  nand (_35795_, _35741_, _33684_);
  nor (_35796_, _35795_, _35722_);
  and (_35797_, _33942_, _35728_);
  nand (_35798_, _33684_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_35799_, _33682_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_35800_, _35799_, _35798_);
  or (_35801_, _35800_, _35797_);
  or (_35802_, _35801_, _35796_);
  and (_35803_, _35802_, _35581_);
  or (_36934_, _35803_, _35794_);
  not (_35804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_35805_, _35581_, _35804_);
  and (_35806_, _35741_, _33700_);
  not (_35807_, _35806_);
  nor (_35808_, _35807_, _35722_);
  nand (_35809_, _34221_, _35728_);
  or (_35810_, _33699_, _35728_);
  and (_35811_, _35810_, _35807_);
  and (_35812_, _35811_, _35809_);
  or (_35813_, _35812_, _35808_);
  and (_35814_, _35813_, _35581_);
  or (_36935_, _35814_, _35805_);
  and (_35815_, _35732_, _34784_);
  and (_35816_, _35566_, _34584_);
  and (_35817_, _35816_, _35571_);
  and (_35818_, _35817_, _35579_);
  and (_35819_, _35818_, _35815_);
  not (_35820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_35821_, _35818_, _35820_);
  or (_37816_, _35821_, _35819_);
  and (_35822_, _35748_, _34784_);
  and (_35823_, _35818_, _35822_);
  not (_35824_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_35825_, _35818_, _35824_);
  or (_37817_, _35825_, _35823_);
  and (_35826_, _35757_, _34784_);
  and (_35827_, _35818_, _35826_);
  not (_35828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_35829_, _35818_, _35828_);
  or (_37818_, _35829_, _35827_);
  and (_35830_, _35767_, _34784_);
  and (_35831_, _35818_, _35830_);
  not (_35832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_35833_, _35818_, _35832_);
  or (_37819_, _35833_, _35831_);
  and (_35834_, _35778_, _34784_);
  and (_35835_, _35818_, _35834_);
  not (_35836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_35837_, _35818_, _35836_);
  or (_37820_, _35837_, _35835_);
  and (_35838_, _35791_, _34784_);
  and (_35839_, _35818_, _35838_);
  not (_35840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_35841_, _35818_, _35840_);
  or (_37821_, _35841_, _35839_);
  and (_35842_, _35802_, _34784_);
  and (_35843_, _35818_, _35842_);
  not (_35844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_35845_, _35818_, _35844_);
  or (_37822_, _35845_, _35843_);
  and (_35846_, _35813_, _34784_);
  and (_35847_, _35818_, _35846_);
  not (_35848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_35849_, _35818_, _35848_);
  or (_37823_, _35849_, _35847_);
  and (_35850_, _35567_, _34477_);
  and (_35851_, _35850_, _35571_);
  and (_35852_, _35851_, _35579_);
  and (_35853_, _35852_, _35815_);
  not (_35854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_35855_, _35852_, _35854_);
  or (_38360_, _35855_, _35853_);
  and (_35856_, _35852_, _35822_);
  not (_35857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_35858_, _35852_, _35857_);
  or (_38361_, _35858_, _35856_);
  and (_35859_, _35852_, _35826_);
  not (_35860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_35861_, _35852_, _35860_);
  or (_38362_, _35861_, _35859_);
  and (_35862_, _35852_, _35830_);
  not (_35863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor (_35864_, _35852_, _35863_);
  or (_38363_, _35864_, _35862_);
  and (_35865_, _35852_, _35834_);
  not (_35866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_35867_, _35852_, _35866_);
  or (_38364_, _35867_, _35865_);
  and (_35868_, _35852_, _35838_);
  not (_35869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_35870_, _35852_, _35869_);
  or (_38365_, _35870_, _35868_);
  and (_35871_, _35852_, _35842_);
  not (_35872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_35873_, _35852_, _35872_);
  or (_38366_, _35873_, _35871_);
  and (_35874_, _35852_, _35846_);
  not (_35875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_35876_, _35852_, _35875_);
  or (_38367_, _35876_, _35874_);
  and (_35877_, _35567_, _35566_);
  and (_35878_, _35877_, _35571_);
  and (_35879_, _35878_, _35579_);
  and (_35880_, _35879_, _35815_);
  not (_35881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_35882_, _35879_, _35881_);
  or (_38448_, _35882_, _35880_);
  and (_35883_, _35879_, _35822_);
  not (_35884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_35885_, _35879_, _35884_);
  or (_38449_, _35885_, _35883_);
  and (_35886_, _35879_, _35826_);
  not (_35887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_35888_, _35879_, _35887_);
  or (_38450_, _35888_, _35886_);
  and (_35889_, _35879_, _35830_);
  not (_35890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_35891_, _35879_, _35890_);
  or (_38451_, _35891_, _35889_);
  and (_35892_, _35879_, _35834_);
  not (_35893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_35894_, _35879_, _35893_);
  or (_38452_, _35894_, _35892_);
  and (_35895_, _35879_, _35838_);
  not (_35896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_35897_, _35879_, _35896_);
  or (_38453_, _35897_, _35895_);
  and (_35898_, _35879_, _35842_);
  not (_35899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_35900_, _35879_, _35899_);
  or (_38454_, _35900_, _35898_);
  and (_35901_, _35879_, _35846_);
  not (_35902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_35903_, _35879_, _35902_);
  or (_38455_, _35903_, _35901_);
  and (_35904_, _35569_, _34716_);
  and (_35905_, _35904_, _35568_);
  and (_35906_, _35905_, _35579_);
  and (_35907_, _35906_, _35815_);
  not (_35908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_35909_, _35906_, _35908_);
  or (_38536_, _35909_, _35907_);
  and (_35910_, _35906_, _35822_);
  not (_35911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_35912_, _35906_, _35911_);
  or (_38537_, _35912_, _35910_);
  and (_35913_, _35906_, _35826_);
  not (_35914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_35915_, _35906_, _35914_);
  or (_38538_, _35915_, _35913_);
  and (_35916_, _35906_, _35830_);
  not (_35917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_35918_, _35906_, _35917_);
  or (_38539_, _35918_, _35916_);
  and (_35919_, _35906_, _35834_);
  not (_35920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_35921_, _35906_, _35920_);
  or (_38540_, _35921_, _35919_);
  and (_35922_, _35906_, _35838_);
  not (_35923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_35924_, _35906_, _35923_);
  or (_38541_, _35924_, _35922_);
  and (_35925_, _35906_, _35842_);
  not (_35926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_35927_, _35906_, _35926_);
  or (_38542_, _35927_, _35925_);
  and (_35928_, _35906_, _35846_);
  not (_35929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_35930_, _35906_, _35929_);
  or (_38543_, _35930_, _35928_);
  and (_35931_, _35904_, _35816_);
  and (_35932_, _35931_, _35579_);
  and (_35933_, _35932_, _35815_);
  not (_35934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_35935_, _35932_, _35934_);
  or (_38624_, _35935_, _35933_);
  and (_35936_, _35932_, _35822_);
  not (_35937_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_35938_, _35932_, _35937_);
  or (_38625_, _35938_, _35936_);
  and (_35939_, _35932_, _35826_);
  not (_35940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_35941_, _35932_, _35940_);
  or (_38626_, _35941_, _35939_);
  and (_35942_, _35932_, _35830_);
  not (_35943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_35944_, _35932_, _35943_);
  or (_38627_, _35944_, _35942_);
  and (_35945_, _35932_, _35834_);
  not (_35946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_35947_, _35932_, _35946_);
  or (_38628_, _35947_, _35945_);
  and (_35948_, _35932_, _35838_);
  not (_35949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_35950_, _35932_, _35949_);
  or (_38629_, _35950_, _35948_);
  and (_35951_, _35932_, _35842_);
  not (_35952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_35953_, _35932_, _35952_);
  or (_38630_, _35953_, _35951_);
  and (_35954_, _35932_, _35846_);
  not (_35955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_35956_, _35932_, _35955_);
  or (_38631_, _35956_, _35954_);
  and (_35957_, _35904_, _35850_);
  and (_35958_, _35957_, _35579_);
  and (_35959_, _35958_, _35815_);
  not (_35960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_35961_, _35958_, _35960_);
  or (_38712_, _35961_, _35959_);
  and (_35962_, _35958_, _35822_);
  not (_35963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_35964_, _35958_, _35963_);
  or (_38713_, _35964_, _35962_);
  and (_35965_, _35958_, _35826_);
  not (_35966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_35967_, _35958_, _35966_);
  or (_38714_, _35967_, _35965_);
  and (_35968_, _35958_, _35830_);
  not (_35969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_35970_, _35958_, _35969_);
  or (_38715_, _35970_, _35968_);
  and (_35971_, _35958_, _35834_);
  not (_35972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_35973_, _35958_, _35972_);
  or (_38716_, _35973_, _35971_);
  and (_35974_, _35958_, _35838_);
  not (_35975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_35976_, _35958_, _35975_);
  or (_38717_, _35976_, _35974_);
  and (_35977_, _35958_, _35842_);
  not (_35978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_35979_, _35958_, _35978_);
  or (_38718_, _35979_, _35977_);
  and (_35980_, _35958_, _35846_);
  not (_35981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_35982_, _35958_, _35981_);
  or (_38719_, _35982_, _35980_);
  and (_35983_, _35904_, _35877_);
  and (_35984_, _35983_, _35579_);
  and (_35985_, _35984_, _35815_);
  not (_35986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_35987_, _35984_, _35986_);
  or (_38800_, _35987_, _35985_);
  and (_35988_, _35984_, _35822_);
  not (_35989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_35990_, _35984_, _35989_);
  or (_38801_, _35990_, _35988_);
  and (_35991_, _35984_, _35826_);
  not (_35992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_35993_, _35984_, _35992_);
  or (_38802_, _35993_, _35991_);
  and (_35994_, _35984_, _35830_);
  not (_35995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_35996_, _35984_, _35995_);
  or (_38803_, _35996_, _35994_);
  and (_35997_, _35984_, _35834_);
  not (_35998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_35999_, _35984_, _35998_);
  or (_38804_, _35999_, _35997_);
  and (_36000_, _35984_, _35838_);
  not (_36001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_36002_, _35984_, _36001_);
  or (_38805_, _36002_, _36000_);
  and (_36003_, _35984_, _35842_);
  not (_36004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_36005_, _35984_, _36004_);
  or (_38806_, _36005_, _36003_);
  and (_36006_, _35984_, _35846_);
  not (_36007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_36008_, _35984_, _36007_);
  or (_38807_, _36008_, _36006_);
  and (_36009_, _35570_, _34775_);
  and (_36010_, _36009_, _35568_);
  and (_36011_, _36010_, _35579_);
  and (_36012_, _36011_, _35815_);
  not (_36013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_36014_, _36011_, _36013_);
  or (_38888_, _36014_, _36012_);
  and (_36015_, _36011_, _35822_);
  not (_36016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_36017_, _36011_, _36016_);
  or (_38889_, _36017_, _36015_);
  and (_36018_, _36011_, _35826_);
  not (_36019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_36020_, _36011_, _36019_);
  or (_38890_, _36020_, _36018_);
  and (_36021_, _36011_, _35830_);
  not (_36022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_36023_, _36011_, _36022_);
  or (_38891_, _36023_, _36021_);
  and (_36024_, _36011_, _35834_);
  not (_36025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_36026_, _36011_, _36025_);
  or (_38892_, _36026_, _36024_);
  and (_36027_, _36011_, _35838_);
  not (_36028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_36029_, _36011_, _36028_);
  or (_38893_, _36029_, _36027_);
  and (_36030_, _36011_, _35842_);
  not (_36031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_36032_, _36011_, _36031_);
  or (_38894_, _36032_, _36030_);
  and (_36033_, _36011_, _35846_);
  not (_36034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_36035_, _36011_, _36034_);
  or (_38895_, _36035_, _36033_);
  and (_36036_, _36009_, _35816_);
  and (_36037_, _36036_, _35579_);
  and (_36038_, _36037_, _35815_);
  not (_36039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_36040_, _36037_, _36039_);
  or (_38976_, _36040_, _36038_);
  and (_36041_, _36037_, _35822_);
  not (_36042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_36043_, _36037_, _36042_);
  or (_38977_, _36043_, _36041_);
  and (_36044_, _36037_, _35826_);
  not (_36045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_36046_, _36037_, _36045_);
  or (_38978_, _36046_, _36044_);
  and (_36047_, _36037_, _35830_);
  not (_36048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_36049_, _36037_, _36048_);
  or (_38979_, _36049_, _36047_);
  and (_36050_, _36037_, _35834_);
  not (_36051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_36052_, _36037_, _36051_);
  or (_38980_, _36052_, _36050_);
  and (_36053_, _36037_, _35838_);
  not (_36054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_36055_, _36037_, _36054_);
  or (_38981_, _36055_, _36053_);
  and (_36056_, _36037_, _35842_);
  not (_36057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_36058_, _36037_, _36057_);
  or (_38982_, _36058_, _36056_);
  and (_36059_, _36037_, _35846_);
  not (_36060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_36061_, _36037_, _36060_);
  or (_38983_, _36061_, _36059_);
  and (_36062_, _36009_, _35850_);
  and (_36063_, _36062_, _35579_);
  and (_36064_, _36063_, _35815_);
  not (_36065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_36066_, _36063_, _36065_);
  or (_37016_, _36066_, _36064_);
  and (_36067_, _36063_, _35822_);
  not (_36068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_36069_, _36063_, _36068_);
  or (_37017_, _36069_, _36067_);
  and (_36070_, _36063_, _35826_);
  not (_36071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_36072_, _36063_, _36071_);
  or (_37018_, _36072_, _36070_);
  and (_36073_, _36063_, _35830_);
  not (_36074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_36075_, _36063_, _36074_);
  or (_37019_, _36075_, _36073_);
  and (_36076_, _36063_, _35834_);
  not (_36077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_36078_, _36063_, _36077_);
  or (_37020_, _36078_, _36076_);
  and (_36079_, _36063_, _35838_);
  not (_36080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_36081_, _36063_, _36080_);
  or (_37021_, _36081_, _36079_);
  and (_36082_, _36063_, _35842_);
  not (_36083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_36084_, _36063_, _36083_);
  or (_37022_, _36084_, _36082_);
  and (_36085_, _36063_, _35846_);
  not (_36086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor (_36087_, _36063_, _36086_);
  or (_37023_, _36087_, _36085_);
  and (_36088_, _36009_, _35877_);
  and (_36089_, _36088_, _35579_);
  and (_36090_, _36089_, _35815_);
  not (_36091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_36092_, _36089_, _36091_);
  or (_37104_, _36092_, _36090_);
  and (_36093_, _36089_, _35822_);
  not (_36094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_36095_, _36089_, _36094_);
  or (_37105_, _36095_, _36093_);
  and (_36096_, _36089_, _35826_);
  not (_36097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_36098_, _36089_, _36097_);
  or (_37106_, _36098_, _36096_);
  and (_36099_, _36089_, _35830_);
  not (_36100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_36101_, _36089_, _36100_);
  or (_37107_, _36101_, _36099_);
  and (_36102_, _36089_, _35834_);
  not (_36103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_36104_, _36089_, _36103_);
  or (_37108_, _36104_, _36102_);
  and (_36105_, _36089_, _35838_);
  not (_36106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_36107_, _36089_, _36106_);
  or (_37109_, _36107_, _36105_);
  and (_36108_, _36089_, _35842_);
  not (_36109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_36110_, _36089_, _36109_);
  or (_37110_, _36110_, _36108_);
  and (_36111_, _36089_, _35846_);
  not (_36112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_36113_, _36089_, _36112_);
  or (_37111_, _36113_, _36111_);
  and (_36114_, _35570_, _35569_);
  and (_36115_, _36114_, _35568_);
  and (_36116_, _36115_, _35579_);
  and (_36117_, _36116_, _35815_);
  not (_36118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_36119_, _36116_, _36118_);
  or (_37192_, _36119_, _36117_);
  and (_36120_, _36116_, _35822_);
  not (_36121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_36122_, _36116_, _36121_);
  or (_37193_, _36122_, _36120_);
  and (_36123_, _36116_, _35826_);
  not (_36124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_36125_, _36116_, _36124_);
  or (_37194_, _36125_, _36123_);
  and (_36126_, _36116_, _35830_);
  not (_36127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_36128_, _36116_, _36127_);
  or (_37195_, _36128_, _36126_);
  and (_36129_, _36116_, _35834_);
  not (_36130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_36131_, _36116_, _36130_);
  or (_37196_, _36131_, _36129_);
  and (_36132_, _36116_, _35838_);
  not (_36133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_36134_, _36116_, _36133_);
  or (_37197_, _36134_, _36132_);
  and (_36135_, _36116_, _35842_);
  not (_36136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_36137_, _36116_, _36136_);
  or (_37198_, _36137_, _36135_);
  and (_36138_, _36116_, _35846_);
  not (_36139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_36140_, _36116_, _36139_);
  or (_37199_, _36140_, _36138_);
  and (_36141_, _36114_, _35816_);
  and (_36142_, _36141_, _35579_);
  and (_36143_, _36142_, _35815_);
  not (_36144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_36145_, _36142_, _36144_);
  or (_37280_, _36145_, _36143_);
  and (_36146_, _36142_, _35822_);
  not (_36147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_36148_, _36142_, _36147_);
  or (_37281_, _36148_, _36146_);
  and (_36149_, _36142_, _35826_);
  not (_36150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_36151_, _36142_, _36150_);
  or (_37282_, _36151_, _36149_);
  and (_36152_, _36142_, _35830_);
  not (_36153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_36154_, _36142_, _36153_);
  or (_37283_, _36154_, _36152_);
  and (_36155_, _36142_, _35834_);
  not (_36156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_36157_, _36142_, _36156_);
  or (_37284_, _36157_, _36155_);
  and (_36158_, _36142_, _35838_);
  not (_36159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_36160_, _36142_, _36159_);
  or (_37285_, _36160_, _36158_);
  and (_36161_, _36142_, _35842_);
  not (_36162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_36163_, _36142_, _36162_);
  or (_37286_, _36163_, _36161_);
  and (_36164_, _36142_, _35846_);
  not (_36165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_36166_, _36142_, _36165_);
  or (_37287_, _36166_, _36164_);
  and (_36167_, _36114_, _35850_);
  and (_36168_, _36167_, _35579_);
  and (_36169_, _36168_, _35815_);
  not (_36170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_36171_, _36168_, _36170_);
  or (_37368_, _36171_, _36169_);
  and (_36172_, _36168_, _35822_);
  not (_36173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_36174_, _36168_, _36173_);
  or (_37369_, _36174_, _36172_);
  and (_36175_, _36168_, _35826_);
  not (_36176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_36177_, _36168_, _36176_);
  or (_37370_, _36177_, _36175_);
  and (_36178_, _36168_, _35830_);
  not (_36179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_36180_, _36168_, _36179_);
  or (_37371_, _36180_, _36178_);
  and (_36181_, _36168_, _35834_);
  not (_36182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_36183_, _36168_, _36182_);
  or (_37372_, _36183_, _36181_);
  and (_36184_, _36168_, _35838_);
  not (_36185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_36186_, _36168_, _36185_);
  or (_37373_, _36186_, _36184_);
  and (_36187_, _36168_, _35842_);
  not (_36188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_36189_, _36168_, _36188_);
  or (_37374_, _36189_, _36187_);
  and (_36190_, _36168_, _35846_);
  not (_36191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor (_36192_, _36168_, _36191_);
  or (_37375_, _36192_, _36190_);
  and (_36193_, _36114_, _35877_);
  and (_36194_, _36193_, _35579_);
  and (_36195_, _36194_, _35815_);
  not (_36196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_36197_, _36194_, _36196_);
  or (_37456_, _36197_, _36195_);
  and (_36198_, _36194_, _35822_);
  not (_36199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_36200_, _36194_, _36199_);
  or (_37457_, _36200_, _36198_);
  and (_36201_, _36194_, _35826_);
  not (_36202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_36203_, _36194_, _36202_);
  or (_37458_, _36203_, _36201_);
  and (_36204_, _36194_, _35830_);
  not (_36205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_36206_, _36194_, _36205_);
  or (_37459_, _36206_, _36204_);
  and (_36207_, _36194_, _35834_);
  not (_36208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_36209_, _36194_, _36208_);
  or (_37460_, _36209_, _36207_);
  and (_36210_, _36194_, _35838_);
  not (_36211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_36212_, _36194_, _36211_);
  or (_37461_, _36212_, _36210_);
  and (_36213_, _36194_, _35842_);
  not (_36214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_36215_, _36194_, _36214_);
  or (_37462_, _36215_, _36213_);
  and (_36216_, _36194_, _35846_);
  not (_36217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_36218_, _36194_, _36217_);
  or (_37463_, _36218_, _36216_);
  not (_36219_, _35576_);
  and (_36220_, _35573_, _33591_);
  and (_36221_, _36220_, _36219_);
  and (_36222_, _36221_, _35572_);
  and (_36223_, _36222_, _35815_);
  not (_36224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nor (_36225_, _36222_, _36224_);
  or (_37544_, _36225_, _36223_);
  and (_36226_, _36222_, _35822_);
  not (_36227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nor (_36228_, _36222_, _36227_);
  or (_37545_, _36228_, _36226_);
  and (_36229_, _36222_, _35826_);
  not (_36230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nor (_36231_, _36222_, _36230_);
  or (_37546_, _36231_, _36229_);
  and (_36232_, _36222_, _35830_);
  not (_36233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  nor (_36234_, _36222_, _36233_);
  or (_37547_, _36234_, _36232_);
  and (_36235_, _36222_, _35834_);
  not (_36236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nor (_36237_, _36222_, _36236_);
  or (_37548_, _36237_, _36235_);
  and (_36238_, _36222_, _35838_);
  not (_36239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  nor (_36240_, _36222_, _36239_);
  or (_37549_, _36240_, _36238_);
  and (_36241_, _36222_, _35842_);
  not (_36242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nor (_36243_, _36222_, _36242_);
  or (_37550_, _36243_, _36241_);
  and (_36244_, _36222_, _35846_);
  not (_36245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  nor (_36246_, _36222_, _36245_);
  or (_37551_, _36246_, _36244_);
  and (_36247_, _36221_, _35817_);
  and (_36248_, _36247_, _35815_);
  not (_36249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nor (_36250_, _36247_, _36249_);
  or (_37632_, _36250_, _36248_);
  and (_36251_, _36247_, _35822_);
  not (_36252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nor (_36253_, _36247_, _36252_);
  or (_37633_, _36253_, _36251_);
  and (_36254_, _36247_, _35826_);
  not (_36255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nor (_36256_, _36247_, _36255_);
  or (_37634_, _36256_, _36254_);
  and (_36257_, _36247_, _35830_);
  not (_36258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nor (_36259_, _36247_, _36258_);
  or (_37635_, _36259_, _36257_);
  and (_36260_, _36247_, _35834_);
  not (_36261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  nor (_36262_, _36247_, _36261_);
  or (_37636_, _36262_, _36260_);
  and (_36263_, _36247_, _35838_);
  not (_36264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  nor (_36265_, _36247_, _36264_);
  or (_37637_, _36265_, _36263_);
  and (_36266_, _36247_, _35842_);
  not (_36267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  nor (_36268_, _36247_, _36267_);
  or (_37638_, _36268_, _36266_);
  and (_36269_, _36247_, _35846_);
  not (_36270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  nor (_36271_, _36247_, _36270_);
  or (_37639_, _36271_, _36269_);
  and (_36272_, _36221_, _35851_);
  and (_36273_, _36272_, _35815_);
  not (_36274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  nor (_36275_, _36272_, _36274_);
  or (_37720_, _36275_, _36273_);
  and (_36276_, _36272_, _35822_);
  not (_36277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  nor (_36278_, _36272_, _36277_);
  or (_37721_, _36278_, _36276_);
  and (_36279_, _36272_, _35826_);
  not (_36280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  nor (_36281_, _36272_, _36280_);
  or (_37722_, _36281_, _36279_);
  and (_36282_, _36272_, _35830_);
  not (_36283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  nor (_36284_, _36272_, _36283_);
  or (_37723_, _36284_, _36282_);
  and (_36285_, _36272_, _35834_);
  not (_36286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nor (_36287_, _36272_, _36286_);
  or (_37724_, _36287_, _36285_);
  and (_36288_, _36272_, _35838_);
  not (_36289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  nor (_36290_, _36272_, _36289_);
  or (_37725_, _36290_, _36288_);
  and (_36291_, _36272_, _35842_);
  not (_36292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nor (_36293_, _36272_, _36292_);
  or (_37726_, _36293_, _36291_);
  and (_36294_, _36272_, _35846_);
  not (_36295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  nor (_36296_, _36272_, _36295_);
  or (_37727_, _36296_, _36294_);
  and (_36297_, _36221_, _35878_);
  and (_36298_, _36297_, _35815_);
  not (_36299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nor (_36300_, _36297_, _36299_);
  or (_37808_, _36300_, _36298_);
  and (_36301_, _36297_, _35822_);
  not (_36302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  nor (_36303_, _36297_, _36302_);
  or (_37809_, _36303_, _36301_);
  and (_36304_, _36297_, _35826_);
  not (_36305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nor (_36306_, _36297_, _36305_);
  or (_37810_, _36306_, _36304_);
  and (_36307_, _36297_, _35830_);
  not (_36308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nor (_36309_, _36297_, _36308_);
  or (_37811_, _36309_, _36307_);
  and (_36310_, _36297_, _35834_);
  not (_36311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nor (_36312_, _36297_, _36311_);
  or (_37812_, _36312_, _36310_);
  and (_36313_, _36297_, _35838_);
  not (_36314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  nor (_36315_, _36297_, _36314_);
  or (_37813_, _36315_, _36313_);
  and (_36316_, _36297_, _35842_);
  not (_36317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  nor (_36318_, _36297_, _36317_);
  or (_37814_, _36318_, _36316_);
  and (_36319_, _36297_, _35846_);
  not (_36320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  nor (_36321_, _36297_, _36320_);
  or (_37815_, _36321_, _36319_);
  and (_36322_, _36221_, _35905_);
  and (_36323_, _36322_, _35815_);
  not (_36324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  nor (_36325_, _36322_, _36324_);
  or (_37904_, _36325_, _36323_);
  and (_36326_, _36322_, _35822_);
  not (_36327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nor (_36328_, _36322_, _36327_);
  or (_37905_, _36328_, _36326_);
  and (_36329_, _36322_, _35826_);
  not (_36330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  nor (_36331_, _36322_, _36330_);
  or (_37906_, _36331_, _36329_);
  and (_36332_, _36322_, _35830_);
  not (_36333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  nor (_36334_, _36322_, _36333_);
  or (_37907_, _36334_, _36332_);
  and (_36335_, _36322_, _35834_);
  not (_36336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  nor (_36337_, _36322_, _36336_);
  or (_37908_, _36337_, _36335_);
  and (_36338_, _36322_, _35838_);
  not (_36339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  nor (_36340_, _36322_, _36339_);
  or (_37909_, _36340_, _36338_);
  and (_36341_, _36322_, _35842_);
  not (_36342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nor (_36343_, _36322_, _36342_);
  or (_37910_, _36343_, _36341_);
  and (_36344_, _36322_, _35846_);
  not (_36345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  nor (_36346_, _36322_, _36345_);
  or (_37911_, _36346_, _36344_);
  and (_36347_, _36221_, _35931_);
  and (_36348_, _36347_, _35815_);
  not (_36349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nor (_36350_, _36347_, _36349_);
  or (_37992_, _36350_, _36348_);
  and (_36351_, _36347_, _35822_);
  not (_36352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  nor (_36353_, _36347_, _36352_);
  or (_37993_, _36353_, _36351_);
  and (_36354_, _36347_, _35826_);
  not (_36355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  nor (_36356_, _36347_, _36355_);
  or (_37994_, _36356_, _36354_);
  and (_36357_, _36347_, _35830_);
  not (_36358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nor (_36359_, _36347_, _36358_);
  or (_37995_, _36359_, _36357_);
  and (_36360_, _36347_, _35834_);
  not (_36361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  nor (_36362_, _36347_, _36361_);
  or (_37996_, _36362_, _36360_);
  and (_36363_, _36347_, _35838_);
  not (_36364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  nor (_36365_, _36347_, _36364_);
  or (_37997_, _36365_, _36363_);
  and (_36366_, _36347_, _35842_);
  not (_36367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nor (_36368_, _36347_, _36367_);
  or (_37998_, _36368_, _36366_);
  and (_36369_, _36347_, _35846_);
  not (_36370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  nor (_36371_, _36347_, _36370_);
  or (_37999_, _36371_, _36369_);
  and (_36372_, _36221_, _35957_);
  and (_36373_, _36372_, _35815_);
  not (_36374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  nor (_36375_, _36372_, _36374_);
  or (_38080_, _36375_, _36373_);
  and (_36376_, _36372_, _35822_);
  not (_36377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nor (_36378_, _36372_, _36377_);
  or (_38081_, _36378_, _36376_);
  and (_36379_, _36372_, _35826_);
  not (_36380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nor (_36381_, _36372_, _36380_);
  or (_38082_, _36381_, _36379_);
  and (_36382_, _36372_, _35830_);
  not (_36383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  nor (_36384_, _36372_, _36383_);
  or (_38083_, _36384_, _36382_);
  and (_36385_, _36372_, _35834_);
  not (_36386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nor (_36387_, _36372_, _36386_);
  or (_38084_, _36387_, _36385_);
  and (_36388_, _36372_, _35838_);
  not (_36389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  nor (_36390_, _36372_, _36389_);
  or (_38085_, _36390_, _36388_);
  and (_36391_, _36372_, _35842_);
  not (_36392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  nor (_36393_, _36372_, _36392_);
  or (_38086_, _36393_, _36391_);
  and (_36394_, _36372_, _35846_);
  not (_36395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  nor (_36396_, _36372_, _36395_);
  or (_38087_, _36396_, _36394_);
  and (_36397_, _36221_, _35983_);
  and (_36398_, _36397_, _35815_);
  not (_36399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nor (_36400_, _36397_, _36399_);
  or (_38168_, _36400_, _36398_);
  and (_36401_, _36397_, _35822_);
  not (_36402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  nor (_36403_, _36397_, _36402_);
  or (_38169_, _36403_, _36401_);
  and (_36404_, _36397_, _35826_);
  not (_36405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  nor (_36406_, _36397_, _36405_);
  or (_38170_, _36406_, _36404_);
  and (_36407_, _36397_, _35830_);
  not (_36408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nor (_36409_, _36397_, _36408_);
  or (_38171_, _36409_, _36407_);
  and (_36410_, _36397_, _35834_);
  not (_36411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nor (_36412_, _36397_, _36411_);
  or (_38172_, _36412_, _36410_);
  and (_36413_, _36397_, _35838_);
  not (_36414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nor (_36415_, _36397_, _36414_);
  or (_38173_, _36415_, _36413_);
  and (_36416_, _36397_, _35842_);
  not (_36417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nor (_36418_, _36397_, _36417_);
  or (_38174_, _36418_, _36416_);
  and (_36419_, _36397_, _35846_);
  not (_36420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  nor (_36421_, _36397_, _36420_);
  or (_38175_, _36421_, _36419_);
  and (_36422_, _36221_, _36010_);
  and (_36423_, _36422_, _35815_);
  not (_36424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  nor (_36425_, _36422_, _36424_);
  or (_38256_, _36425_, _36423_);
  and (_36426_, _36422_, _35822_);
  not (_36427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor (_36428_, _36422_, _36427_);
  or (_38257_, _36428_, _36426_);
  and (_36429_, _36422_, _35826_);
  not (_36430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor (_36431_, _36422_, _36430_);
  or (_38258_, _36431_, _36429_);
  and (_36432_, _36422_, _35830_);
  not (_36433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  nor (_36434_, _36422_, _36433_);
  or (_38259_, _36434_, _36432_);
  and (_36435_, _36422_, _35834_);
  not (_36436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  nor (_36437_, _36422_, _36436_);
  or (_38260_, _36437_, _36435_);
  and (_36438_, _36422_, _35838_);
  not (_36439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  nor (_36440_, _36422_, _36439_);
  or (_38261_, _36440_, _36438_);
  and (_36441_, _36422_, _35842_);
  not (_36442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  nor (_36443_, _36422_, _36442_);
  or (_38262_, _36443_, _36441_);
  and (_36444_, _36422_, _35846_);
  not (_36445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  nor (_36446_, _36422_, _36445_);
  or (_38263_, _36446_, _36444_);
  and (_36447_, _36221_, _36036_);
  and (_36448_, _36447_, _35815_);
  not (_36449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor (_36450_, _36447_, _36449_);
  or (_38320_, _36450_, _36448_);
  and (_36451_, _36447_, _35822_);
  not (_36452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nor (_36453_, _36447_, _36452_);
  or (_38321_, _36453_, _36451_);
  and (_36454_, _36447_, _35826_);
  not (_36455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nor (_36456_, _36447_, _36455_);
  or (_38322_, _36456_, _36454_);
  and (_36457_, _36447_, _35830_);
  not (_36458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor (_36459_, _36447_, _36458_);
  or (_38323_, _36459_, _36457_);
  and (_36460_, _36447_, _35834_);
  not (_36461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor (_36462_, _36447_, _36461_);
  or (_38324_, _36462_, _36460_);
  and (_36463_, _36447_, _35838_);
  not (_36464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nor (_36465_, _36447_, _36464_);
  or (_38325_, _36465_, _36463_);
  and (_36466_, _36447_, _35842_);
  not (_36467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor (_36468_, _36447_, _36467_);
  or (_38326_, _36468_, _36466_);
  and (_36469_, _36447_, _35846_);
  not (_36470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  nor (_36471_, _36447_, _36470_);
  or (_38327_, _36471_, _36469_);
  and (_36472_, _36221_, _36062_);
  and (_36473_, _36472_, _35815_);
  not (_36474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  nor (_36475_, _36472_, _36474_);
  or (_38328_, _36475_, _36473_);
  and (_36476_, _36472_, _35822_);
  not (_36477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  nor (_36478_, _36472_, _36477_);
  or (_38329_, _36478_, _36476_);
  and (_36479_, _36472_, _35826_);
  not (_36480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  nor (_36481_, _36472_, _36480_);
  or (_38330_, _36481_, _36479_);
  and (_36482_, _36472_, _35830_);
  not (_36483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  nor (_36484_, _36472_, _36483_);
  or (_38331_, _36484_, _36482_);
  and (_36485_, _36472_, _35834_);
  not (_36486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  nor (_36487_, _36472_, _36486_);
  or (_38332_, _36487_, _36485_);
  and (_36488_, _36472_, _35838_);
  not (_36489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  nor (_36490_, _36472_, _36489_);
  or (_38333_, _36490_, _36488_);
  and (_36491_, _36472_, _35842_);
  not (_36492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  nor (_36493_, _36472_, _36492_);
  or (_38334_, _36493_, _36491_);
  and (_36494_, _36472_, _35846_);
  not (_36495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  nor (_36496_, _36472_, _36495_);
  or (_38335_, _36496_, _36494_);
  and (_36497_, _36221_, _36088_);
  and (_36498_, _36497_, _35815_);
  not (_36499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor (_36500_, _36497_, _36499_);
  or (_38336_, _36500_, _36498_);
  and (_36501_, _36497_, _35822_);
  not (_36502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  nor (_36503_, _36497_, _36502_);
  or (_38337_, _36503_, _36501_);
  and (_36504_, _36497_, _35826_);
  not (_36505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  nor (_36506_, _36497_, _36505_);
  or (_38338_, _36506_, _36504_);
  and (_36507_, _36497_, _35830_);
  not (_36508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor (_36509_, _36497_, _36508_);
  or (_38339_, _36509_, _36507_);
  and (_36510_, _36497_, _35834_);
  not (_36511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor (_36512_, _36497_, _36511_);
  or (_38340_, _36512_, _36510_);
  and (_36513_, _36497_, _35838_);
  not (_36514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  nor (_36515_, _36497_, _36514_);
  or (_38341_, _36515_, _36513_);
  and (_36516_, _36497_, _35842_);
  not (_36517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  nor (_36518_, _36497_, _36517_);
  or (_38342_, _36518_, _36516_);
  and (_36519_, _36497_, _35846_);
  not (_36520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  nor (_36521_, _36497_, _36520_);
  or (_38343_, _36521_, _36519_);
  and (_36522_, _36221_, _36115_);
  and (_36523_, _36522_, _35815_);
  not (_36524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  nor (_36525_, _36522_, _36524_);
  or (_38344_, _36525_, _36523_);
  and (_36526_, _36522_, _35822_);
  not (_36527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor (_36528_, _36522_, _36527_);
  or (_38345_, _36528_, _36526_);
  and (_36529_, _36522_, _35826_);
  not (_36530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor (_36531_, _36522_, _36530_);
  or (_38346_, _36531_, _36529_);
  and (_36532_, _36522_, _35830_);
  not (_36533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  nor (_36534_, _36522_, _36533_);
  or (_38347_, _36534_, _36532_);
  and (_36535_, _36522_, _35834_);
  not (_36536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  nor (_36537_, _36522_, _36536_);
  or (_38348_, _36537_, _36535_);
  and (_36538_, _36522_, _35838_);
  not (_36539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  nor (_36540_, _36522_, _36539_);
  or (_38349_, _36540_, _36538_);
  and (_36541_, _36522_, _35842_);
  not (_36542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor (_36543_, _36522_, _36542_);
  or (_38350_, _36543_, _36541_);
  and (_36544_, _36522_, _35846_);
  not (_36545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  nor (_36546_, _36522_, _36545_);
  or (_38351_, _36546_, _36544_);
  and (_36547_, _36221_, _36141_);
  and (_36548_, _36547_, _35815_);
  not (_36549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor (_36550_, _36547_, _36549_);
  or (_38352_, _36550_, _36548_);
  and (_36551_, _36547_, _35822_);
  not (_36552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  nor (_36553_, _36547_, _36552_);
  or (_38353_, _36553_, _36551_);
  and (_36554_, _36547_, _35826_);
  not (_36555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  nor (_36556_, _36547_, _36555_);
  or (_38354_, _36556_, _36554_);
  and (_36557_, _36547_, _35830_);
  not (_36558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor (_36559_, _36547_, _36558_);
  or (_38355_, _36559_, _36557_);
  and (_36560_, _36547_, _35834_);
  not (_36561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  nor (_36562_, _36547_, _36561_);
  or (_38356_, _36562_, _36560_);
  and (_36563_, _36547_, _35838_);
  not (_36564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor (_36565_, _36547_, _36564_);
  or (_38357_, _36565_, _36563_);
  and (_36566_, _36547_, _35842_);
  not (_36567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nor (_36568_, _36547_, _36567_);
  or (_38358_, _36568_, _36566_);
  and (_36569_, _36547_, _35846_);
  not (_36570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  nor (_36571_, _36547_, _36570_);
  or (_38359_, _36571_, _36569_);
  and (_36572_, _36221_, _36167_);
  and (_36573_, _36572_, _35815_);
  not (_36574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  nor (_36575_, _36572_, _36574_);
  or (_38368_, _36575_, _36573_);
  and (_36576_, _36572_, _35822_);
  not (_36577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor (_36578_, _36572_, _36577_);
  or (_38369_, _36578_, _36576_);
  and (_36579_, _36572_, _35826_);
  not (_36580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nor (_36581_, _36572_, _36580_);
  or (_38370_, _36581_, _36579_);
  and (_36582_, _36572_, _35830_);
  not (_36583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  nor (_36584_, _36572_, _36583_);
  or (_38371_, _36584_, _36582_);
  and (_36585_, _36572_, _35834_);
  not (_36586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor (_36587_, _36572_, _36586_);
  or (_38372_, _36587_, _36585_);
  and (_36588_, _36572_, _35838_);
  not (_36589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  nor (_36590_, _36572_, _36589_);
  or (_38373_, _36590_, _36588_);
  and (_36591_, _36572_, _35842_);
  not (_36592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  nor (_36593_, _36572_, _36592_);
  or (_38374_, _36593_, _36591_);
  and (_36594_, _36572_, _35846_);
  not (_36595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  nor (_36596_, _36572_, _36595_);
  or (_38375_, _36596_, _36594_);
  and (_36597_, _36221_, _36193_);
  and (_36598_, _36597_, _35815_);
  not (_36599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor (_36600_, _36597_, _36599_);
  or (_38376_, _36600_, _36598_);
  and (_36601_, _36597_, _35822_);
  not (_36602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor (_36603_, _36597_, _36602_);
  or (_38377_, _36603_, _36601_);
  and (_36604_, _36597_, _35826_);
  not (_36605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor (_36606_, _36597_, _36605_);
  or (_38378_, _36606_, _36604_);
  and (_36607_, _36597_, _35830_);
  not (_36608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  nor (_36609_, _36597_, _36608_);
  or (_38379_, _36609_, _36607_);
  and (_36610_, _36597_, _35834_);
  not (_36611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor (_36612_, _36597_, _36611_);
  or (_38380_, _36612_, _36610_);
  and (_36613_, _36597_, _35838_);
  not (_36614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  nor (_36615_, _36597_, _36614_);
  or (_38381_, _36615_, _36613_);
  and (_36616_, _36597_, _35842_);
  not (_36617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nor (_36618_, _36597_, _36617_);
  or (_38382_, _36618_, _36616_);
  and (_36619_, _36597_, _35846_);
  not (_36620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor (_36621_, _36597_, _36620_);
  or (_38383_, _36621_, _36619_);
  and (_36622_, _35574_, _34702_);
  and (_36623_, _36622_, _36219_);
  and (_36624_, _36623_, _35572_);
  and (_36625_, _36624_, _35815_);
  not (_36626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  nor (_36627_, _36624_, _36626_);
  or (_38384_, _36627_, _36625_);
  and (_36628_, _36624_, _35822_);
  not (_36629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  nor (_36630_, _36624_, _36629_);
  or (_38385_, _36630_, _36628_);
  and (_36631_, _36624_, _35826_);
  not (_36632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  nor (_36633_, _36624_, _36632_);
  or (_38386_, _36633_, _36631_);
  and (_36634_, _36624_, _35830_);
  not (_36635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nor (_36636_, _36624_, _36635_);
  or (_38387_, _36636_, _36634_);
  and (_36637_, _36624_, _35834_);
  not (_36638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  nor (_36639_, _36624_, _36638_);
  or (_38388_, _36639_, _36637_);
  and (_36640_, _36624_, _35838_);
  not (_36641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  nor (_36642_, _36624_, _36641_);
  or (_38389_, _36642_, _36640_);
  and (_36643_, _36624_, _35842_);
  not (_36644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  nor (_36645_, _36624_, _36644_);
  or (_38390_, _36645_, _36643_);
  and (_36646_, _36624_, _35846_);
  not (_36647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  nor (_36648_, _36624_, _36647_);
  or (_38391_, _36648_, _36646_);
  and (_36649_, _36623_, _35817_);
  and (_36650_, _36649_, _35815_);
  not (_36651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  nor (_36652_, _36649_, _36651_);
  or (_38392_, _36652_, _36650_);
  and (_36653_, _36649_, _35822_);
  not (_36654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  nor (_36655_, _36649_, _36654_);
  or (_38393_, _36655_, _36653_);
  and (_36656_, _36649_, _35826_);
  not (_36657_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nor (_36658_, _36649_, _36657_);
  or (_38394_, _36658_, _36656_);
  and (_36659_, _36649_, _35830_);
  not (_36660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nor (_36661_, _36649_, _36660_);
  or (_38395_, _36661_, _36659_);
  and (_36662_, _36649_, _35834_);
  not (_36663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  nor (_36664_, _36649_, _36663_);
  or (_38396_, _36664_, _36662_);
  and (_36665_, _36649_, _35838_);
  not (_36666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  nor (_36667_, _36649_, _36666_);
  or (_38397_, _36667_, _36665_);
  and (_36668_, _36649_, _35842_);
  not (_36669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  nor (_36670_, _36649_, _36669_);
  or (_38398_, _36670_, _36668_);
  and (_36671_, _36649_, _35846_);
  not (_36672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  nor (_36673_, _36649_, _36672_);
  or (_38399_, _36673_, _36671_);
  and (_36674_, _36623_, _35851_);
  and (_36675_, _36674_, _35815_);
  not (_36676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nor (_36677_, _36674_, _36676_);
  or (_38400_, _36677_, _36675_);
  and (_36678_, _36674_, _35822_);
  not (_36679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nor (_36680_, _36674_, _36679_);
  or (_38401_, _36680_, _36678_);
  and (_36681_, _36674_, _35826_);
  not (_36682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  nor (_36683_, _36674_, _36682_);
  or (_38402_, _36683_, _36681_);
  and (_36684_, _36674_, _35830_);
  not (_36685_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  nor (_36686_, _36674_, _36685_);
  or (_38403_, _36686_, _36684_);
  and (_36687_, _36674_, _35834_);
  not (_36688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nor (_36689_, _36674_, _36688_);
  or (_38404_, _36689_, _36687_);
  and (_36690_, _36674_, _35838_);
  not (_36691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  nor (_36692_, _36674_, _36691_);
  or (_38405_, _36692_, _36690_);
  and (_36693_, _36674_, _35842_);
  not (_36694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nor (_36695_, _36674_, _36694_);
  or (_38406_, _36695_, _36693_);
  and (_36696_, _36674_, _35846_);
  not (_36697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  nor (_36698_, _36674_, _36697_);
  or (_38407_, _36698_, _36696_);
  and (_36699_, _36623_, _35878_);
  and (_36700_, _36699_, _35815_);
  not (_36701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nor (_36702_, _36699_, _36701_);
  or (_38408_, _36702_, _36700_);
  and (_36703_, _36699_, _35822_);
  not (_36704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nor (_36705_, _36699_, _36704_);
  or (_38409_, _36705_, _36703_);
  and (_36706_, _36699_, _35826_);
  not (_36707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nor (_36708_, _36699_, _36707_);
  or (_38410_, _36708_, _36706_);
  and (_36709_, _36699_, _35830_);
  not (_36710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  nor (_36711_, _36699_, _36710_);
  or (_38411_, _36711_, _36709_);
  and (_36712_, _36699_, _35834_);
  not (_36713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  nor (_36714_, _36699_, _36713_);
  or (_38412_, _36714_, _36712_);
  and (_36715_, _36699_, _35838_);
  not (_36716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  nor (_36717_, _36699_, _36716_);
  or (_38413_, _36717_, _36715_);
  and (_36718_, _36699_, _35842_);
  not (_36719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nor (_36720_, _36699_, _36719_);
  or (_38414_, _36720_, _36718_);
  and (_36721_, _36699_, _35846_);
  not (_36722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  nor (_36723_, _36699_, _36722_);
  or (_38415_, _36723_, _36721_);
  and (_36724_, _36623_, _35905_);
  and (_36725_, _36724_, _35815_);
  not (_36726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  nor (_36727_, _36724_, _36726_);
  or (_38416_, _36727_, _36725_);
  and (_36728_, _36724_, _35822_);
  not (_00009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  nor (_00010_, _36724_, _00009_);
  or (_38417_, _00010_, _36728_);
  and (_00011_, _36724_, _35826_);
  not (_00012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  nor (_00013_, _36724_, _00012_);
  or (_38418_, _00013_, _00011_);
  and (_00014_, _36724_, _35830_);
  not (_00015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nor (_00016_, _36724_, _00015_);
  or (_38419_, _00016_, _00014_);
  and (_00017_, _36724_, _35834_);
  not (_00018_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nor (_00019_, _36724_, _00018_);
  or (_38420_, _00019_, _00017_);
  and (_00020_, _36724_, _35838_);
  not (_00021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  nor (_00022_, _36724_, _00021_);
  or (_38421_, _00022_, _00020_);
  and (_00023_, _36724_, _35842_);
  not (_00024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  nor (_00025_, _36724_, _00024_);
  or (_38422_, _00025_, _00023_);
  and (_00026_, _36724_, _35846_);
  not (_00027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  nor (_00028_, _36724_, _00027_);
  or (_38423_, _00028_, _00026_);
  and (_00029_, _36623_, _35931_);
  and (_00030_, _00029_, _35815_);
  not (_00031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  nor (_00032_, _00029_, _00031_);
  or (_38424_, _00032_, _00030_);
  and (_00033_, _00029_, _35822_);
  not (_00034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nor (_00035_, _00029_, _00034_);
  or (_38425_, _00035_, _00033_);
  and (_00036_, _00029_, _35826_);
  not (_00037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  nor (_00038_, _00029_, _00037_);
  or (_38426_, _00038_, _00036_);
  and (_00039_, _00029_, _35830_);
  not (_00040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nor (_00041_, _00029_, _00040_);
  or (_38427_, _00041_, _00039_);
  and (_00042_, _00029_, _35834_);
  not (_00043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  nor (_00044_, _00029_, _00043_);
  or (_38428_, _00044_, _00042_);
  and (_00045_, _00029_, _35838_);
  not (_00046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  nor (_00047_, _00029_, _00046_);
  or (_38429_, _00047_, _00045_);
  and (_00048_, _00029_, _35842_);
  not (_00049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  nor (_00050_, _00029_, _00049_);
  or (_38430_, _00050_, _00048_);
  and (_00051_, _00029_, _35846_);
  not (_00052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  nor (_00053_, _00029_, _00052_);
  or (_38431_, _00053_, _00051_);
  and (_00054_, _36623_, _35957_);
  and (_00055_, _00054_, _35815_);
  not (_00056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nor (_00057_, _00054_, _00056_);
  or (_38432_, _00057_, _00055_);
  and (_00058_, _00054_, _35822_);
  not (_00059_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  nor (_00060_, _00054_, _00059_);
  or (_38433_, _00060_, _00058_);
  and (_00061_, _00054_, _35826_);
  not (_00062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nor (_00063_, _00054_, _00062_);
  or (_38434_, _00063_, _00061_);
  and (_00064_, _00054_, _35830_);
  not (_00065_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  nor (_00066_, _00054_, _00065_);
  or (_38435_, _00066_, _00064_);
  and (_00067_, _00054_, _35834_);
  not (_00068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nor (_00069_, _00054_, _00068_);
  or (_38436_, _00069_, _00067_);
  and (_00070_, _00054_, _35838_);
  not (_00071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  nor (_00072_, _00054_, _00071_);
  or (_38437_, _00072_, _00070_);
  and (_00073_, _00054_, _35842_);
  not (_00074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nor (_00075_, _00054_, _00074_);
  or (_38438_, _00075_, _00073_);
  and (_00076_, _00054_, _35846_);
  not (_00077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  nor (_00078_, _00054_, _00077_);
  or (_38439_, _00078_, _00076_);
  and (_00079_, _36623_, _35983_);
  and (_00080_, _00079_, _35815_);
  not (_00081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nor (_00082_, _00079_, _00081_);
  or (_38440_, _00082_, _00080_);
  and (_00083_, _00079_, _35822_);
  not (_00084_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nor (_00085_, _00079_, _00084_);
  or (_38441_, _00085_, _00083_);
  and (_00086_, _00079_, _35826_);
  not (_00087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  nor (_00088_, _00079_, _00087_);
  or (_38442_, _00088_, _00086_);
  and (_00089_, _00079_, _35830_);
  not (_00090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nor (_00091_, _00079_, _00090_);
  or (_38443_, _00091_, _00089_);
  and (_00092_, _00079_, _35834_);
  not (_00093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  nor (_00094_, _00079_, _00093_);
  or (_38444_, _00094_, _00092_);
  and (_00095_, _00079_, _35838_);
  not (_00096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  nor (_00097_, _00079_, _00096_);
  or (_38445_, _00097_, _00095_);
  and (_00098_, _00079_, _35842_);
  not (_00099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nor (_00100_, _00079_, _00099_);
  or (_38446_, _00100_, _00098_);
  and (_00101_, _00079_, _35846_);
  not (_00102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  nor (_00103_, _00079_, _00102_);
  or (_38447_, _00103_, _00101_);
  and (_00104_, _36623_, _36010_);
  and (_00105_, _00104_, _35815_);
  not (_00106_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  nor (_00107_, _00104_, _00106_);
  or (_38456_, _00107_, _00105_);
  and (_00108_, _00104_, _35822_);
  not (_00109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  nor (_00110_, _00104_, _00109_);
  or (_38457_, _00110_, _00108_);
  and (_00111_, _00104_, _35826_);
  not (_00112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nor (_00113_, _00104_, _00112_);
  or (_38458_, _00113_, _00111_);
  and (_00114_, _00104_, _35830_);
  not (_00115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  nor (_00116_, _00104_, _00115_);
  or (_38459_, _00116_, _00114_);
  and (_00117_, _00104_, _35834_);
  not (_00118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nor (_00119_, _00104_, _00118_);
  or (_38460_, _00119_, _00117_);
  and (_00120_, _00104_, _35838_);
  not (_00121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  nor (_00122_, _00104_, _00121_);
  or (_38461_, _00122_, _00120_);
  and (_00123_, _00104_, _35842_);
  not (_00124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  nor (_00125_, _00104_, _00124_);
  or (_38462_, _00125_, _00123_);
  and (_00126_, _00104_, _35846_);
  not (_00127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  nor (_00128_, _00104_, _00127_);
  or (_38463_, _00128_, _00126_);
  and (_00129_, _36623_, _36036_);
  and (_00130_, _00129_, _35815_);
  not (_00131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  nor (_00132_, _00129_, _00131_);
  or (_38464_, _00132_, _00130_);
  and (_00133_, _00129_, _35822_);
  not (_00134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  nor (_00135_, _00129_, _00134_);
  or (_38465_, _00135_, _00133_);
  and (_00136_, _00129_, _35826_);
  not (_00137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  nor (_00138_, _00129_, _00137_);
  or (_38466_, _00138_, _00136_);
  and (_00139_, _00129_, _35830_);
  not (_00140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  nor (_00141_, _00129_, _00140_);
  or (_38467_, _00141_, _00139_);
  and (_00142_, _00129_, _35834_);
  not (_00143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nor (_00144_, _00129_, _00143_);
  or (_38468_, _00144_, _00142_);
  and (_00145_, _00129_, _35838_);
  not (_00146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  nor (_00147_, _00129_, _00146_);
  or (_38469_, _00147_, _00145_);
  and (_00148_, _00129_, _35842_);
  not (_00149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nor (_00150_, _00129_, _00149_);
  or (_38470_, _00150_, _00148_);
  and (_00151_, _00129_, _35846_);
  not (_00152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  nor (_00153_, _00129_, _00152_);
  or (_38471_, _00153_, _00151_);
  and (_00154_, _36623_, _36062_);
  and (_00155_, _00154_, _35815_);
  not (_00156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor (_00157_, _00154_, _00156_);
  or (_38472_, _00157_, _00155_);
  and (_00158_, _00154_, _35822_);
  not (_00159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nor (_00160_, _00154_, _00159_);
  or (_38473_, _00160_, _00158_);
  and (_00161_, _00154_, _35826_);
  not (_00162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor (_00163_, _00154_, _00162_);
  or (_38474_, _00163_, _00161_);
  and (_00164_, _00154_, _35830_);
  not (_00165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor (_00166_, _00154_, _00165_);
  or (_38475_, _00166_, _00164_);
  and (_00167_, _00154_, _35834_);
  not (_00168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  nor (_00169_, _00154_, _00168_);
  or (_38476_, _00169_, _00167_);
  and (_00170_, _00154_, _35838_);
  not (_00171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  nor (_00172_, _00154_, _00171_);
  or (_38477_, _00172_, _00170_);
  and (_00173_, _00154_, _35842_);
  not (_00174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  nor (_00175_, _00154_, _00174_);
  or (_38478_, _00175_, _00173_);
  and (_00176_, _00154_, _35846_);
  not (_00177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  nor (_00178_, _00154_, _00177_);
  or (_38479_, _00178_, _00176_);
  and (_00179_, _36623_, _36088_);
  and (_00180_, _00179_, _35815_);
  not (_00181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor (_00182_, _00179_, _00181_);
  or (_38480_, _00182_, _00180_);
  and (_00183_, _00179_, _35822_);
  not (_00184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor (_00185_, _00179_, _00184_);
  or (_38481_, _00185_, _00183_);
  and (_00186_, _00179_, _35826_);
  not (_00187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor (_00188_, _00179_, _00187_);
  or (_38482_, _00188_, _00186_);
  and (_00189_, _00179_, _35830_);
  not (_00190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  nor (_00191_, _00179_, _00190_);
  or (_38483_, _00191_, _00189_);
  and (_00192_, _00179_, _35834_);
  not (_00193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  nor (_00194_, _00179_, _00193_);
  or (_38484_, _00194_, _00192_);
  and (_00195_, _00179_, _35838_);
  not (_00196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  nor (_00197_, _00179_, _00196_);
  or (_38485_, _00197_, _00195_);
  and (_00198_, _00179_, _35842_);
  not (_00199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  nor (_00200_, _00179_, _00199_);
  or (_38486_, _00200_, _00198_);
  and (_00201_, _00179_, _35846_);
  not (_00202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  nor (_00203_, _00179_, _00202_);
  or (_38487_, _00203_, _00201_);
  and (_00204_, _36623_, _36115_);
  and (_00205_, _00204_, _35815_);
  not (_00206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  nor (_00207_, _00204_, _00206_);
  or (_38488_, _00207_, _00205_);
  and (_00208_, _00204_, _35822_);
  not (_00209_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  nor (_00210_, _00204_, _00209_);
  or (_38489_, _00210_, _00208_);
  and (_00211_, _00204_, _35826_);
  not (_00212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  nor (_00213_, _00204_, _00212_);
  or (_38490_, _00213_, _00211_);
  and (_00214_, _00204_, _35830_);
  not (_00215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nor (_00216_, _00204_, _00215_);
  or (_38491_, _00216_, _00214_);
  and (_00217_, _00204_, _35834_);
  not (_00218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nor (_00219_, _00204_, _00218_);
  or (_38492_, _00219_, _00217_);
  and (_00220_, _00204_, _35838_);
  not (_00221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  nor (_00222_, _00204_, _00221_);
  or (_38493_, _00222_, _00220_);
  and (_00223_, _00204_, _35842_);
  not (_00224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nor (_00225_, _00204_, _00224_);
  or (_38494_, _00225_, _00223_);
  and (_00226_, _00204_, _35846_);
  not (_00227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  nor (_00228_, _00204_, _00227_);
  or (_38495_, _00228_, _00226_);
  and (_00229_, _36623_, _36141_);
  and (_00230_, _00229_, _35815_);
  not (_00231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  nor (_00232_, _00229_, _00231_);
  or (_38496_, _00232_, _00230_);
  and (_00233_, _00229_, _35822_);
  not (_00234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nor (_00235_, _00229_, _00234_);
  or (_38497_, _00235_, _00233_);
  and (_00236_, _00229_, _35826_);
  not (_00237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nor (_00238_, _00229_, _00237_);
  or (_38498_, _00238_, _00236_);
  and (_00239_, _00229_, _35830_);
  not (_00240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  nor (_00241_, _00229_, _00240_);
  or (_38499_, _00241_, _00239_);
  and (_00242_, _00229_, _35834_);
  not (_00243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  nor (_00244_, _00229_, _00243_);
  or (_38500_, _00244_, _00242_);
  and (_00245_, _00229_, _35838_);
  not (_00246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  nor (_00247_, _00229_, _00246_);
  or (_38501_, _00247_, _00245_);
  and (_00248_, _00229_, _35842_);
  not (_00249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nor (_00250_, _00229_, _00249_);
  or (_38502_, _00250_, _00248_);
  and (_00251_, _00229_, _35846_);
  not (_00252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  nor (_00253_, _00229_, _00252_);
  or (_38503_, _00253_, _00251_);
  and (_00254_, _36623_, _36167_);
  and (_00255_, _00254_, _35815_);
  not (_00256_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor (_00257_, _00254_, _00256_);
  or (_38504_, _00257_, _00255_);
  and (_00258_, _00254_, _35822_);
  not (_00259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  nor (_00260_, _00254_, _00259_);
  or (_38505_, _00260_, _00258_);
  and (_00261_, _00254_, _35826_);
  not (_00262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  nor (_00263_, _00254_, _00262_);
  or (_38506_, _00263_, _00261_);
  and (_00264_, _00254_, _35830_);
  not (_00265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor (_00266_, _00254_, _00265_);
  or (_38507_, _00266_, _00264_);
  and (_00267_, _00254_, _35834_);
  not (_00268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor (_00269_, _00254_, _00268_);
  or (_38508_, _00269_, _00267_);
  and (_00270_, _00254_, _35838_);
  not (_00271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  nor (_00272_, _00254_, _00271_);
  or (_38509_, _00272_, _00270_);
  and (_00273_, _00254_, _35842_);
  not (_00274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  nor (_00275_, _00254_, _00274_);
  or (_38510_, _00275_, _00273_);
  and (_00276_, _00254_, _35846_);
  not (_00277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  nor (_00278_, _00254_, _00277_);
  or (_38511_, _00278_, _00276_);
  and (_00279_, _36623_, _36193_);
  and (_00280_, _00279_, _35815_);
  not (_00281_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  nor (_00282_, _00279_, _00281_);
  or (_38512_, _00282_, _00280_);
  and (_00283_, _00279_, _35822_);
  not (_00284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor (_00285_, _00279_, _00284_);
  or (_38513_, _00285_, _00283_);
  and (_00286_, _00279_, _35826_);
  not (_00287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  nor (_00288_, _00279_, _00287_);
  or (_38514_, _00288_, _00286_);
  and (_00289_, _00279_, _35830_);
  not (_00290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor (_00291_, _00279_, _00290_);
  or (_38515_, _00291_, _00289_);
  and (_00292_, _00279_, _35834_);
  not (_00293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor (_00294_, _00279_, _00293_);
  or (_38516_, _00294_, _00292_);
  and (_00295_, _00279_, _35838_);
  not (_00296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  nor (_00297_, _00279_, _00296_);
  or (_38517_, _00297_, _00295_);
  and (_00298_, _00279_, _35842_);
  not (_00299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  nor (_00300_, _00279_, _00299_);
  or (_38518_, _00300_, _00298_);
  and (_00301_, _00279_, _35846_);
  not (_00302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  nor (_00303_, _00279_, _00302_);
  or (_38519_, _00303_, _00301_);
  and (_00304_, _35573_, _34640_);
  and (_00305_, _00304_, _36219_);
  and (_00306_, _00305_, _35572_);
  and (_00307_, _00306_, _35815_);
  not (_00308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nor (_00309_, _00306_, _00308_);
  or (_38520_, _00309_, _00307_);
  and (_00310_, _00306_, _35822_);
  not (_00311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  nor (_00312_, _00306_, _00311_);
  or (_38521_, _00312_, _00310_);
  and (_00313_, _00306_, _35826_);
  not (_00314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nor (_00315_, _00306_, _00314_);
  or (_38522_, _00315_, _00313_);
  and (_00316_, _00306_, _35830_);
  not (_00317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  nor (_00318_, _00306_, _00317_);
  or (_38523_, _00318_, _00316_);
  and (_00319_, _00306_, _35834_);
  not (_00320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  nor (_00321_, _00306_, _00320_);
  or (_38524_, _00321_, _00319_);
  and (_00322_, _00306_, _35838_);
  not (_00323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  nor (_00324_, _00306_, _00323_);
  or (_38525_, _00324_, _00322_);
  and (_00325_, _00306_, _35842_);
  not (_00326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nor (_00327_, _00306_, _00326_);
  or (_38526_, _00327_, _00325_);
  and (_00328_, _00306_, _35846_);
  not (_00329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  nor (_00330_, _00306_, _00329_);
  or (_38527_, _00330_, _00328_);
  and (_00331_, _00305_, _35817_);
  and (_00332_, _00331_, _35815_);
  not (_00333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nor (_00334_, _00331_, _00333_);
  or (_38528_, _00334_, _00332_);
  and (_00335_, _00331_, _35822_);
  not (_00336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nor (_00337_, _00331_, _00336_);
  or (_38529_, _00337_, _00335_);
  and (_00338_, _00331_, _35826_);
  not (_00339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nor (_00340_, _00331_, _00339_);
  or (_38530_, _00340_, _00338_);
  and (_00341_, _00331_, _35830_);
  not (_00342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nor (_00343_, _00331_, _00342_);
  or (_38531_, _00343_, _00341_);
  and (_00344_, _00331_, _35834_);
  not (_00345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nor (_00346_, _00331_, _00345_);
  or (_38532_, _00346_, _00344_);
  and (_00347_, _00331_, _35838_);
  not (_00348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  nor (_00349_, _00331_, _00348_);
  or (_38533_, _00349_, _00347_);
  and (_00350_, _00331_, _35842_);
  not (_00351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nor (_00352_, _00331_, _00351_);
  or (_38534_, _00352_, _00350_);
  and (_00353_, _00331_, _35846_);
  not (_00354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  nor (_00355_, _00331_, _00354_);
  or (_38535_, _00355_, _00353_);
  and (_00356_, _00305_, _35851_);
  and (_00357_, _00356_, _35815_);
  not (_00358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  nor (_00359_, _00356_, _00358_);
  or (_38544_, _00359_, _00357_);
  and (_00360_, _00356_, _35822_);
  not (_00361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  nor (_00362_, _00356_, _00361_);
  or (_38545_, _00362_, _00360_);
  and (_00363_, _00356_, _35826_);
  not (_00364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  nor (_00365_, _00356_, _00364_);
  or (_38546_, _00365_, _00363_);
  and (_00366_, _00356_, _35830_);
  not (_00367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  nor (_00368_, _00356_, _00367_);
  or (_38547_, _00368_, _00366_);
  and (_00369_, _00356_, _35834_);
  not (_00370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  nor (_00371_, _00356_, _00370_);
  or (_38548_, _00371_, _00369_);
  and (_00372_, _00356_, _35838_);
  not (_00373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  nor (_00374_, _00356_, _00373_);
  or (_38549_, _00374_, _00372_);
  and (_00375_, _00356_, _35842_);
  not (_00376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  nor (_00377_, _00356_, _00376_);
  or (_38550_, _00377_, _00375_);
  and (_00378_, _00356_, _35846_);
  not (_00379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  nor (_00380_, _00356_, _00379_);
  or (_38551_, _00380_, _00378_);
  and (_00381_, _00305_, _35878_);
  and (_00382_, _00381_, _35815_);
  not (_00383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nor (_00384_, _00381_, _00383_);
  or (_38552_, _00384_, _00382_);
  and (_00385_, _00381_, _35822_);
  not (_00386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nor (_00387_, _00381_, _00386_);
  or (_38553_, _00387_, _00385_);
  and (_00388_, _00381_, _35826_);
  not (_00389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  nor (_00390_, _00381_, _00389_);
  or (_38554_, _00390_, _00388_);
  and (_00391_, _00381_, _35830_);
  not (_00392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  nor (_00393_, _00381_, _00392_);
  or (_38555_, _00393_, _00391_);
  and (_00394_, _00381_, _35834_);
  not (_00395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nor (_00396_, _00381_, _00395_);
  or (_38556_, _00396_, _00394_);
  and (_00397_, _00381_, _35838_);
  not (_00398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  nor (_00399_, _00381_, _00398_);
  or (_38557_, _00399_, _00397_);
  and (_00400_, _00381_, _35842_);
  not (_00401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  nor (_00402_, _00381_, _00401_);
  or (_38558_, _00402_, _00400_);
  and (_00403_, _00381_, _35846_);
  not (_00404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  nor (_00405_, _00381_, _00404_);
  or (_38559_, _00405_, _00403_);
  and (_00406_, _00305_, _35905_);
  and (_00407_, _00406_, _35815_);
  not (_00408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  nor (_00409_, _00406_, _00408_);
  or (_38560_, _00409_, _00407_);
  and (_00410_, _00406_, _35822_);
  not (_00411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  nor (_00412_, _00406_, _00411_);
  or (_38561_, _00412_, _00410_);
  and (_00413_, _00406_, _35826_);
  not (_00414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nor (_00415_, _00406_, _00414_);
  or (_38562_, _00415_, _00413_);
  and (_00416_, _00406_, _35830_);
  not (_00417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nor (_00418_, _00406_, _00417_);
  or (_38563_, _00418_, _00416_);
  and (_00419_, _00406_, _35834_);
  not (_00420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  nor (_00421_, _00406_, _00420_);
  or (_38564_, _00421_, _00419_);
  and (_00422_, _00406_, _35838_);
  not (_00423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  nor (_00424_, _00406_, _00423_);
  or (_38565_, _00424_, _00422_);
  and (_00425_, _00406_, _35842_);
  not (_00426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nor (_00427_, _00406_, _00426_);
  or (_38566_, _00427_, _00425_);
  and (_00428_, _00406_, _35846_);
  not (_00429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  nor (_00430_, _00406_, _00429_);
  or (_38567_, _00430_, _00428_);
  and (_00431_, _00305_, _35931_);
  and (_00432_, _00431_, _35815_);
  not (_00433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nor (_00434_, _00431_, _00433_);
  or (_38568_, _00434_, _00432_);
  and (_00435_, _00431_, _35822_);
  not (_00436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nor (_00437_, _00431_, _00436_);
  or (_38569_, _00437_, _00435_);
  and (_00438_, _00431_, _35826_);
  not (_00439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  nor (_00440_, _00431_, _00439_);
  or (_38570_, _00440_, _00438_);
  and (_00441_, _00431_, _35830_);
  not (_00442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  nor (_00443_, _00431_, _00442_);
  or (_38571_, _00443_, _00441_);
  and (_00444_, _00431_, _35834_);
  not (_00445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  nor (_00446_, _00431_, _00445_);
  or (_38572_, _00446_, _00444_);
  and (_00447_, _00431_, _35838_);
  not (_00448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  nor (_00449_, _00431_, _00448_);
  or (_38573_, _00449_, _00447_);
  and (_00450_, _00431_, _35842_);
  not (_00451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nor (_00452_, _00431_, _00451_);
  or (_38574_, _00452_, _00450_);
  and (_00453_, _00431_, _35846_);
  not (_00454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  nor (_00455_, _00431_, _00454_);
  or (_38575_, _00455_, _00453_);
  and (_00456_, _00305_, _35957_);
  and (_00457_, _00456_, _35815_);
  not (_00458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  nor (_00459_, _00456_, _00458_);
  or (_38576_, _00459_, _00457_);
  and (_00460_, _00456_, _35822_);
  not (_00461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  nor (_00462_, _00456_, _00461_);
  or (_38577_, _00462_, _00460_);
  and (_00463_, _00456_, _35826_);
  not (_00464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nor (_00465_, _00456_, _00464_);
  or (_38578_, _00465_, _00463_);
  and (_00466_, _00456_, _35830_);
  not (_00467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nor (_00468_, _00456_, _00467_);
  or (_38579_, _00468_, _00466_);
  and (_00469_, _00456_, _35834_);
  not (_00470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nor (_00471_, _00456_, _00470_);
  or (_38580_, _00471_, _00469_);
  and (_00472_, _00456_, _35838_);
  not (_00473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  nor (_00474_, _00456_, _00473_);
  or (_38581_, _00474_, _00472_);
  and (_00475_, _00456_, _35842_);
  not (_00476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  nor (_00477_, _00456_, _00476_);
  or (_38582_, _00477_, _00475_);
  and (_00478_, _00456_, _35846_);
  not (_00479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  nor (_00480_, _00456_, _00479_);
  or (_38583_, _00480_, _00478_);
  and (_00481_, _00305_, _35983_);
  and (_00482_, _00481_, _35815_);
  not (_00483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  nor (_00484_, _00481_, _00483_);
  or (_38584_, _00484_, _00482_);
  and (_00485_, _00481_, _35822_);
  not (_00486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nor (_00487_, _00481_, _00486_);
  or (_38585_, _00487_, _00485_);
  and (_00488_, _00481_, _35826_);
  not (_00489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  nor (_00490_, _00481_, _00489_);
  or (_38586_, _00490_, _00488_);
  and (_00491_, _00481_, _35830_);
  not (_00492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nor (_00493_, _00481_, _00492_);
  or (_38587_, _00493_, _00491_);
  and (_00494_, _00481_, _35834_);
  not (_00495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nor (_00496_, _00481_, _00495_);
  or (_38588_, _00496_, _00494_);
  and (_00497_, _00481_, _35838_);
  not (_00498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nor (_00499_, _00481_, _00498_);
  or (_38589_, _00499_, _00497_);
  and (_00500_, _00481_, _35842_);
  not (_00501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nor (_00502_, _00481_, _00501_);
  or (_38590_, _00502_, _00500_);
  and (_00503_, _00481_, _35846_);
  not (_00504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  nor (_00505_, _00481_, _00504_);
  or (_38591_, _00505_, _00503_);
  and (_00506_, _00305_, _36010_);
  and (_00507_, _00506_, _35815_);
  not (_00508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor (_00509_, _00506_, _00508_);
  or (_38592_, _00509_, _00507_);
  and (_00510_, _00506_, _35822_);
  not (_00511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  nor (_00512_, _00506_, _00511_);
  or (_38593_, _00512_, _00510_);
  and (_00513_, _00506_, _35826_);
  not (_00514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nor (_00515_, _00506_, _00514_);
  or (_38594_, _00515_, _00513_);
  and (_00516_, _00506_, _35830_);
  not (_00517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  nor (_00518_, _00506_, _00517_);
  or (_38595_, _00518_, _00516_);
  and (_00519_, _00506_, _35834_);
  not (_00520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  nor (_00521_, _00506_, _00520_);
  or (_38596_, _00521_, _00519_);
  and (_00522_, _00506_, _35838_);
  not (_00523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  nor (_00524_, _00506_, _00523_);
  or (_38597_, _00524_, _00522_);
  and (_00525_, _00506_, _35842_);
  not (_00526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  nor (_00527_, _00506_, _00526_);
  or (_38598_, _00527_, _00525_);
  and (_00528_, _00506_, _35846_);
  not (_00529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  nor (_00530_, _00506_, _00529_);
  or (_38599_, _00530_, _00528_);
  and (_00531_, _00305_, _36036_);
  and (_00532_, _00531_, _35815_);
  not (_00533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor (_00534_, _00531_, _00533_);
  or (_38600_, _00534_, _00532_);
  and (_00535_, _00531_, _35822_);
  not (_00536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor (_00537_, _00531_, _00536_);
  or (_38601_, _00537_, _00535_);
  and (_00538_, _00531_, _35826_);
  not (_00539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nor (_00540_, _00531_, _00539_);
  or (_38602_, _00540_, _00538_);
  and (_00541_, _00531_, _35830_);
  not (_00542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor (_00543_, _00531_, _00542_);
  or (_38603_, _00543_, _00541_);
  and (_00544_, _00531_, _35834_);
  not (_00545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  nor (_00546_, _00531_, _00545_);
  or (_38604_, _00546_, _00544_);
  and (_00547_, _00531_, _35838_);
  not (_00548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  nor (_00549_, _00531_, _00548_);
  or (_38605_, _00549_, _00547_);
  and (_00550_, _00531_, _35842_);
  not (_00551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor (_00552_, _00531_, _00551_);
  or (_38606_, _00552_, _00550_);
  and (_00553_, _00531_, _35846_);
  not (_00554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  nor (_00555_, _00531_, _00554_);
  or (_38607_, _00555_, _00553_);
  and (_00556_, _00305_, _36062_);
  and (_00557_, _00556_, _35815_);
  not (_00558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  nor (_00559_, _00556_, _00558_);
  or (_38608_, _00559_, _00557_);
  and (_00560_, _00556_, _35822_);
  not (_00561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  nor (_00562_, _00556_, _00561_);
  or (_38609_, _00562_, _00560_);
  and (_00563_, _00556_, _35826_);
  not (_00564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  nor (_00565_, _00556_, _00564_);
  or (_38610_, _00565_, _00563_);
  and (_00566_, _00556_, _35830_);
  not (_00567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  nor (_00568_, _00556_, _00567_);
  or (_38611_, _00568_, _00566_);
  and (_00569_, _00556_, _35834_);
  not (_00570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor (_00571_, _00556_, _00570_);
  or (_38612_, _00571_, _00569_);
  and (_00572_, _00556_, _35838_);
  not (_00573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  nor (_00574_, _00556_, _00573_);
  or (_38613_, _00574_, _00572_);
  and (_00575_, _00556_, _35842_);
  not (_00576_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  nor (_00577_, _00556_, _00576_);
  or (_38614_, _00577_, _00575_);
  and (_00578_, _00556_, _35846_);
  not (_00579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  nor (_00580_, _00556_, _00579_);
  or (_38615_, _00580_, _00578_);
  and (_00581_, _00305_, _36088_);
  and (_00582_, _00581_, _35815_);
  not (_00583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor (_00584_, _00581_, _00583_);
  or (_38616_, _00584_, _00582_);
  and (_00585_, _00581_, _35822_);
  not (_00586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor (_00587_, _00581_, _00586_);
  or (_38617_, _00587_, _00585_);
  and (_00588_, _00581_, _35826_);
  not (_00589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  nor (_00590_, _00581_, _00589_);
  or (_38618_, _00590_, _00588_);
  and (_00591_, _00581_, _35830_);
  not (_00592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor (_00593_, _00581_, _00592_);
  or (_38619_, _00593_, _00591_);
  and (_00594_, _00581_, _35834_);
  not (_00595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  nor (_00596_, _00581_, _00595_);
  or (_38620_, _00596_, _00594_);
  and (_00597_, _00581_, _35838_);
  not (_00598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  nor (_00599_, _00581_, _00598_);
  or (_38621_, _00599_, _00597_);
  and (_00600_, _00581_, _35842_);
  not (_00601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  nor (_00602_, _00581_, _00601_);
  or (_38622_, _00602_, _00600_);
  and (_00603_, _00581_, _35846_);
  not (_00604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  nor (_00605_, _00581_, _00604_);
  or (_38623_, _00605_, _00603_);
  and (_00606_, _00305_, _36115_);
  and (_00607_, _00606_, _35815_);
  not (_00608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  nor (_00609_, _00606_, _00608_);
  or (_38632_, _00609_, _00607_);
  and (_00610_, _00606_, _35822_);
  not (_00611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  nor (_00612_, _00606_, _00611_);
  or (_38633_, _00612_, _00610_);
  and (_00613_, _00606_, _35826_);
  not (_00614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor (_00615_, _00606_, _00614_);
  or (_38634_, _00615_, _00613_);
  and (_00616_, _00606_, _35830_);
  not (_00617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  nor (_00618_, _00606_, _00617_);
  or (_38635_, _00618_, _00616_);
  and (_00619_, _00606_, _35834_);
  not (_00620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor (_00621_, _00606_, _00620_);
  or (_38636_, _00621_, _00619_);
  and (_00622_, _00606_, _35838_);
  not (_00623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  nor (_00624_, _00606_, _00623_);
  or (_38637_, _00624_, _00622_);
  and (_00625_, _00606_, _35842_);
  not (_00626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor (_00627_, _00606_, _00626_);
  or (_38638_, _00627_, _00625_);
  and (_00628_, _00606_, _35846_);
  not (_00629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  nor (_00630_, _00606_, _00629_);
  or (_38639_, _00630_, _00628_);
  and (_00631_, _00305_, _36141_);
  and (_00632_, _00631_, _35815_);
  not (_00633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  nor (_00634_, _00631_, _00633_);
  or (_38640_, _00634_, _00632_);
  and (_00635_, _00631_, _35822_);
  not (_00636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor (_00637_, _00631_, _00636_);
  or (_38641_, _00637_, _00635_);
  and (_00638_, _00631_, _35826_);
  not (_00639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor (_00640_, _00631_, _00639_);
  or (_38642_, _00640_, _00638_);
  and (_00641_, _00631_, _35830_);
  not (_00642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor (_00643_, _00631_, _00642_);
  or (_38643_, _00643_, _00641_);
  and (_00644_, _00631_, _35834_);
  not (_00645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nor (_00646_, _00631_, _00645_);
  or (_38644_, _00646_, _00644_);
  and (_00647_, _00631_, _35838_);
  not (_00648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor (_00649_, _00631_, _00648_);
  or (_38645_, _00649_, _00647_);
  and (_00650_, _00631_, _35842_);
  not (_00651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor (_00652_, _00631_, _00651_);
  or (_38646_, _00652_, _00650_);
  and (_00653_, _00631_, _35846_);
  not (_00654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  nor (_00655_, _00631_, _00654_);
  or (_38647_, _00655_, _00653_);
  and (_00656_, _00305_, _36167_);
  and (_00657_, _00656_, _35815_);
  not (_00658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor (_00659_, _00656_, _00658_);
  or (_38648_, _00659_, _00657_);
  and (_00660_, _00656_, _35822_);
  not (_00661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  nor (_00662_, _00656_, _00661_);
  or (_38649_, _00662_, _00660_);
  and (_00663_, _00656_, _35826_);
  not (_00664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  nor (_00665_, _00656_, _00664_);
  or (_38650_, _00665_, _00663_);
  and (_00666_, _00656_, _35830_);
  not (_00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  nor (_00668_, _00656_, _00667_);
  or (_38651_, _00668_, _00666_);
  and (_00669_, _00656_, _35834_);
  not (_00670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  nor (_00671_, _00656_, _00670_);
  or (_38652_, _00671_, _00669_);
  and (_00672_, _00656_, _35838_);
  not (_00673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  nor (_00674_, _00656_, _00673_);
  or (_38653_, _00674_, _00672_);
  and (_00675_, _00656_, _35842_);
  not (_00676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  nor (_00677_, _00656_, _00676_);
  or (_38654_, _00677_, _00675_);
  and (_00678_, _00656_, _35846_);
  not (_00679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor (_00680_, _00656_, _00679_);
  or (_38655_, _00680_, _00678_);
  and (_00681_, _00305_, _36193_);
  and (_00682_, _00681_, _35815_);
  not (_00683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor (_00684_, _00681_, _00683_);
  or (_38656_, _00684_, _00682_);
  and (_00685_, _00681_, _35822_);
  not (_00686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  nor (_00687_, _00681_, _00686_);
  or (_38657_, _00687_, _00685_);
  and (_00688_, _00681_, _35826_);
  not (_00689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor (_00690_, _00681_, _00689_);
  or (_38658_, _00690_, _00688_);
  and (_00691_, _00681_, _35830_);
  not (_00692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  nor (_00693_, _00681_, _00692_);
  or (_38659_, _00693_, _00691_);
  and (_00694_, _00681_, _35834_);
  not (_00695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  nor (_00696_, _00681_, _00695_);
  or (_38660_, _00696_, _00694_);
  and (_00697_, _00681_, _35838_);
  not (_00698_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  nor (_00699_, _00681_, _00698_);
  or (_38661_, _00699_, _00697_);
  and (_00700_, _00681_, _35842_);
  not (_00701_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor (_00702_, _00681_, _00701_);
  or (_38662_, _00702_, _00700_);
  and (_00703_, _00681_, _35846_);
  not (_00704_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  nor (_00705_, _00681_, _00704_);
  or (_38663_, _00705_, _00703_);
  and (_00706_, _33659_, _33618_);
  and (_00707_, _00706_, _34693_);
  and (_00708_, _00707_, _35575_);
  and (_00709_, _00708_, _35572_);
  and (_00710_, _00709_, _35815_);
  not (_00711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  nor (_00712_, _00709_, _00711_);
  or (_38664_, _00712_, _00710_);
  and (_00713_, _00709_, _35822_);
  not (_00714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nor (_00715_, _00709_, _00714_);
  or (_38665_, _00715_, _00713_);
  and (_00716_, _00709_, _35826_);
  not (_00717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  nor (_00718_, _00709_, _00717_);
  or (_38666_, _00718_, _00716_);
  and (_00719_, _00709_, _35830_);
  not (_00720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  nor (_00721_, _00709_, _00720_);
  or (_38667_, _00721_, _00719_);
  and (_00722_, _00709_, _35834_);
  not (_00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nor (_00724_, _00709_, _00723_);
  or (_38668_, _00724_, _00722_);
  and (_00725_, _00709_, _35838_);
  not (_00726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nor (_00727_, _00709_, _00726_);
  or (_38669_, _00727_, _00725_);
  and (_00728_, _00709_, _35842_);
  not (_00729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  nor (_00730_, _00709_, _00729_);
  or (_38670_, _00730_, _00728_);
  and (_00731_, _00709_, _35846_);
  not (_00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  nor (_00733_, _00709_, _00732_);
  or (_38671_, _00733_, _00731_);
  and (_00734_, _00708_, _35817_);
  and (_00735_, _00734_, _35815_);
  not (_00736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nor (_00737_, _00734_, _00736_);
  or (_38672_, _00737_, _00735_);
  and (_00738_, _00734_, _35822_);
  not (_00739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  nor (_00740_, _00734_, _00739_);
  or (_38673_, _00740_, _00738_);
  and (_00741_, _00734_, _35826_);
  not (_00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nor (_00743_, _00734_, _00742_);
  or (_38674_, _00743_, _00741_);
  and (_00744_, _00734_, _35830_);
  not (_00745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nor (_00746_, _00734_, _00745_);
  or (_38675_, _00746_, _00744_);
  and (_00747_, _00734_, _35834_);
  not (_00748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  nor (_00749_, _00734_, _00748_);
  or (_38676_, _00749_, _00747_);
  and (_00750_, _00734_, _35838_);
  not (_00751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  nor (_00752_, _00734_, _00751_);
  or (_38677_, _00752_, _00750_);
  and (_00753_, _00734_, _35842_);
  not (_00754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nor (_00755_, _00734_, _00754_);
  or (_38678_, _00755_, _00753_);
  and (_00756_, _00734_, _35846_);
  not (_00757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  nor (_00758_, _00734_, _00757_);
  or (_38679_, _00758_, _00756_);
  and (_00759_, _00708_, _35851_);
  and (_00760_, _00759_, _35815_);
  not (_00761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  nor (_00762_, _00759_, _00761_);
  or (_38680_, _00762_, _00760_);
  and (_00763_, _00759_, _35822_);
  not (_00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nor (_00765_, _00759_, _00764_);
  or (_38681_, _00765_, _00763_);
  and (_00766_, _00759_, _35826_);
  not (_00767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  nor (_00768_, _00759_, _00767_);
  or (_38682_, _00768_, _00766_);
  and (_00769_, _00759_, _35830_);
  not (_00770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  nor (_00771_, _00759_, _00770_);
  or (_38683_, _00771_, _00769_);
  and (_00772_, _00759_, _35834_);
  not (_00773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nor (_00774_, _00759_, _00773_);
  or (_38684_, _00774_, _00772_);
  and (_00775_, _00759_, _35838_);
  not (_00776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  nor (_00777_, _00759_, _00776_);
  or (_38685_, _00777_, _00775_);
  and (_00778_, _00759_, _35842_);
  not (_00779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  nor (_00780_, _00759_, _00779_);
  or (_38686_, _00780_, _00778_);
  and (_00781_, _00759_, _35846_);
  not (_00782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  nor (_00783_, _00759_, _00782_);
  or (_38687_, _00783_, _00781_);
  and (_00784_, _00708_, _35878_);
  and (_00785_, _00784_, _35815_);
  not (_00786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nor (_00787_, _00784_, _00786_);
  or (_38688_, _00787_, _00785_);
  and (_00788_, _00784_, _35822_);
  not (_00789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  nor (_00790_, _00784_, _00789_);
  or (_38689_, _00790_, _00788_);
  and (_00791_, _00784_, _35826_);
  not (_00792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nor (_00793_, _00784_, _00792_);
  or (_38690_, _00793_, _00791_);
  and (_00794_, _00784_, _35830_);
  not (_00795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nor (_00796_, _00784_, _00795_);
  or (_38691_, _00796_, _00794_);
  and (_00797_, _00784_, _35834_);
  not (_00798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  nor (_00799_, _00784_, _00798_);
  or (_38692_, _00799_, _00797_);
  and (_00800_, _00784_, _35838_);
  not (_00801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  nor (_00802_, _00784_, _00801_);
  or (_38693_, _00802_, _00800_);
  and (_00803_, _00784_, _35842_);
  not (_00804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nor (_00805_, _00784_, _00804_);
  or (_38694_, _00805_, _00803_);
  and (_00806_, _00784_, _35846_);
  not (_00807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  nor (_00808_, _00784_, _00807_);
  or (_38695_, _00808_, _00806_);
  and (_00809_, _00708_, _35905_);
  and (_00810_, _00809_, _35815_);
  not (_00811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  nor (_00812_, _00809_, _00811_);
  or (_38696_, _00812_, _00810_);
  and (_00813_, _00809_, _35822_);
  not (_00814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nor (_00815_, _00809_, _00814_);
  or (_38697_, _00815_, _00813_);
  and (_00816_, _00809_, _35826_);
  not (_00817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  nor (_00818_, _00809_, _00817_);
  or (_38698_, _00818_, _00816_);
  and (_00819_, _00809_, _35830_);
  not (_00820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  nor (_00821_, _00809_, _00820_);
  or (_38699_, _00821_, _00819_);
  and (_00822_, _00809_, _35834_);
  not (_00823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nor (_00824_, _00809_, _00823_);
  or (_38700_, _00824_, _00822_);
  and (_00825_, _00809_, _35838_);
  not (_00826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  nor (_00827_, _00809_, _00826_);
  or (_38701_, _00827_, _00825_);
  and (_00828_, _00809_, _35842_);
  not (_00829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  nor (_00830_, _00809_, _00829_);
  or (_38702_, _00830_, _00828_);
  and (_00831_, _00809_, _35846_);
  not (_00832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  nor (_00833_, _00809_, _00832_);
  or (_38703_, _00833_, _00831_);
  and (_00834_, _00708_, _35931_);
  and (_00835_, _00834_, _35815_);
  not (_00836_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  nor (_00837_, _00834_, _00836_);
  or (_38704_, _00837_, _00835_);
  and (_00838_, _00834_, _35822_);
  not (_00839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  nor (_00840_, _00834_, _00839_);
  or (_38705_, _00840_, _00838_);
  and (_00841_, _00834_, _35826_);
  not (_00842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  nor (_00843_, _00834_, _00842_);
  or (_38706_, _00843_, _00841_);
  and (_00844_, _00834_, _35830_);
  not (_00845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nor (_00846_, _00834_, _00845_);
  or (_38707_, _00846_, _00844_);
  and (_00847_, _00834_, _35834_);
  not (_00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nor (_00849_, _00834_, _00848_);
  or (_38708_, _00849_, _00847_);
  and (_00850_, _00834_, _35838_);
  not (_00851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  nor (_00852_, _00834_, _00851_);
  or (_38709_, _00852_, _00850_);
  and (_00853_, _00834_, _35842_);
  not (_00854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  nor (_00855_, _00834_, _00854_);
  or (_38710_, _00855_, _00853_);
  and (_00856_, _00834_, _35846_);
  not (_00857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  nor (_00858_, _00834_, _00857_);
  or (_38711_, _00858_, _00856_);
  and (_00859_, _00708_, _35957_);
  and (_00860_, _00859_, _35815_);
  not (_00861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nor (_00862_, _00859_, _00861_);
  or (_38720_, _00862_, _00860_);
  and (_00863_, _00859_, _35822_);
  not (_00864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nor (_00865_, _00859_, _00864_);
  or (_38721_, _00865_, _00863_);
  and (_00866_, _00859_, _35826_);
  not (_00867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nor (_00868_, _00859_, _00867_);
  or (_38722_, _00868_, _00866_);
  and (_00869_, _00859_, _35830_);
  not (_00870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  nor (_00871_, _00859_, _00870_);
  or (_38723_, _00871_, _00869_);
  and (_00872_, _00859_, _35834_);
  not (_00873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  nor (_00874_, _00859_, _00873_);
  or (_38724_, _00874_, _00872_);
  and (_00875_, _00859_, _35838_);
  not (_00876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  nor (_00877_, _00859_, _00876_);
  or (_38725_, _00877_, _00875_);
  and (_00878_, _00859_, _35842_);
  not (_00879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nor (_00880_, _00859_, _00879_);
  or (_38726_, _00880_, _00878_);
  and (_00881_, _00859_, _35846_);
  not (_00882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  nor (_00883_, _00859_, _00882_);
  or (_38727_, _00883_, _00881_);
  and (_00884_, _00708_, _35983_);
  and (_00885_, _00884_, _35815_);
  not (_00886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  nor (_00887_, _00884_, _00886_);
  or (_38728_, _00887_, _00885_);
  and (_00888_, _00884_, _35822_);
  not (_00889_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  nor (_00890_, _00884_, _00889_);
  or (_38729_, _00890_, _00888_);
  and (_00891_, _00884_, _35826_);
  not (_00892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nor (_00893_, _00884_, _00892_);
  or (_38730_, _00893_, _00891_);
  and (_00894_, _00884_, _35830_);
  not (_00895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  nor (_00896_, _00884_, _00895_);
  or (_38731_, _00896_, _00894_);
  and (_00897_, _00884_, _35834_);
  not (_00898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  nor (_00899_, _00884_, _00898_);
  or (_38732_, _00899_, _00897_);
  and (_00900_, _00884_, _35838_);
  not (_00901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  nor (_00902_, _00884_, _00901_);
  or (_38733_, _00902_, _00900_);
  and (_00903_, _00884_, _35842_);
  not (_00904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  nor (_00905_, _00884_, _00904_);
  or (_38734_, _00905_, _00903_);
  and (_00906_, _00884_, _35846_);
  not (_00907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  nor (_00908_, _00884_, _00907_);
  or (_38735_, _00908_, _00906_);
  and (_00909_, _00708_, _36010_);
  and (_00910_, _00909_, _35815_);
  not (_00911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nor (_00912_, _00909_, _00911_);
  or (_38736_, _00912_, _00910_);
  and (_00913_, _00909_, _35822_);
  not (_00914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor (_00915_, _00909_, _00914_);
  or (_38737_, _00915_, _00913_);
  and (_00916_, _00909_, _35826_);
  not (_00917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  nor (_00918_, _00909_, _00917_);
  or (_38738_, _00918_, _00916_);
  and (_00919_, _00909_, _35830_);
  not (_00920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nor (_00921_, _00909_, _00920_);
  or (_38739_, _00921_, _00919_);
  and (_00922_, _00909_, _35834_);
  not (_00923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nor (_00924_, _00909_, _00923_);
  or (_38740_, _00924_, _00922_);
  and (_00925_, _00909_, _35838_);
  not (_00926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  nor (_00927_, _00909_, _00926_);
  or (_38741_, _00927_, _00925_);
  and (_00928_, _00909_, _35842_);
  not (_00929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nor (_00930_, _00909_, _00929_);
  or (_38742_, _00930_, _00928_);
  and (_00931_, _00909_, _35846_);
  not (_00932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  nor (_00933_, _00909_, _00932_);
  or (_38743_, _00933_, _00931_);
  and (_00934_, _00708_, _36036_);
  and (_00935_, _00934_, _35815_);
  not (_00936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  nor (_00937_, _00934_, _00936_);
  or (_38744_, _00937_, _00935_);
  and (_00938_, _00934_, _35822_);
  not (_00939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  nor (_00940_, _00934_, _00939_);
  or (_38745_, _00940_, _00938_);
  and (_00941_, _00934_, _35826_);
  not (_00942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  nor (_00943_, _00934_, _00942_);
  or (_38746_, _00943_, _00941_);
  and (_00944_, _00934_, _35830_);
  not (_00945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nor (_00946_, _00934_, _00945_);
  or (_38747_, _00946_, _00944_);
  and (_00947_, _00934_, _35834_);
  not (_00948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  nor (_00949_, _00934_, _00948_);
  or (_38748_, _00949_, _00947_);
  and (_00950_, _00934_, _35838_);
  not (_00951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  nor (_00952_, _00934_, _00951_);
  or (_38749_, _00952_, _00950_);
  and (_00953_, _00934_, _35842_);
  not (_00954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  nor (_00955_, _00934_, _00954_);
  or (_38750_, _00955_, _00953_);
  and (_00956_, _00934_, _35846_);
  not (_00957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  nor (_00958_, _00934_, _00957_);
  or (_38751_, _00958_, _00956_);
  and (_00959_, _00708_, _36062_);
  and (_00960_, _00959_, _35815_);
  not (_00961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor (_00962_, _00959_, _00961_);
  or (_38752_, _00962_, _00960_);
  and (_00963_, _00959_, _35822_);
  not (_00964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor (_00965_, _00959_, _00964_);
  or (_38753_, _00965_, _00963_);
  and (_00966_, _00959_, _35826_);
  not (_00967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor (_00968_, _00959_, _00967_);
  or (_38754_, _00968_, _00966_);
  and (_00969_, _00959_, _35830_);
  not (_00970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  nor (_00971_, _00959_, _00970_);
  or (_38755_, _00971_, _00969_);
  and (_00972_, _00959_, _35834_);
  not (_00973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nor (_00974_, _00959_, _00973_);
  or (_38756_, _00974_, _00972_);
  and (_00975_, _00959_, _35838_);
  not (_00976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  nor (_00977_, _00959_, _00976_);
  or (_38757_, _00977_, _00975_);
  and (_00978_, _00959_, _35842_);
  not (_00979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor (_00980_, _00959_, _00979_);
  or (_38758_, _00980_, _00978_);
  and (_00981_, _00959_, _35846_);
  not (_00982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  nor (_00983_, _00959_, _00982_);
  or (_38759_, _00983_, _00981_);
  and (_00984_, _00708_, _36088_);
  and (_00985_, _00984_, _35815_);
  not (_00986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nor (_00987_, _00984_, _00986_);
  or (_38760_, _00987_, _00985_);
  and (_00988_, _00984_, _35822_);
  not (_00989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor (_00990_, _00984_, _00989_);
  or (_38761_, _00990_, _00988_);
  and (_00991_, _00984_, _35826_);
  not (_00992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor (_00993_, _00984_, _00992_);
  or (_38762_, _00993_, _00991_);
  and (_00994_, _00984_, _35830_);
  not (_00995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  nor (_00996_, _00984_, _00995_);
  or (_38763_, _00996_, _00994_);
  and (_00997_, _00984_, _35834_);
  not (_00998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  nor (_00999_, _00984_, _00998_);
  or (_38764_, _00999_, _00997_);
  and (_01000_, _00984_, _35838_);
  not (_01001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  nor (_01002_, _00984_, _01001_);
  or (_38765_, _01002_, _01000_);
  and (_01003_, _00984_, _35842_);
  not (_01004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor (_01005_, _00984_, _01004_);
  or (_38766_, _01005_, _01003_);
  and (_01006_, _00984_, _35846_);
  not (_01007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  nor (_01008_, _00984_, _01007_);
  or (_38767_, _01008_, _01006_);
  and (_01009_, _00708_, _36115_);
  and (_01010_, _01009_, _35815_);
  not (_01011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  nor (_01012_, _01009_, _01011_);
  or (_38768_, _01012_, _01010_);
  and (_01013_, _01009_, _35822_);
  not (_01014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  nor (_01015_, _01009_, _01014_);
  or (_38769_, _01015_, _01013_);
  and (_01016_, _01009_, _35826_);
  not (_01017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  nor (_01018_, _01009_, _01017_);
  or (_38770_, _01018_, _01016_);
  and (_01019_, _01009_, _35830_);
  not (_01020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nor (_01021_, _01009_, _01020_);
  or (_38771_, _01021_, _01019_);
  and (_01022_, _01009_, _35834_);
  not (_01023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nor (_01024_, _01009_, _01023_);
  or (_38772_, _01024_, _01022_);
  and (_01025_, _01009_, _35838_);
  not (_01026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  nor (_01027_, _01009_, _01026_);
  or (_38773_, _01027_, _01025_);
  and (_01028_, _01009_, _35842_);
  not (_01029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  nor (_01030_, _01009_, _01029_);
  or (_38774_, _01030_, _01028_);
  and (_01031_, _01009_, _35846_);
  not (_01032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  nor (_01033_, _01009_, _01032_);
  or (_38775_, _01033_, _01031_);
  and (_01034_, _00708_, _36141_);
  and (_01035_, _01034_, _35815_);
  not (_01036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nor (_01037_, _01034_, _01036_);
  or (_38776_, _01037_, _01035_);
  and (_01038_, _01034_, _35822_);
  not (_01039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nor (_01040_, _01034_, _01039_);
  or (_38777_, _01040_, _01038_);
  and (_01041_, _01034_, _35826_);
  not (_01042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  nor (_01043_, _01034_, _01042_);
  or (_38778_, _01043_, _01041_);
  and (_01044_, _01034_, _35830_);
  not (_01045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nor (_01046_, _01034_, _01045_);
  or (_38779_, _01046_, _01044_);
  and (_01047_, _01034_, _35834_);
  not (_01048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  nor (_01049_, _01034_, _01048_);
  or (_38780_, _01049_, _01047_);
  and (_01050_, _01034_, _35838_);
  not (_01051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  nor (_01052_, _01034_, _01051_);
  or (_38781_, _01052_, _01050_);
  and (_01053_, _01034_, _35842_);
  not (_01054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nor (_01055_, _01034_, _01054_);
  or (_38782_, _01055_, _01053_);
  and (_01056_, _01034_, _35846_);
  not (_01057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  nor (_01058_, _01034_, _01057_);
  or (_38783_, _01058_, _01056_);
  and (_01059_, _00708_, _36167_);
  and (_01060_, _01059_, _35815_);
  not (_01061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  nor (_01062_, _01059_, _01061_);
  or (_38784_, _01062_, _01060_);
  and (_01063_, _01059_, _35822_);
  not (_01064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  nor (_01065_, _01059_, _01064_);
  or (_38785_, _01065_, _01063_);
  and (_01066_, _01059_, _35826_);
  not (_01067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nor (_01068_, _01059_, _01067_);
  or (_38786_, _01068_, _01066_);
  and (_01069_, _01059_, _35830_);
  not (_01070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  nor (_01071_, _01059_, _01070_);
  or (_38787_, _01071_, _01069_);
  and (_01072_, _01059_, _35834_);
  not (_01073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor (_01074_, _01059_, _01073_);
  or (_38788_, _01074_, _01072_);
  and (_01075_, _01059_, _35838_);
  not (_01076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  nor (_01077_, _01059_, _01076_);
  or (_38789_, _01077_, _01075_);
  and (_01078_, _01059_, _35842_);
  not (_01079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  nor (_01080_, _01059_, _01079_);
  or (_38790_, _01080_, _01078_);
  and (_01081_, _01059_, _35846_);
  not (_01082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  nor (_01083_, _01059_, _01082_);
  or (_38791_, _01083_, _01081_);
  and (_01084_, _00708_, _36193_);
  and (_01085_, _01084_, _35815_);
  not (_01086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  nor (_01087_, _01084_, _01086_);
  or (_38792_, _01087_, _01085_);
  and (_01088_, _01084_, _35822_);
  not (_01089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor (_01090_, _01084_, _01089_);
  or (_38793_, _01090_, _01088_);
  and (_01091_, _01084_, _35826_);
  not (_01092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  nor (_01093_, _01084_, _01092_);
  or (_38794_, _01093_, _01091_);
  and (_01094_, _01084_, _35830_);
  not (_01095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor (_01096_, _01084_, _01095_);
  or (_38795_, _01096_, _01094_);
  and (_01097_, _01084_, _35834_);
  not (_01098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  nor (_01099_, _01084_, _01098_);
  or (_38796_, _01099_, _01097_);
  and (_01100_, _01084_, _35838_);
  not (_01101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  nor (_01102_, _01084_, _01101_);
  or (_38797_, _01102_, _01100_);
  and (_01103_, _01084_, _35842_);
  not (_01104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor (_01105_, _01084_, _01104_);
  or (_38798_, _01105_, _01103_);
  and (_01106_, _01084_, _35846_);
  not (_01107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  nor (_01108_, _01084_, _01107_);
  or (_38799_, _01108_, _01106_);
  and (_01109_, _00707_, _36220_);
  and (_01110_, _01109_, _35572_);
  and (_01111_, _01110_, _35815_);
  not (_01112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nor (_01113_, _01110_, _01112_);
  or (_38808_, _01113_, _01111_);
  and (_01114_, _01110_, _35822_);
  not (_01115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  nor (_01116_, _01110_, _01115_);
  or (_38809_, _01116_, _01114_);
  and (_01117_, _01110_, _35826_);
  not (_01118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nor (_01119_, _01110_, _01118_);
  or (_38810_, _01119_, _01117_);
  and (_01120_, _01110_, _35830_);
  not (_01121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  nor (_01122_, _01110_, _01121_);
  or (_38811_, _01122_, _01120_);
  and (_01123_, _01110_, _35834_);
  not (_01124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nor (_01125_, _01110_, _01124_);
  or (_38812_, _01125_, _01123_);
  and (_01126_, _01110_, _35838_);
  not (_01127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  nor (_01128_, _01110_, _01127_);
  or (_38813_, _01128_, _01126_);
  and (_01129_, _01110_, _35842_);
  not (_01130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  nor (_01131_, _01110_, _01130_);
  or (_38814_, _01131_, _01129_);
  and (_01132_, _01110_, _35846_);
  not (_01133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  nor (_01134_, _01110_, _01133_);
  or (_38815_, _01134_, _01132_);
  and (_01135_, _01109_, _35817_);
  and (_01136_, _01135_, _35815_);
  not (_01137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nor (_01138_, _01135_, _01137_);
  or (_38816_, _01138_, _01136_);
  and (_01139_, _01135_, _35822_);
  not (_01140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  nor (_01141_, _01135_, _01140_);
  or (_38817_, _01141_, _01139_);
  and (_01142_, _01135_, _35826_);
  not (_01143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nor (_01144_, _01135_, _01143_);
  or (_38818_, _01144_, _01142_);
  and (_01145_, _01135_, _35830_);
  not (_01146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nor (_01147_, _01135_, _01146_);
  or (_38819_, _01147_, _01145_);
  and (_01148_, _01135_, _35834_);
  not (_01149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  nor (_01150_, _01135_, _01149_);
  or (_38820_, _01150_, _01148_);
  and (_01151_, _01135_, _35838_);
  not (_01152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nor (_01153_, _01135_, _01152_);
  or (_38821_, _01153_, _01151_);
  and (_01154_, _01135_, _35842_);
  not (_01155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  nor (_01156_, _01135_, _01155_);
  or (_38822_, _01156_, _01154_);
  and (_01157_, _01135_, _35846_);
  not (_01158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  nor (_01159_, _01135_, _01158_);
  or (_38823_, _01159_, _01157_);
  and (_01160_, _01109_, _35851_);
  and (_01161_, _01160_, _35815_);
  not (_01162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  nor (_01163_, _01160_, _01162_);
  or (_38824_, _01163_, _01161_);
  and (_01164_, _01160_, _35822_);
  not (_01165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nor (_01166_, _01160_, _01165_);
  or (_38825_, _01166_, _01164_);
  and (_01167_, _01160_, _35826_);
  not (_01168_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  nor (_01169_, _01160_, _01168_);
  or (_38826_, _01169_, _01167_);
  and (_01170_, _01160_, _35830_);
  not (_01171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  nor (_01172_, _01160_, _01171_);
  or (_38827_, _01172_, _01170_);
  and (_01173_, _01160_, _35834_);
  not (_01174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nor (_01175_, _01160_, _01174_);
  or (_38828_, _01175_, _01173_);
  and (_01176_, _01160_, _35838_);
  not (_01177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  nor (_01178_, _01160_, _01177_);
  or (_38829_, _01178_, _01176_);
  and (_01179_, _01160_, _35842_);
  not (_01180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nor (_01181_, _01160_, _01180_);
  or (_38830_, _01181_, _01179_);
  and (_01182_, _01160_, _35846_);
  not (_01183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nor (_01184_, _01160_, _01183_);
  or (_38831_, _01184_, _01182_);
  and (_01185_, _01109_, _35878_);
  and (_01186_, _01185_, _35815_);
  not (_01187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nor (_01188_, _01185_, _01187_);
  or (_38832_, _01188_, _01186_);
  and (_01189_, _01185_, _35822_);
  not (_01190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nor (_01191_, _01185_, _01190_);
  or (_38833_, _01191_, _01189_);
  and (_01192_, _01185_, _35826_);
  not (_01193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nor (_01194_, _01185_, _01193_);
  or (_38834_, _01194_, _01192_);
  and (_01195_, _01185_, _35830_);
  not (_01196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  nor (_01197_, _01185_, _01196_);
  or (_38835_, _01197_, _01195_);
  and (_01198_, _01185_, _35834_);
  not (_01199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nor (_01200_, _01185_, _01199_);
  or (_38836_, _01200_, _01198_);
  and (_01201_, _01185_, _35838_);
  not (_01202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  nor (_01203_, _01185_, _01202_);
  or (_38837_, _01203_, _01201_);
  and (_01204_, _01185_, _35842_);
  not (_01205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nor (_01206_, _01185_, _01205_);
  or (_38838_, _01206_, _01204_);
  and (_01207_, _01185_, _35846_);
  not (_01208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  nor (_01209_, _01185_, _01208_);
  or (_38839_, _01209_, _01207_);
  and (_01210_, _01109_, _35905_);
  and (_01211_, _01210_, _35815_);
  not (_01212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  nor (_01213_, _01210_, _01212_);
  or (_38840_, _01213_, _01211_);
  and (_01214_, _01210_, _35822_);
  not (_01215_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  nor (_01216_, _01210_, _01215_);
  or (_38841_, _01216_, _01214_);
  and (_01217_, _01210_, _35826_);
  not (_01218_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  nor (_01219_, _01210_, _01218_);
  or (_38842_, _01219_, _01217_);
  and (_01220_, _01210_, _35830_);
  not (_01221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nor (_01222_, _01210_, _01221_);
  or (_38843_, _01222_, _01220_);
  and (_01223_, _01210_, _35834_);
  not (_01224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  nor (_01225_, _01210_, _01224_);
  or (_38844_, _01225_, _01223_);
  and (_01226_, _01210_, _35838_);
  not (_01227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  nor (_01228_, _01210_, _01227_);
  or (_38845_, _01228_, _01226_);
  and (_01229_, _01210_, _35842_);
  not (_01230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  nor (_01231_, _01210_, _01230_);
  or (_38846_, _01231_, _01229_);
  and (_01232_, _01210_, _35846_);
  not (_01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  nor (_01234_, _01210_, _01233_);
  or (_38847_, _01234_, _01232_);
  and (_01235_, _01109_, _35931_);
  and (_01236_, _01235_, _35815_);
  not (_01237_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nor (_01238_, _01235_, _01237_);
  or (_38848_, _01238_, _01236_);
  and (_01239_, _01235_, _35822_);
  not (_01240_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  nor (_01241_, _01235_, _01240_);
  or (_38849_, _01241_, _01239_);
  and (_01242_, _01235_, _35826_);
  not (_01243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nor (_01244_, _01235_, _01243_);
  or (_38850_, _01244_, _01242_);
  and (_01245_, _01235_, _35830_);
  not (_01246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  nor (_01247_, _01235_, _01246_);
  or (_38851_, _01247_, _01245_);
  and (_01248_, _01235_, _35834_);
  not (_01249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  nor (_01250_, _01235_, _01249_);
  or (_38852_, _01250_, _01248_);
  and (_01251_, _01235_, _35838_);
  not (_01252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  nor (_01253_, _01235_, _01252_);
  or (_38853_, _01253_, _01251_);
  and (_01254_, _01235_, _35842_);
  not (_01255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nor (_01256_, _01235_, _01255_);
  or (_38854_, _01256_, _01254_);
  and (_01257_, _01235_, _35846_);
  not (_01258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  nor (_01259_, _01235_, _01258_);
  or (_38855_, _01259_, _01257_);
  and (_01260_, _01109_, _35957_);
  and (_01261_, _01260_, _35815_);
  not (_01262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  nor (_01263_, _01260_, _01262_);
  or (_38856_, _01263_, _01261_);
  and (_01264_, _01260_, _35822_);
  not (_01265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nor (_01266_, _01260_, _01265_);
  or (_38857_, _01266_, _01264_);
  and (_01267_, _01260_, _35826_);
  not (_01268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  nor (_01269_, _01260_, _01268_);
  or (_38858_, _01269_, _01267_);
  and (_01270_, _01260_, _35830_);
  not (_01271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nor (_01272_, _01260_, _01271_);
  or (_38859_, _01272_, _01270_);
  and (_01273_, _01260_, _35834_);
  not (_01274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nor (_01275_, _01260_, _01274_);
  or (_38860_, _01275_, _01273_);
  and (_01276_, _01260_, _35838_);
  not (_01277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  nor (_01278_, _01260_, _01277_);
  or (_38861_, _01278_, _01276_);
  and (_01279_, _01260_, _35842_);
  not (_01280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  nor (_01281_, _01260_, _01280_);
  or (_38862_, _01281_, _01279_);
  and (_01282_, _01260_, _35846_);
  not (_01283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  nor (_01284_, _01260_, _01283_);
  or (_38863_, _01284_, _01282_);
  and (_01285_, _01109_, _35983_);
  and (_01286_, _01285_, _35815_);
  not (_01287_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nor (_01288_, _01285_, _01287_);
  or (_38864_, _01288_, _01286_);
  and (_01289_, _01285_, _35822_);
  not (_01290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nor (_01291_, _01285_, _01290_);
  or (_38865_, _01291_, _01289_);
  and (_01292_, _01285_, _35826_);
  not (_01293_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  nor (_01294_, _01285_, _01293_);
  or (_38866_, _01294_, _01292_);
  and (_01295_, _01285_, _35830_);
  not (_01296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  nor (_01297_, _01285_, _01296_);
  or (_38867_, _01297_, _01295_);
  and (_01298_, _01285_, _35834_);
  not (_01299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  nor (_01300_, _01285_, _01299_);
  or (_38868_, _01300_, _01298_);
  and (_01301_, _01285_, _35838_);
  not (_01302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  nor (_01303_, _01285_, _01302_);
  or (_38869_, _01303_, _01301_);
  and (_01304_, _01285_, _35842_);
  not (_01305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nor (_01306_, _01285_, _01305_);
  or (_38870_, _01306_, _01304_);
  and (_01307_, _01285_, _35846_);
  not (_01308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  nor (_01309_, _01285_, _01308_);
  or (_38871_, _01309_, _01307_);
  and (_01310_, _01109_, _36010_);
  and (_01311_, _01310_, _35815_);
  not (_01312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  nor (_01313_, _01310_, _01312_);
  or (_38872_, _01313_, _01311_);
  and (_01314_, _01310_, _35822_);
  not (_01315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  nor (_01316_, _01310_, _01315_);
  or (_38873_, _01316_, _01314_);
  and (_01317_, _01310_, _35826_);
  not (_01318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor (_01319_, _01310_, _01318_);
  or (_38874_, _01319_, _01317_);
  and (_01320_, _01310_, _35830_);
  not (_01321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor (_01322_, _01310_, _01321_);
  or (_38875_, _01322_, _01320_);
  and (_01323_, _01310_, _35834_);
  not (_01324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor (_01325_, _01310_, _01324_);
  or (_38876_, _01325_, _01323_);
  and (_01326_, _01310_, _35838_);
  not (_01327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  nor (_01328_, _01310_, _01327_);
  or (_38877_, _01328_, _01326_);
  and (_01329_, _01310_, _35842_);
  not (_01330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  nor (_01331_, _01310_, _01330_);
  or (_38878_, _01331_, _01329_);
  and (_01332_, _01310_, _35846_);
  not (_01333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor (_01334_, _01310_, _01333_);
  or (_38879_, _01334_, _01332_);
  and (_01335_, _01109_, _36036_);
  and (_01336_, _01335_, _35815_);
  not (_01337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  nor (_01338_, _01335_, _01337_);
  or (_38880_, _01338_, _01336_);
  and (_01339_, _01335_, _35822_);
  not (_01340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  nor (_01341_, _01335_, _01340_);
  or (_38881_, _01341_, _01339_);
  and (_01342_, _01335_, _35826_);
  not (_01343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  nor (_01344_, _01335_, _01343_);
  or (_38882_, _01344_, _01342_);
  and (_01345_, _01335_, _35830_);
  not (_01346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  nor (_01347_, _01335_, _01346_);
  or (_38883_, _01347_, _01345_);
  and (_01348_, _01335_, _35834_);
  not (_01349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  nor (_01350_, _01335_, _01349_);
  or (_38884_, _01350_, _01348_);
  and (_01351_, _01335_, _35838_);
  not (_01352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  nor (_01353_, _01335_, _01352_);
  or (_38885_, _01353_, _01351_);
  and (_01354_, _01335_, _35842_);
  not (_01355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  nor (_01356_, _01335_, _01355_);
  or (_38886_, _01356_, _01354_);
  and (_01357_, _01335_, _35846_);
  not (_01358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  nor (_01359_, _01335_, _01358_);
  or (_38887_, _01359_, _01357_);
  and (_01360_, _01109_, _36062_);
  and (_01361_, _01360_, _35815_);
  not (_01362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor (_01363_, _01360_, _01362_);
  or (_38896_, _01363_, _01361_);
  and (_01364_, _01360_, _35822_);
  not (_01365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor (_01366_, _01360_, _01365_);
  or (_38897_, _01366_, _01364_);
  and (_01367_, _01360_, _35826_);
  not (_01368_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor (_01369_, _01360_, _01368_);
  or (_38898_, _01369_, _01367_);
  and (_01370_, _01360_, _35830_);
  not (_01371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor (_01372_, _01360_, _01371_);
  or (_38899_, _01372_, _01370_);
  and (_01373_, _01360_, _35834_);
  not (_01374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor (_01375_, _01360_, _01374_);
  or (_38900_, _01375_, _01373_);
  and (_01376_, _01360_, _35838_);
  not (_01377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  nor (_01378_, _01360_, _01377_);
  or (_38901_, _01378_, _01376_);
  and (_01379_, _01360_, _35842_);
  not (_01380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor (_01381_, _01360_, _01380_);
  or (_38902_, _01381_, _01379_);
  and (_01382_, _01360_, _35846_);
  not (_01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  nor (_01384_, _01360_, _01383_);
  or (_38903_, _01384_, _01382_);
  and (_01385_, _01109_, _36088_);
  and (_01386_, _01385_, _35815_);
  not (_01387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nor (_01388_, _01385_, _01387_);
  or (_38904_, _01388_, _01386_);
  and (_01389_, _01385_, _35822_);
  not (_01390_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  nor (_01391_, _01385_, _01390_);
  or (_38905_, _01391_, _01389_);
  and (_01392_, _01385_, _35826_);
  not (_01393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  nor (_01394_, _01385_, _01393_);
  or (_38906_, _01394_, _01392_);
  and (_01395_, _01385_, _35830_);
  not (_01396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor (_01397_, _01385_, _01396_);
  or (_38907_, _01397_, _01395_);
  and (_01398_, _01385_, _35834_);
  not (_01399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor (_01400_, _01385_, _01399_);
  or (_38908_, _01400_, _01398_);
  and (_01401_, _01385_, _35838_);
  not (_01402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  nor (_01403_, _01385_, _01402_);
  or (_38909_, _01403_, _01401_);
  and (_01404_, _01385_, _35842_);
  not (_01405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  nor (_01406_, _01385_, _01405_);
  or (_38910_, _01406_, _01404_);
  and (_01407_, _01385_, _35846_);
  not (_01408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  nor (_01409_, _01385_, _01408_);
  or (_38911_, _01409_, _01407_);
  and (_01410_, _01109_, _36115_);
  and (_01411_, _01410_, _35815_);
  not (_01412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  nor (_01413_, _01410_, _01412_);
  or (_38912_, _01413_, _01411_);
  and (_01414_, _01410_, _35822_);
  not (_01415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor (_01416_, _01410_, _01415_);
  or (_38913_, _01416_, _01414_);
  and (_01417_, _01410_, _35826_);
  not (_01418_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor (_01419_, _01410_, _01418_);
  or (_38914_, _01419_, _01417_);
  and (_01420_, _01410_, _35830_);
  not (_01421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  nor (_01422_, _01410_, _01421_);
  or (_38915_, _01422_, _01420_);
  and (_01423_, _01410_, _35834_);
  not (_01424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  nor (_01425_, _01410_, _01424_);
  or (_38916_, _01425_, _01423_);
  and (_01426_, _01410_, _35838_);
  not (_01427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  nor (_01428_, _01410_, _01427_);
  or (_38917_, _01428_, _01426_);
  and (_01429_, _01410_, _35842_);
  not (_01430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor (_01431_, _01410_, _01430_);
  or (_38918_, _01431_, _01429_);
  and (_01432_, _01410_, _35846_);
  not (_01433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor (_01434_, _01410_, _01433_);
  or (_38919_, _01434_, _01432_);
  and (_01435_, _01109_, _36141_);
  and (_01436_, _01435_, _35815_);
  not (_01437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor (_01438_, _01435_, _01437_);
  or (_38920_, _01438_, _01436_);
  and (_01439_, _01435_, _35822_);
  not (_01440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  nor (_01441_, _01435_, _01440_);
  or (_38921_, _01441_, _01439_);
  and (_01442_, _01435_, _35826_);
  not (_01443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  nor (_01444_, _01435_, _01443_);
  or (_38922_, _01444_, _01442_);
  and (_01445_, _01435_, _35830_);
  not (_01446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  nor (_01447_, _01435_, _01446_);
  or (_38923_, _01447_, _01445_);
  and (_01448_, _01435_, _35834_);
  not (_01449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor (_01450_, _01435_, _01449_);
  or (_38924_, _01450_, _01448_);
  and (_01451_, _01435_, _35838_);
  not (_01452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  nor (_01453_, _01435_, _01452_);
  or (_38925_, _01453_, _01451_);
  and (_01454_, _01435_, _35842_);
  not (_01455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  nor (_01456_, _01435_, _01455_);
  or (_38926_, _01456_, _01454_);
  and (_01457_, _01435_, _35846_);
  not (_01458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  nor (_01459_, _01435_, _01458_);
  or (_38927_, _01459_, _01457_);
  and (_01460_, _01109_, _36167_);
  and (_01461_, _01460_, _35815_);
  not (_01462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  nor (_01463_, _01460_, _01462_);
  or (_38928_, _01463_, _01461_);
  and (_01464_, _01460_, _35822_);
  not (_01465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor (_01466_, _01460_, _01465_);
  or (_38929_, _01466_, _01464_);
  and (_01467_, _01460_, _35826_);
  not (_01468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor (_01469_, _01460_, _01468_);
  or (_38930_, _01469_, _01467_);
  and (_01470_, _01460_, _35830_);
  not (_01471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor (_01472_, _01460_, _01471_);
  or (_38931_, _01472_, _01470_);
  and (_01473_, _01460_, _35834_);
  not (_01474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  nor (_01475_, _01460_, _01474_);
  or (_38932_, _01475_, _01473_);
  and (_01476_, _01460_, _35838_);
  not (_01477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  nor (_01478_, _01460_, _01477_);
  or (_38933_, _01478_, _01476_);
  and (_01479_, _01460_, _35842_);
  not (_01480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor (_01481_, _01460_, _01480_);
  or (_38934_, _01481_, _01479_);
  and (_01482_, _01460_, _35846_);
  not (_01483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  nor (_01484_, _01460_, _01483_);
  or (_38935_, _01484_, _01482_);
  and (_01485_, _01109_, _36193_);
  and (_01486_, _01485_, _35815_);
  not (_01487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  nor (_01488_, _01485_, _01487_);
  or (_38936_, _01488_, _01486_);
  and (_01489_, _01485_, _35822_);
  not (_01490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nor (_01491_, _01485_, _01490_);
  or (_38937_, _01491_, _01489_);
  and (_01492_, _01485_, _35826_);
  not (_01493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  nor (_01494_, _01485_, _01493_);
  or (_38938_, _01494_, _01492_);
  and (_01495_, _01485_, _35830_);
  not (_01496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor (_01497_, _01485_, _01496_);
  or (_38939_, _01497_, _01495_);
  and (_01498_, _01485_, _35834_);
  not (_01499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor (_01500_, _01485_, _01499_);
  or (_38940_, _01500_, _01498_);
  and (_01501_, _01485_, _35838_);
  not (_01502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  nor (_01503_, _01485_, _01502_);
  or (_38941_, _01503_, _01501_);
  and (_01504_, _01485_, _35842_);
  not (_01505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  nor (_01506_, _01485_, _01505_);
  or (_38942_, _01506_, _01504_);
  and (_01507_, _01485_, _35846_);
  not (_01508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  nor (_01509_, _01485_, _01508_);
  or (_38943_, _01509_, _01507_);
  and (_01510_, _00707_, _36622_);
  and (_01511_, _01510_, _35572_);
  and (_01512_, _01511_, _35815_);
  not (_01513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nor (_01514_, _01511_, _01513_);
  or (_38944_, _01514_, _01512_);
  and (_01515_, _01511_, _35822_);
  not (_01516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  nor (_01517_, _01511_, _01516_);
  or (_38945_, _01517_, _01515_);
  and (_01518_, _01511_, _35826_);
  not (_01519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nor (_01520_, _01511_, _01519_);
  or (_38946_, _01520_, _01518_);
  and (_01521_, _01511_, _35830_);
  not (_01522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  nor (_01523_, _01511_, _01522_);
  or (_38947_, _01523_, _01521_);
  and (_01524_, _01511_, _35834_);
  not (_01525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  nor (_01526_, _01511_, _01525_);
  or (_38948_, _01526_, _01524_);
  and (_01527_, _01511_, _35838_);
  not (_01528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  nor (_01529_, _01511_, _01528_);
  or (_38949_, _01529_, _01527_);
  and (_01530_, _01511_, _35842_);
  not (_01531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nor (_01532_, _01511_, _01531_);
  or (_38950_, _01532_, _01530_);
  and (_01533_, _01511_, _35846_);
  not (_01534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  nor (_01535_, _01511_, _01534_);
  or (_38951_, _01535_, _01533_);
  and (_01536_, _01510_, _35817_);
  and (_01537_, _01536_, _35815_);
  not (_01538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  nor (_01539_, _01536_, _01538_);
  or (_38952_, _01539_, _01537_);
  and (_01540_, _01536_, _35822_);
  not (_01541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nor (_01542_, _01536_, _01541_);
  or (_38953_, _01542_, _01540_);
  and (_01543_, _01536_, _35826_);
  not (_01544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nor (_01545_, _01536_, _01544_);
  or (_38954_, _01545_, _01543_);
  and (_01546_, _01536_, _35830_);
  not (_01547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  nor (_01548_, _01536_, _01547_);
  or (_38955_, _01548_, _01546_);
  and (_01549_, _01536_, _35834_);
  not (_01550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nor (_01551_, _01536_, _01550_);
  or (_38956_, _01551_, _01549_);
  and (_01552_, _01536_, _35838_);
  not (_01553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  nor (_01554_, _01536_, _01553_);
  or (_38957_, _01554_, _01552_);
  and (_01555_, _01536_, _35842_);
  not (_01556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nor (_01557_, _01536_, _01556_);
  or (_38958_, _01557_, _01555_);
  and (_01558_, _01536_, _35846_);
  not (_01559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  nor (_01560_, _01536_, _01559_);
  or (_38959_, _01560_, _01558_);
  and (_01561_, _01510_, _35851_);
  and (_01562_, _01561_, _35815_);
  not (_01563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nor (_01564_, _01561_, _01563_);
  or (_38960_, _01564_, _01562_);
  and (_01565_, _01561_, _35822_);
  not (_01566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  nor (_01567_, _01561_, _01566_);
  or (_38961_, _01567_, _01565_);
  and (_01568_, _01561_, _35826_);
  not (_01569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  nor (_01570_, _01561_, _01569_);
  or (_38962_, _01570_, _01568_);
  and (_01571_, _01561_, _35830_);
  not (_01572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nor (_01573_, _01561_, _01572_);
  or (_38963_, _01573_, _01571_);
  and (_01574_, _01561_, _35834_);
  not (_01575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  nor (_01576_, _01561_, _01575_);
  or (_38964_, _01576_, _01574_);
  and (_01577_, _01561_, _35838_);
  not (_01578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  nor (_01579_, _01561_, _01578_);
  or (_38965_, _01579_, _01577_);
  and (_01580_, _01561_, _35842_);
  not (_01581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  nor (_01582_, _01561_, _01581_);
  or (_38966_, _01582_, _01580_);
  and (_01583_, _01561_, _35846_);
  not (_01584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  nor (_01585_, _01561_, _01584_);
  or (_38967_, _01585_, _01583_);
  and (_01586_, _01510_, _35878_);
  and (_01587_, _01586_, _35815_);
  not (_01588_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nor (_01589_, _01586_, _01588_);
  or (_38968_, _01589_, _01587_);
  and (_01590_, _01586_, _35822_);
  not (_01591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nor (_01592_, _01586_, _01591_);
  or (_38969_, _01592_, _01590_);
  and (_01593_, _01586_, _35826_);
  not (_01594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nor (_01595_, _01586_, _01594_);
  or (_38970_, _01595_, _01593_);
  and (_01596_, _01586_, _35830_);
  not (_01597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  nor (_01598_, _01586_, _01597_);
  or (_38971_, _01598_, _01596_);
  and (_01599_, _01586_, _35834_);
  not (_01600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  nor (_01601_, _01586_, _01600_);
  or (_38972_, _01601_, _01599_);
  and (_01602_, _01586_, _35838_);
  not (_01603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  nor (_01604_, _01586_, _01603_);
  or (_38973_, _01604_, _01602_);
  and (_01605_, _01586_, _35842_);
  not (_01606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  nor (_01607_, _01586_, _01606_);
  or (_38974_, _01607_, _01605_);
  and (_01608_, _01586_, _35846_);
  not (_01609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nor (_01610_, _01586_, _01609_);
  or (_38975_, _01610_, _01608_);
  and (_01611_, _01510_, _35905_);
  and (_01612_, _01611_, _35815_);
  not (_01613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  nor (_01614_, _01611_, _01613_);
  or (_36936_, _01614_, _01612_);
  and (_01615_, _01611_, _35822_);
  not (_01616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  nor (_01617_, _01611_, _01616_);
  or (_36937_, _01617_, _01615_);
  and (_01618_, _01611_, _35826_);
  not (_01619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  nor (_01620_, _01611_, _01619_);
  or (_36938_, _01620_, _01618_);
  and (_01621_, _01611_, _35830_);
  not (_01622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nor (_01623_, _01611_, _01622_);
  or (_36939_, _01623_, _01621_);
  and (_01624_, _01611_, _35834_);
  not (_01625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nor (_01626_, _01611_, _01625_);
  or (_36940_, _01626_, _01624_);
  and (_01627_, _01611_, _35838_);
  not (_01628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  nor (_01629_, _01611_, _01628_);
  or (_36941_, _01629_, _01627_);
  and (_01630_, _01611_, _35842_);
  not (_01631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nor (_01632_, _01611_, _01631_);
  or (_36942_, _01632_, _01630_);
  and (_01633_, _01611_, _35846_);
  not (_01634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  nor (_01635_, _01611_, _01634_);
  or (_36943_, _01635_, _01633_);
  and (_01636_, _01510_, _35931_);
  and (_01637_, _01636_, _35815_);
  not (_01638_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nor (_01639_, _01636_, _01638_);
  or (_36944_, _01639_, _01637_);
  and (_01640_, _01636_, _35822_);
  not (_01641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nor (_01642_, _01636_, _01641_);
  or (_36945_, _01642_, _01640_);
  and (_01643_, _01636_, _35826_);
  not (_01644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nor (_01645_, _01636_, _01644_);
  or (_36946_, _01645_, _01643_);
  and (_01646_, _01636_, _35830_);
  not (_01647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nor (_01648_, _01636_, _01647_);
  or (_36947_, _01648_, _01646_);
  and (_01649_, _01636_, _35834_);
  not (_01650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  nor (_01651_, _01636_, _01650_);
  or (_36948_, _01651_, _01649_);
  and (_01652_, _01636_, _35838_);
  not (_01653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  nor (_01654_, _01636_, _01653_);
  or (_36949_, _01654_, _01652_);
  and (_01655_, _01636_, _35842_);
  not (_01656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  nor (_01657_, _01636_, _01656_);
  or (_36950_, _01657_, _01655_);
  and (_01658_, _01636_, _35846_);
  not (_01659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  nor (_01660_, _01636_, _01659_);
  or (_36951_, _01660_, _01658_);
  and (_01661_, _01510_, _35957_);
  and (_01662_, _01661_, _35815_);
  not (_01663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  nor (_01664_, _01661_, _01663_);
  or (_36952_, _01664_, _01662_);
  and (_01665_, _01661_, _35822_);
  not (_01666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  nor (_01667_, _01661_, _01666_);
  or (_36953_, _01667_, _01665_);
  and (_01668_, _01661_, _35826_);
  not (_01669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  nor (_01670_, _01661_, _01669_);
  or (_36954_, _01670_, _01668_);
  and (_01671_, _01661_, _35830_);
  not (_01672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  nor (_01673_, _01661_, _01672_);
  or (_36955_, _01673_, _01671_);
  and (_01674_, _01661_, _35834_);
  not (_01675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nor (_01676_, _01661_, _01675_);
  or (_36956_, _01676_, _01674_);
  and (_01677_, _01661_, _35838_);
  not (_01678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  nor (_01679_, _01661_, _01678_);
  or (_36957_, _01679_, _01677_);
  and (_01680_, _01661_, _35842_);
  not (_01681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nor (_01682_, _01661_, _01681_);
  or (_36958_, _01682_, _01680_);
  and (_01683_, _01661_, _35846_);
  not (_01684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  nor (_01685_, _01661_, _01684_);
  or (_36959_, _01685_, _01683_);
  and (_01686_, _01510_, _35983_);
  and (_01687_, _01686_, _35815_);
  not (_01688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nor (_01689_, _01686_, _01688_);
  or (_36960_, _01689_, _01687_);
  and (_01690_, _01686_, _35822_);
  not (_01691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  nor (_01692_, _01686_, _01691_);
  or (_36961_, _01692_, _01690_);
  and (_01693_, _01686_, _35826_);
  not (_01694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nor (_01695_, _01686_, _01694_);
  or (_36962_, _01695_, _01693_);
  and (_01696_, _01686_, _35830_);
  not (_01697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nor (_01698_, _01686_, _01697_);
  or (_36963_, _01698_, _01696_);
  and (_01699_, _01686_, _35834_);
  not (_01700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nor (_01701_, _01686_, _01700_);
  or (_36964_, _01701_, _01699_);
  and (_01702_, _01686_, _35838_);
  not (_01703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  nor (_01704_, _01686_, _01703_);
  or (_36965_, _01704_, _01702_);
  and (_01705_, _01686_, _35842_);
  not (_01706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  nor (_01707_, _01686_, _01706_);
  or (_36966_, _01707_, _01705_);
  and (_01708_, _01686_, _35846_);
  not (_01709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  nor (_01710_, _01686_, _01709_);
  or (_36967_, _01710_, _01708_);
  and (_01711_, _01510_, _36010_);
  and (_01712_, _01711_, _35815_);
  not (_01713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  nor (_01714_, _01711_, _01713_);
  or (_36968_, _01714_, _01712_);
  and (_01715_, _01711_, _35822_);
  not (_01716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nor (_01717_, _01711_, _01716_);
  or (_36969_, _01717_, _01715_);
  and (_01718_, _01711_, _35826_);
  not (_01719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  nor (_01720_, _01711_, _01719_);
  or (_36970_, _01720_, _01718_);
  and (_01721_, _01711_, _35830_);
  not (_01722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  nor (_01723_, _01711_, _01722_);
  or (_36971_, _01723_, _01721_);
  and (_01724_, _01711_, _35834_);
  not (_01725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  nor (_01726_, _01711_, _01725_);
  or (_36972_, _01726_, _01724_);
  and (_01727_, _01711_, _35838_);
  not (_01728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  nor (_01729_, _01711_, _01728_);
  or (_36973_, _01729_, _01727_);
  and (_01730_, _01711_, _35842_);
  not (_01731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nor (_01732_, _01711_, _01731_);
  or (_36974_, _01732_, _01730_);
  and (_01733_, _01711_, _35846_);
  not (_01734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  nor (_01735_, _01711_, _01734_);
  or (_36975_, _01735_, _01733_);
  and (_01736_, _01510_, _36036_);
  and (_01737_, _01736_, _35815_);
  not (_01738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nor (_01739_, _01736_, _01738_);
  or (_36976_, _01739_, _01737_);
  and (_01740_, _01736_, _35822_);
  not (_01741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  nor (_01742_, _01736_, _01741_);
  or (_36977_, _01742_, _01740_);
  and (_01743_, _01736_, _35826_);
  not (_01744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nor (_01745_, _01736_, _01744_);
  or (_36978_, _01745_, _01743_);
  and (_01746_, _01736_, _35830_);
  not (_01747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nor (_01748_, _01736_, _01747_);
  or (_36979_, _01748_, _01746_);
  and (_01749_, _01736_, _35834_);
  not (_01750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nor (_01751_, _01736_, _01750_);
  or (_36980_, _01751_, _01749_);
  and (_01752_, _01736_, _35838_);
  not (_01753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  nor (_01754_, _01736_, _01753_);
  or (_36981_, _01754_, _01752_);
  and (_01755_, _01736_, _35842_);
  not (_01756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  nor (_01757_, _01736_, _01756_);
  or (_36982_, _01757_, _01755_);
  and (_01758_, _01736_, _35846_);
  not (_01759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  nor (_01760_, _01736_, _01759_);
  or (_36983_, _01760_, _01758_);
  and (_01761_, _01510_, _36062_);
  and (_01762_, _01761_, _35815_);
  not (_01763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  nor (_01764_, _01761_, _01763_);
  or (_36984_, _01764_, _01762_);
  and (_01765_, _01761_, _35822_);
  not (_01766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor (_01767_, _01761_, _01766_);
  or (_36985_, _01767_, _01765_);
  and (_01768_, _01761_, _35826_);
  not (_01769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  nor (_01770_, _01761_, _01769_);
  or (_36986_, _01770_, _01768_);
  and (_01771_, _01761_, _35830_);
  not (_01772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  nor (_01773_, _01761_, _01772_);
  or (_36987_, _01773_, _01771_);
  and (_01774_, _01761_, _35834_);
  not (_01775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  nor (_01776_, _01761_, _01775_);
  or (_36988_, _01776_, _01774_);
  and (_01777_, _01761_, _35838_);
  not (_01778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  nor (_01779_, _01761_, _01778_);
  or (_36989_, _01779_, _01777_);
  and (_01780_, _01761_, _35842_);
  not (_01781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor (_01782_, _01761_, _01781_);
  or (_36990_, _01782_, _01780_);
  and (_01783_, _01761_, _35846_);
  not (_01784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  nor (_01785_, _01761_, _01784_);
  or (_36991_, _01785_, _01783_);
  and (_01786_, _01510_, _36088_);
  and (_01787_, _01786_, _35815_);
  not (_01788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nor (_01789_, _01786_, _01788_);
  or (_36992_, _01789_, _01787_);
  and (_01790_, _01786_, _35822_);
  not (_01791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  nor (_01792_, _01786_, _01791_);
  or (_36993_, _01792_, _01790_);
  and (_01793_, _01786_, _35826_);
  not (_01794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  nor (_01795_, _01786_, _01794_);
  or (_36994_, _01795_, _01793_);
  and (_01796_, _01786_, _35830_);
  not (_01797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor (_01798_, _01786_, _01797_);
  or (_36995_, _01798_, _01796_);
  and (_01799_, _01786_, _35834_);
  not (_01800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  nor (_01801_, _01786_, _01800_);
  or (_36996_, _01801_, _01799_);
  and (_01802_, _01786_, _35838_);
  not (_01803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  nor (_01804_, _01786_, _01803_);
  or (_36997_, _01804_, _01802_);
  and (_01805_, _01786_, _35842_);
  not (_01806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  nor (_01807_, _01786_, _01806_);
  or (_36998_, _01807_, _01805_);
  and (_01808_, _01786_, _35846_);
  not (_01809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  nor (_01810_, _01786_, _01809_);
  or (_36999_, _01810_, _01808_);
  and (_01811_, _01510_, _36115_);
  and (_01812_, _01811_, _35815_);
  not (_01813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  nor (_01814_, _01811_, _01813_);
  or (_37000_, _01814_, _01812_);
  and (_01815_, _01811_, _35822_);
  not (_01816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nor (_01817_, _01811_, _01816_);
  or (_37001_, _01817_, _01815_);
  and (_01818_, _01811_, _35826_);
  not (_01819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nor (_01820_, _01811_, _01819_);
  or (_37002_, _01820_, _01818_);
  and (_01821_, _01811_, _35830_);
  not (_01822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  nor (_01823_, _01811_, _01822_);
  or (_37003_, _01823_, _01821_);
  and (_01824_, _01811_, _35834_);
  not (_01825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nor (_01826_, _01811_, _01825_);
  or (_37004_, _01826_, _01824_);
  and (_01827_, _01811_, _35838_);
  not (_01828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  nor (_01829_, _01811_, _01828_);
  or (_37005_, _01829_, _01827_);
  and (_01830_, _01811_, _35842_);
  not (_01831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nor (_01832_, _01811_, _01831_);
  or (_37006_, _01832_, _01830_);
  and (_01833_, _01811_, _35846_);
  not (_01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  nor (_01835_, _01811_, _01834_);
  or (_37007_, _01835_, _01833_);
  and (_01836_, _01510_, _36141_);
  and (_01837_, _01836_, _35815_);
  not (_01838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  nor (_01839_, _01836_, _01838_);
  or (_37008_, _01839_, _01837_);
  and (_01840_, _01836_, _35822_);
  not (_01841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nor (_01842_, _01836_, _01841_);
  or (_37009_, _01842_, _01840_);
  and (_01843_, _01836_, _35826_);
  not (_01844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  nor (_01845_, _01836_, _01844_);
  or (_37010_, _01845_, _01843_);
  and (_01846_, _01836_, _35830_);
  not (_01847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nor (_01848_, _01836_, _01847_);
  or (_37011_, _01848_, _01846_);
  and (_01849_, _01836_, _35834_);
  not (_01850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  nor (_01851_, _01836_, _01850_);
  or (_37012_, _01851_, _01849_);
  and (_01852_, _01836_, _35838_);
  not (_01853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  nor (_01854_, _01836_, _01853_);
  or (_37013_, _01854_, _01852_);
  and (_01855_, _01836_, _35842_);
  not (_01856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nor (_01857_, _01836_, _01856_);
  or (_37014_, _01857_, _01855_);
  and (_01858_, _01836_, _35846_);
  not (_01859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  nor (_01860_, _01836_, _01859_);
  or (_37015_, _01860_, _01858_);
  and (_01861_, _01510_, _36167_);
  and (_01862_, _01861_, _35815_);
  not (_01863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor (_01864_, _01861_, _01863_);
  or (_37024_, _01864_, _01862_);
  and (_01865_, _01861_, _35822_);
  not (_01866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  nor (_01867_, _01861_, _01866_);
  or (_37025_, _01867_, _01865_);
  and (_01868_, _01861_, _35826_);
  not (_01869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor (_01870_, _01861_, _01869_);
  or (_37026_, _01870_, _01868_);
  and (_01871_, _01861_, _35830_);
  not (_01872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  nor (_01873_, _01861_, _01872_);
  or (_37027_, _01873_, _01871_);
  and (_01874_, _01861_, _35834_);
  not (_01875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor (_01876_, _01861_, _01875_);
  or (_37028_, _01876_, _01874_);
  and (_01877_, _01861_, _35838_);
  not (_01878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  nor (_01879_, _01861_, _01878_);
  or (_37029_, _01879_, _01877_);
  and (_01880_, _01861_, _35842_);
  not (_01881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  nor (_01882_, _01861_, _01881_);
  or (_37030_, _01882_, _01880_);
  and (_01883_, _01861_, _35846_);
  not (_01884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  nor (_01885_, _01861_, _01884_);
  or (_37031_, _01885_, _01883_);
  and (_01886_, _01510_, _36193_);
  and (_01887_, _01886_, _35815_);
  not (_01888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor (_01889_, _01886_, _01888_);
  or (_37032_, _01889_, _01887_);
  and (_01890_, _01886_, _35822_);
  not (_01891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor (_01892_, _01886_, _01891_);
  or (_37033_, _01892_, _01890_);
  and (_01893_, _01886_, _35826_);
  not (_01894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  nor (_01895_, _01886_, _01894_);
  or (_37034_, _01895_, _01893_);
  and (_01896_, _01886_, _35830_);
  not (_01897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor (_01898_, _01886_, _01897_);
  or (_37035_, _01898_, _01896_);
  and (_01899_, _01886_, _35834_);
  not (_01900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  nor (_01901_, _01886_, _01900_);
  or (_37036_, _01901_, _01899_);
  and (_01902_, _01886_, _35838_);
  not (_01903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor (_01904_, _01886_, _01903_);
  or (_37037_, _01904_, _01902_);
  and (_01905_, _01886_, _35842_);
  not (_01906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor (_01907_, _01886_, _01906_);
  or (_37038_, _01907_, _01905_);
  and (_01908_, _01886_, _35846_);
  not (_01909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  nor (_01910_, _01886_, _01909_);
  or (_37039_, _01910_, _01908_);
  and (_01911_, _00707_, _00304_);
  and (_01912_, _01911_, _35572_);
  and (_01913_, _01912_, _35815_);
  not (_01914_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  nor (_01915_, _01912_, _01914_);
  or (_37040_, _01915_, _01913_);
  and (_01916_, _01912_, _35822_);
  not (_01917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  nor (_01918_, _01912_, _01917_);
  or (_37041_, _01918_, _01916_);
  and (_01919_, _01912_, _35826_);
  not (_01920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nor (_01921_, _01912_, _01920_);
  or (_37042_, _01921_, _01919_);
  and (_01922_, _01912_, _35830_);
  not (_01923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  nor (_01924_, _01912_, _01923_);
  or (_37043_, _01924_, _01922_);
  and (_01925_, _01912_, _35834_);
  not (_01926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nor (_01927_, _01912_, _01926_);
  or (_37044_, _01927_, _01925_);
  and (_01928_, _01912_, _35838_);
  not (_01929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  nor (_01930_, _01912_, _01929_);
  or (_37045_, _01930_, _01928_);
  and (_01931_, _01912_, _35842_);
  not (_01932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  nor (_01933_, _01912_, _01932_);
  or (_37046_, _01933_, _01931_);
  and (_01934_, _01912_, _35846_);
  not (_01935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  nor (_01936_, _01912_, _01935_);
  or (_37047_, _01936_, _01934_);
  and (_01937_, _01911_, _35817_);
  and (_01938_, _01937_, _35815_);
  not (_01939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  nor (_01940_, _01937_, _01939_);
  or (_37048_, _01940_, _01938_);
  and (_01941_, _01937_, _35822_);
  not (_01942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  nor (_01943_, _01937_, _01942_);
  or (_37049_, _01943_, _01941_);
  and (_01944_, _01937_, _35826_);
  not (_01945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  nor (_01946_, _01937_, _01945_);
  or (_37050_, _01946_, _01944_);
  and (_01947_, _01937_, _35830_);
  not (_01948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nor (_01949_, _01937_, _01948_);
  or (_37051_, _01949_, _01947_);
  and (_01950_, _01937_, _35834_);
  not (_01951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  nor (_01952_, _01937_, _01951_);
  or (_37052_, _01952_, _01950_);
  and (_01953_, _01937_, _35838_);
  not (_01954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nor (_01955_, _01937_, _01954_);
  or (_37053_, _01955_, _01953_);
  and (_01956_, _01937_, _35842_);
  not (_01957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nor (_01958_, _01937_, _01957_);
  or (_37054_, _01958_, _01956_);
  and (_01959_, _01937_, _35846_);
  not (_01960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nor (_01961_, _01937_, _01960_);
  or (_37055_, _01961_, _01959_);
  and (_01962_, _01911_, _35851_);
  and (_01963_, _01962_, _35815_);
  not (_01964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nor (_01965_, _01962_, _01964_);
  or (_37056_, _01965_, _01963_);
  and (_01966_, _01962_, _35822_);
  not (_01967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nor (_01968_, _01962_, _01967_);
  or (_37057_, _01968_, _01966_);
  and (_01969_, _01962_, _35826_);
  not (_01970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nor (_01971_, _01962_, _01970_);
  or (_37058_, _01971_, _01969_);
  and (_01972_, _01962_, _35830_);
  not (_01973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  nor (_01974_, _01962_, _01973_);
  or (_37059_, _01974_, _01972_);
  and (_01975_, _01962_, _35834_);
  not (_01976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nor (_01977_, _01962_, _01976_);
  or (_37060_, _01977_, _01975_);
  and (_01978_, _01962_, _35838_);
  not (_01979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  nor (_01980_, _01962_, _01979_);
  or (_37061_, _01980_, _01978_);
  and (_01981_, _01962_, _35842_);
  not (_01982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  nor (_01983_, _01962_, _01982_);
  or (_37062_, _01983_, _01981_);
  and (_01984_, _01962_, _35846_);
  not (_01985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  nor (_01986_, _01962_, _01985_);
  or (_37063_, _01986_, _01984_);
  and (_01987_, _01911_, _35878_);
  and (_01988_, _01987_, _35815_);
  not (_01989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  nor (_01990_, _01987_, _01989_);
  or (_37064_, _01990_, _01988_);
  and (_01991_, _01987_, _35822_);
  not (_01992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  nor (_01993_, _01987_, _01992_);
  or (_37065_, _01993_, _01991_);
  and (_01994_, _01987_, _35826_);
  not (_01995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  nor (_01996_, _01987_, _01995_);
  or (_37066_, _01996_, _01994_);
  and (_01997_, _01987_, _35830_);
  not (_01998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  nor (_01999_, _01987_, _01998_);
  or (_37067_, _01999_, _01997_);
  and (_02000_, _01987_, _35834_);
  not (_02001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nor (_02002_, _01987_, _02001_);
  or (_37068_, _02002_, _02000_);
  and (_02003_, _01987_, _35838_);
  not (_02004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  nor (_02005_, _01987_, _02004_);
  or (_37069_, _02005_, _02003_);
  and (_02006_, _01987_, _35842_);
  not (_02007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  nor (_02008_, _01987_, _02007_);
  or (_37070_, _02008_, _02006_);
  and (_02009_, _01987_, _35846_);
  not (_02010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  nor (_02011_, _01987_, _02010_);
  or (_37071_, _02011_, _02009_);
  and (_02012_, _01911_, _35905_);
  and (_02013_, _02012_, _35815_);
  not (_02014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nor (_02015_, _02012_, _02014_);
  or (_37072_, _02015_, _02013_);
  and (_02016_, _02012_, _35822_);
  not (_02017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nor (_02018_, _02012_, _02017_);
  or (_37073_, _02018_, _02016_);
  and (_02019_, _02012_, _35826_);
  not (_02020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nor (_02021_, _02012_, _02020_);
  or (_37074_, _02021_, _02019_);
  and (_02022_, _02012_, _35830_);
  not (_02023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nor (_02024_, _02012_, _02023_);
  or (_37075_, _02024_, _02022_);
  and (_02025_, _02012_, _35834_);
  not (_02026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  nor (_02027_, _02012_, _02026_);
  or (_37076_, _02027_, _02025_);
  and (_02028_, _02012_, _35838_);
  not (_02029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  nor (_02030_, _02012_, _02029_);
  or (_37077_, _02030_, _02028_);
  and (_02031_, _02012_, _35842_);
  not (_02032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nor (_02033_, _02012_, _02032_);
  or (_37078_, _02033_, _02031_);
  and (_02034_, _02012_, _35846_);
  not (_02035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  nor (_02036_, _02012_, _02035_);
  or (_37079_, _02036_, _02034_);
  and (_02037_, _01911_, _35931_);
  and (_02038_, _02037_, _35815_);
  not (_02039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  nor (_02040_, _02037_, _02039_);
  or (_37080_, _02040_, _02038_);
  and (_02041_, _02037_, _35822_);
  not (_02042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nor (_02043_, _02037_, _02042_);
  or (_37081_, _02043_, _02041_);
  and (_02044_, _02037_, _35826_);
  not (_02045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  nor (_02046_, _02037_, _02045_);
  or (_37082_, _02046_, _02044_);
  and (_02047_, _02037_, _35830_);
  not (_02048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  nor (_02049_, _02037_, _02048_);
  or (_37083_, _02049_, _02047_);
  and (_02050_, _02037_, _35834_);
  not (_02051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nor (_02052_, _02037_, _02051_);
  or (_37084_, _02052_, _02050_);
  and (_02053_, _02037_, _35838_);
  not (_02054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  nor (_02055_, _02037_, _02054_);
  or (_37085_, _02055_, _02053_);
  and (_02056_, _02037_, _35842_);
  not (_02057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nor (_02058_, _02037_, _02057_);
  or (_37086_, _02058_, _02056_);
  and (_02059_, _02037_, _35846_);
  not (_02060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  nor (_02061_, _02037_, _02060_);
  or (_37087_, _02061_, _02059_);
  and (_02062_, _01911_, _35957_);
  and (_02063_, _02062_, _35815_);
  not (_02064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nor (_02065_, _02062_, _02064_);
  or (_37088_, _02065_, _02063_);
  and (_02066_, _02062_, _35822_);
  not (_02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  nor (_02068_, _02062_, _02067_);
  or (_37089_, _02068_, _02066_);
  and (_02069_, _02062_, _35826_);
  not (_02070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nor (_02071_, _02062_, _02070_);
  or (_37090_, _02071_, _02069_);
  and (_02072_, _02062_, _35830_);
  not (_02073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nor (_02074_, _02062_, _02073_);
  or (_37091_, _02074_, _02072_);
  and (_02075_, _02062_, _35834_);
  not (_02076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  nor (_02077_, _02062_, _02076_);
  or (_37092_, _02077_, _02075_);
  and (_02078_, _02062_, _35838_);
  not (_02079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  nor (_02080_, _02062_, _02079_);
  or (_37093_, _02080_, _02078_);
  and (_02081_, _02062_, _35842_);
  not (_02082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  nor (_02083_, _02062_, _02082_);
  or (_37094_, _02083_, _02081_);
  and (_02084_, _02062_, _35846_);
  not (_02085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  nor (_02086_, _02062_, _02085_);
  or (_37095_, _02086_, _02084_);
  and (_02087_, _01911_, _35983_);
  and (_02088_, _02087_, _35815_);
  not (_02089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  nor (_02090_, _02087_, _02089_);
  or (_37096_, _02090_, _02088_);
  and (_02091_, _02087_, _35822_);
  not (_02092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nor (_02093_, _02087_, _02092_);
  or (_37097_, _02093_, _02091_);
  and (_02094_, _02087_, _35826_);
  not (_02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nor (_02096_, _02087_, _02095_);
  or (_37098_, _02096_, _02094_);
  and (_02097_, _02087_, _35830_);
  not (_02098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  nor (_02099_, _02087_, _02098_);
  or (_37099_, _02099_, _02097_);
  and (_02100_, _02087_, _35834_);
  not (_02101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  nor (_02102_, _02087_, _02101_);
  or (_37100_, _02102_, _02100_);
  and (_02103_, _02087_, _35838_);
  not (_02104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  nor (_02105_, _02087_, _02104_);
  or (_37101_, _02105_, _02103_);
  and (_02106_, _02087_, _35842_);
  not (_02107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  nor (_02108_, _02087_, _02107_);
  or (_37102_, _02108_, _02106_);
  and (_02109_, _02087_, _35846_);
  not (_02110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  nor (_02111_, _02087_, _02110_);
  or (_37103_, _02111_, _02109_);
  and (_02112_, _01911_, _36010_);
  and (_02113_, _02112_, _35815_);
  not (_02114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor (_02115_, _02112_, _02114_);
  or (_37112_, _02115_, _02113_);
  and (_02116_, _02112_, _35822_);
  not (_02117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  nor (_02118_, _02112_, _02117_);
  or (_37113_, _02118_, _02116_);
  and (_02119_, _02112_, _35826_);
  not (_02120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  nor (_02121_, _02112_, _02120_);
  or (_37114_, _02121_, _02119_);
  and (_02122_, _02112_, _35830_);
  not (_02123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor (_02124_, _02112_, _02123_);
  or (_37115_, _02124_, _02122_);
  and (_02125_, _02112_, _35834_);
  not (_02126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor (_02127_, _02112_, _02126_);
  or (_37116_, _02127_, _02125_);
  and (_02128_, _02112_, _35838_);
  not (_02129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  nor (_02130_, _02112_, _02129_);
  or (_37117_, _02130_, _02128_);
  and (_02131_, _02112_, _35842_);
  not (_02132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor (_02133_, _02112_, _02132_);
  or (_37118_, _02133_, _02131_);
  and (_02134_, _02112_, _35846_);
  not (_02135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  nor (_02136_, _02112_, _02135_);
  or (_37119_, _02136_, _02134_);
  and (_02137_, _01911_, _36036_);
  and (_02138_, _02137_, _35815_);
  not (_02139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  nor (_02140_, _02137_, _02139_);
  or (_37120_, _02140_, _02138_);
  and (_02141_, _02137_, _35822_);
  not (_02142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor (_02143_, _02137_, _02142_);
  or (_37121_, _02143_, _02141_);
  and (_02144_, _02137_, _35826_);
  not (_02145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor (_02146_, _02137_, _02145_);
  or (_37122_, _02146_, _02144_);
  and (_02147_, _02137_, _35830_);
  not (_02148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  nor (_02149_, _02137_, _02148_);
  or (_37123_, _02149_, _02147_);
  and (_02150_, _02137_, _35834_);
  not (_02151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor (_02152_, _02137_, _02151_);
  or (_37124_, _02152_, _02150_);
  and (_02153_, _02137_, _35838_);
  not (_02154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor (_02155_, _02137_, _02154_);
  or (_37125_, _02155_, _02153_);
  and (_02156_, _02137_, _35842_);
  not (_02157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  nor (_02158_, _02137_, _02157_);
  or (_37126_, _02158_, _02156_);
  and (_02159_, _02137_, _35846_);
  not (_02160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  nor (_02161_, _02137_, _02160_);
  or (_37127_, _02161_, _02159_);
  and (_02162_, _01911_, _36062_);
  and (_02163_, _02162_, _35815_);
  not (_02164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor (_02165_, _02162_, _02164_);
  or (_37128_, _02165_, _02163_);
  and (_02166_, _02162_, _35822_);
  not (_02167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  nor (_02168_, _02162_, _02167_);
  or (_37129_, _02168_, _02166_);
  and (_02169_, _02162_, _35826_);
  not (_02170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  nor (_02171_, _02162_, _02170_);
  or (_37130_, _02171_, _02169_);
  and (_02172_, _02162_, _35830_);
  not (_02173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor (_02174_, _02162_, _02173_);
  or (_37131_, _02174_, _02172_);
  and (_02175_, _02162_, _35834_);
  not (_02176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  nor (_02177_, _02162_, _02176_);
  or (_37132_, _02177_, _02175_);
  and (_02178_, _02162_, _35838_);
  not (_02179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  nor (_02180_, _02162_, _02179_);
  or (_37133_, _02180_, _02178_);
  and (_02181_, _02162_, _35842_);
  not (_02182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor (_02183_, _02162_, _02182_);
  or (_37134_, _02183_, _02181_);
  and (_02184_, _02162_, _35846_);
  not (_02185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  nor (_02186_, _02162_, _02185_);
  or (_37135_, _02186_, _02184_);
  and (_02187_, _01911_, _36088_);
  and (_02188_, _02187_, _35815_);
  not (_02189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor (_02190_, _02187_, _02189_);
  or (_37136_, _02190_, _02188_);
  and (_02191_, _02187_, _35822_);
  not (_02192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  nor (_02193_, _02187_, _02192_);
  or (_37137_, _02193_, _02191_);
  and (_02194_, _02187_, _35826_);
  not (_02195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor (_02196_, _02187_, _02195_);
  or (_37138_, _02196_, _02194_);
  and (_02197_, _02187_, _35830_);
  not (_02198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  nor (_02199_, _02187_, _02198_);
  or (_37139_, _02199_, _02197_);
  and (_02200_, _02187_, _35834_);
  not (_02201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor (_02202_, _02187_, _02201_);
  or (_37140_, _02202_, _02200_);
  and (_02203_, _02187_, _35838_);
  not (_02204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  nor (_02205_, _02187_, _02204_);
  or (_37141_, _02205_, _02203_);
  and (_02206_, _02187_, _35842_);
  not (_02207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor (_02208_, _02187_, _02207_);
  or (_37142_, _02208_, _02206_);
  and (_02209_, _02187_, _35846_);
  not (_02210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  nor (_02211_, _02187_, _02210_);
  or (_37143_, _02211_, _02209_);
  and (_02212_, _01911_, _36115_);
  and (_02213_, _02212_, _35815_);
  not (_02214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  nor (_02215_, _02212_, _02214_);
  or (_37144_, _02215_, _02213_);
  and (_02216_, _02212_, _35822_);
  not (_02217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor (_02218_, _02212_, _02217_);
  or (_37145_, _02218_, _02216_);
  and (_02219_, _02212_, _35826_);
  not (_02220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  nor (_02221_, _02212_, _02220_);
  or (_37146_, _02221_, _02219_);
  and (_02222_, _02212_, _35830_);
  not (_02223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor (_02224_, _02212_, _02223_);
  or (_37147_, _02224_, _02222_);
  and (_02225_, _02212_, _35834_);
  not (_02226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  nor (_02227_, _02212_, _02226_);
  or (_37148_, _02227_, _02225_);
  and (_02228_, _02212_, _35838_);
  not (_02229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  nor (_02230_, _02212_, _02229_);
  or (_37149_, _02230_, _02228_);
  and (_02231_, _02212_, _35842_);
  not (_02232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  nor (_02233_, _02212_, _02232_);
  or (_37150_, _02233_, _02231_);
  and (_02234_, _02212_, _35846_);
  not (_02235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  nor (_02236_, _02212_, _02235_);
  or (_37151_, _02236_, _02234_);
  and (_02237_, _01911_, _36141_);
  and (_02238_, _02237_, _35815_);
  not (_02239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor (_02240_, _02237_, _02239_);
  or (_37152_, _02240_, _02238_);
  and (_02241_, _02237_, _35822_);
  not (_02242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor (_02243_, _02237_, _02242_);
  or (_37153_, _02243_, _02241_);
  and (_02244_, _02237_, _35826_);
  not (_02245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor (_02246_, _02237_, _02245_);
  or (_37154_, _02246_, _02244_);
  and (_02247_, _02237_, _35830_);
  not (_02248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor (_02249_, _02237_, _02248_);
  or (_37155_, _02249_, _02247_);
  and (_02250_, _02237_, _35834_);
  not (_02251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor (_02252_, _02237_, _02251_);
  or (_37156_, _02252_, _02250_);
  and (_02253_, _02237_, _35838_);
  not (_02254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  nor (_02255_, _02237_, _02254_);
  or (_37157_, _02255_, _02253_);
  and (_02256_, _02237_, _35842_);
  not (_02257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor (_02258_, _02237_, _02257_);
  or (_37158_, _02258_, _02256_);
  and (_02259_, _02237_, _35846_);
  not (_02260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  nor (_02261_, _02237_, _02260_);
  or (_37159_, _02261_, _02259_);
  and (_02262_, _01911_, _36167_);
  and (_02263_, _02262_, _35815_);
  not (_02264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  nor (_02265_, _02262_, _02264_);
  or (_37160_, _02265_, _02263_);
  and (_02266_, _02262_, _35822_);
  not (_02267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  nor (_02268_, _02262_, _02267_);
  or (_37161_, _02268_, _02266_);
  and (_02269_, _02262_, _35826_);
  not (_02270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  nor (_02271_, _02262_, _02270_);
  or (_37162_, _02271_, _02269_);
  and (_02272_, _02262_, _35830_);
  not (_02273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  nor (_02274_, _02262_, _02273_);
  or (_37163_, _02274_, _02272_);
  and (_02275_, _02262_, _35834_);
  not (_02276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  nor (_02277_, _02262_, _02276_);
  or (_37164_, _02277_, _02275_);
  and (_02278_, _02262_, _35838_);
  not (_02279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor (_02280_, _02262_, _02279_);
  or (_37165_, _02280_, _02278_);
  and (_02281_, _02262_, _35842_);
  not (_02282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  nor (_02283_, _02262_, _02282_);
  or (_37166_, _02283_, _02281_);
  and (_02284_, _02262_, _35846_);
  not (_02285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  nor (_02286_, _02262_, _02285_);
  or (_37167_, _02286_, _02284_);
  and (_02287_, _01911_, _36193_);
  and (_02288_, _02287_, _35815_);
  not (_02289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  nor (_02290_, _02287_, _02289_);
  or (_37168_, _02290_, _02288_);
  and (_02291_, _02287_, _35822_);
  not (_02292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor (_02293_, _02287_, _02292_);
  or (_37169_, _02293_, _02291_);
  and (_02294_, _02287_, _35826_);
  not (_02295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  nor (_02296_, _02287_, _02295_);
  or (_37170_, _02296_, _02294_);
  and (_02297_, _02287_, _35830_);
  not (_02298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  nor (_02299_, _02287_, _02298_);
  or (_37171_, _02299_, _02297_);
  and (_02300_, _02287_, _35834_);
  not (_02301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  nor (_02302_, _02287_, _02301_);
  or (_37172_, _02302_, _02300_);
  and (_02303_, _02287_, _35838_);
  not (_02304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  nor (_02305_, _02287_, _02304_);
  or (_37173_, _02305_, _02303_);
  and (_02306_, _02287_, _35842_);
  not (_02307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor (_02308_, _02287_, _02307_);
  or (_37174_, _02308_, _02306_);
  and (_02309_, _02287_, _35846_);
  not (_02310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  nor (_02311_, _02287_, _02310_);
  or (_37175_, _02311_, _02309_);
  and (_02312_, _34784_, _33632_);
  and (_02313_, _02312_, _35575_);
  and (_02314_, _02313_, _35572_);
  and (_02315_, _02314_, _35815_);
  not (_02316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nor (_02317_, _02314_, _02316_);
  or (_37176_, _02317_, _02315_);
  and (_02318_, _02314_, _35822_);
  not (_02319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  nor (_02320_, _02314_, _02319_);
  or (_37177_, _02320_, _02318_);
  and (_02321_, _02314_, _35826_);
  not (_02322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nor (_02323_, _02314_, _02322_);
  or (_37178_, _02323_, _02321_);
  and (_02324_, _02314_, _35830_);
  not (_02325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nor (_02326_, _02314_, _02325_);
  or (_37179_, _02326_, _02324_);
  and (_02327_, _02314_, _35834_);
  not (_02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nor (_02329_, _02314_, _02328_);
  or (_37180_, _02329_, _02327_);
  and (_02330_, _02314_, _35838_);
  not (_02331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  nor (_02332_, _02314_, _02331_);
  or (_37181_, _02332_, _02330_);
  and (_02333_, _02314_, _35842_);
  not (_02334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  nor (_02335_, _02314_, _02334_);
  or (_37182_, _02335_, _02333_);
  and (_02336_, _02314_, _35846_);
  not (_02337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  nor (_02338_, _02314_, _02337_);
  or (_37183_, _02338_, _02336_);
  and (_02339_, _02313_, _35817_);
  and (_02340_, _02339_, _35815_);
  not (_02341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nor (_02342_, _02339_, _02341_);
  or (_37184_, _02342_, _02340_);
  and (_02343_, _02339_, _35822_);
  not (_02344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nor (_02345_, _02339_, _02344_);
  or (_37185_, _02345_, _02343_);
  and (_02346_, _02339_, _35826_);
  not (_02347_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  nor (_02348_, _02339_, _02347_);
  or (_37186_, _02348_, _02346_);
  and (_02349_, _02339_, _35830_);
  not (_02350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nor (_02351_, _02339_, _02350_);
  or (_37187_, _02351_, _02349_);
  and (_02352_, _02339_, _35834_);
  not (_02353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  nor (_02354_, _02339_, _02353_);
  or (_37188_, _02354_, _02352_);
  and (_02355_, _02339_, _35838_);
  not (_02356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  nor (_02357_, _02339_, _02356_);
  or (_37189_, _02357_, _02355_);
  and (_02358_, _02339_, _35842_);
  not (_02359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nor (_02360_, _02339_, _02359_);
  or (_37190_, _02360_, _02358_);
  and (_02361_, _02339_, _35846_);
  not (_02362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nor (_02363_, _02339_, _02362_);
  or (_37191_, _02363_, _02361_);
  and (_02364_, _02313_, _35851_);
  and (_02365_, _02364_, _35815_);
  not (_02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  nor (_02367_, _02364_, _02366_);
  or (_37200_, _02367_, _02365_);
  and (_02368_, _02364_, _35822_);
  not (_02369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  nor (_02370_, _02364_, _02369_);
  or (_37201_, _02370_, _02368_);
  and (_02371_, _02364_, _35826_);
  not (_02372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nor (_02373_, _02364_, _02372_);
  or (_37202_, _02373_, _02371_);
  and (_02374_, _02364_, _35830_);
  not (_02375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  nor (_02376_, _02364_, _02375_);
  or (_37203_, _02376_, _02374_);
  and (_02377_, _02364_, _35834_);
  not (_02378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nor (_02379_, _02364_, _02378_);
  or (_37204_, _02379_, _02377_);
  and (_02380_, _02364_, _35838_);
  not (_02381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nor (_02382_, _02364_, _02381_);
  or (_37205_, _02382_, _02380_);
  and (_02383_, _02364_, _35842_);
  not (_02384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  nor (_02385_, _02364_, _02384_);
  or (_37206_, _02385_, _02383_);
  and (_02386_, _02364_, _35846_);
  not (_02387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nor (_02388_, _02364_, _02387_);
  or (_37207_, _02388_, _02386_);
  and (_02389_, _02313_, _35878_);
  and (_02390_, _02389_, _35815_);
  not (_02391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nor (_02392_, _02389_, _02391_);
  or (_37208_, _02392_, _02390_);
  and (_02393_, _02389_, _35822_);
  not (_02394_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nor (_02395_, _02389_, _02394_);
  or (_37209_, _02395_, _02393_);
  and (_02396_, _02389_, _35826_);
  not (_02397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nor (_02398_, _02389_, _02397_);
  or (_37210_, _02398_, _02396_);
  and (_02399_, _02389_, _35830_);
  not (_02400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  nor (_02401_, _02389_, _02400_);
  or (_37211_, _02401_, _02399_);
  and (_02402_, _02389_, _35834_);
  not (_02403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  nor (_02404_, _02389_, _02403_);
  or (_37212_, _02404_, _02402_);
  and (_02405_, _02389_, _35838_);
  not (_02406_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  nor (_02407_, _02389_, _02406_);
  or (_37213_, _02407_, _02405_);
  and (_02408_, _02389_, _35842_);
  not (_02409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nor (_02410_, _02389_, _02409_);
  or (_37214_, _02410_, _02408_);
  and (_02411_, _02389_, _35846_);
  not (_02412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nor (_02413_, _02389_, _02412_);
  or (_37215_, _02413_, _02411_);
  and (_02414_, _02313_, _35905_);
  and (_02415_, _02414_, _35815_);
  not (_02416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  nor (_02417_, _02414_, _02416_);
  or (_37216_, _02417_, _02415_);
  and (_02418_, _02414_, _35822_);
  not (_02419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  nor (_02420_, _02414_, _02419_);
  or (_37217_, _02420_, _02418_);
  and (_02421_, _02414_, _35826_);
  not (_02422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  nor (_02423_, _02414_, _02422_);
  or (_37218_, _02423_, _02421_);
  and (_02424_, _02414_, _35830_);
  not (_02425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nor (_02426_, _02414_, _02425_);
  or (_37219_, _02426_, _02424_);
  and (_02427_, _02414_, _35834_);
  not (_02428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nor (_02429_, _02414_, _02428_);
  or (_37220_, _02429_, _02427_);
  and (_02430_, _02414_, _35838_);
  not (_02431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  nor (_02432_, _02414_, _02431_);
  or (_37221_, _02432_, _02430_);
  and (_02433_, _02414_, _35842_);
  not (_02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nor (_02435_, _02414_, _02434_);
  or (_37222_, _02435_, _02433_);
  and (_02436_, _02414_, _35846_);
  not (_02437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nor (_02438_, _02414_, _02437_);
  or (_37223_, _02438_, _02436_);
  and (_02439_, _02313_, _35931_);
  and (_02440_, _02439_, _35815_);
  not (_02441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nor (_02442_, _02439_, _02441_);
  or (_37224_, _02442_, _02440_);
  and (_02443_, _02439_, _35822_);
  not (_02444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  nor (_02445_, _02439_, _02444_);
  or (_37225_, _02445_, _02443_);
  and (_02446_, _02439_, _35826_);
  not (_02447_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nor (_02448_, _02439_, _02447_);
  or (_37226_, _02448_, _02446_);
  and (_02449_, _02439_, _35830_);
  not (_02450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  nor (_02451_, _02439_, _02450_);
  or (_37227_, _02451_, _02449_);
  and (_02452_, _02439_, _35834_);
  not (_02453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nor (_02454_, _02439_, _02453_);
  or (_37228_, _02454_, _02452_);
  and (_02455_, _02439_, _35838_);
  not (_02456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  nor (_02457_, _02439_, _02456_);
  or (_37229_, _02457_, _02455_);
  and (_02458_, _02439_, _35842_);
  not (_02459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  nor (_02460_, _02439_, _02459_);
  or (_37230_, _02460_, _02458_);
  and (_02461_, _02439_, _35846_);
  not (_02462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nor (_02463_, _02439_, _02462_);
  or (_37231_, _02463_, _02461_);
  and (_02464_, _02313_, _35957_);
  and (_02465_, _02464_, _35815_);
  not (_02466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  nor (_02467_, _02464_, _02466_);
  or (_37232_, _02467_, _02465_);
  and (_02468_, _02464_, _35822_);
  not (_02469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nor (_02470_, _02464_, _02469_);
  or (_37233_, _02470_, _02468_);
  and (_02471_, _02464_, _35826_);
  not (_02472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  nor (_02473_, _02464_, _02472_);
  or (_37234_, _02473_, _02471_);
  and (_02474_, _02464_, _35830_);
  not (_02475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nor (_02476_, _02464_, _02475_);
  or (_37235_, _02476_, _02474_);
  and (_02477_, _02464_, _35834_);
  not (_02478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  nor (_02479_, _02464_, _02478_);
  or (_37236_, _02479_, _02477_);
  and (_02480_, _02464_, _35838_);
  not (_02481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  nor (_02482_, _02464_, _02481_);
  or (_37237_, _02482_, _02480_);
  and (_02483_, _02464_, _35842_);
  not (_02484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nor (_02485_, _02464_, _02484_);
  or (_37238_, _02485_, _02483_);
  and (_02486_, _02464_, _35846_);
  not (_02487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nor (_02488_, _02464_, _02487_);
  or (_37239_, _02488_, _02486_);
  and (_02489_, _02313_, _35983_);
  and (_02490_, _02489_, _35815_);
  not (_02491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  nor (_02492_, _02489_, _02491_);
  or (_37240_, _02492_, _02490_);
  and (_02493_, _02489_, _35822_);
  not (_02494_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  nor (_02495_, _02489_, _02494_);
  or (_37241_, _02495_, _02493_);
  and (_02496_, _02489_, _35826_);
  not (_02497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  nor (_02498_, _02489_, _02497_);
  or (_37242_, _02498_, _02496_);
  and (_02499_, _02489_, _35830_);
  not (_02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  nor (_02501_, _02489_, _02500_);
  or (_37243_, _02501_, _02499_);
  and (_02502_, _02489_, _35834_);
  not (_02503_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  nor (_02504_, _02489_, _02503_);
  or (_37244_, _02504_, _02502_);
  and (_02505_, _02489_, _35838_);
  not (_02506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  nor (_02507_, _02489_, _02506_);
  or (_37245_, _02507_, _02505_);
  and (_02508_, _02489_, _35842_);
  not (_02509_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nor (_02510_, _02489_, _02509_);
  or (_37246_, _02510_, _02508_);
  and (_02511_, _02489_, _35846_);
  not (_02512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nor (_02513_, _02489_, _02512_);
  or (_37247_, _02513_, _02511_);
  and (_02514_, _02313_, _36010_);
  and (_02515_, _02514_, _35815_);
  not (_02516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nor (_02517_, _02514_, _02516_);
  or (_37248_, _02517_, _02515_);
  and (_02518_, _02514_, _35822_);
  not (_02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nor (_02520_, _02514_, _02519_);
  or (_37249_, _02520_, _02518_);
  and (_02521_, _02514_, _35826_);
  not (_02522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nor (_02523_, _02514_, _02522_);
  or (_37250_, _02523_, _02521_);
  and (_02524_, _02514_, _35830_);
  not (_02525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nor (_02526_, _02514_, _02525_);
  or (_37251_, _02526_, _02524_);
  and (_02527_, _02514_, _35834_);
  not (_02528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nor (_02529_, _02514_, _02528_);
  or (_37252_, _02529_, _02527_);
  and (_02530_, _02514_, _35838_);
  not (_02531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  nor (_02532_, _02514_, _02531_);
  or (_37253_, _02532_, _02530_);
  and (_02533_, _02514_, _35842_);
  not (_02534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nor (_02535_, _02514_, _02534_);
  or (_37254_, _02535_, _02533_);
  and (_02536_, _02514_, _35846_);
  not (_02537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nor (_02538_, _02514_, _02537_);
  or (_37255_, _02538_, _02536_);
  and (_02539_, _02313_, _36036_);
  and (_02540_, _02539_, _35815_);
  not (_02541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nor (_02542_, _02539_, _02541_);
  or (_37256_, _02542_, _02540_);
  and (_02543_, _02539_, _35822_);
  not (_02544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nor (_02545_, _02539_, _02544_);
  or (_37257_, _02545_, _02543_);
  and (_02546_, _02539_, _35826_);
  not (_02547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nor (_02548_, _02539_, _02547_);
  or (_37258_, _02548_, _02546_);
  and (_02549_, _02539_, _35830_);
  not (_02550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nor (_02551_, _02539_, _02550_);
  or (_37259_, _02551_, _02549_);
  and (_02552_, _02539_, _35834_);
  not (_02553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  nor (_02554_, _02539_, _02553_);
  or (_37260_, _02554_, _02552_);
  and (_02555_, _02539_, _35838_);
  not (_02556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  nor (_02557_, _02539_, _02556_);
  or (_37261_, _02557_, _02555_);
  and (_02558_, _02539_, _35842_);
  not (_02559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nor (_02560_, _02539_, _02559_);
  or (_37262_, _02560_, _02558_);
  and (_02561_, _02539_, _35846_);
  not (_02562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  nor (_02563_, _02539_, _02562_);
  or (_37263_, _02563_, _02561_);
  and (_02564_, _02313_, _36062_);
  and (_02565_, _02564_, _35815_);
  not (_02566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  nor (_02567_, _02564_, _02566_);
  or (_37264_, _02567_, _02565_);
  and (_02568_, _02564_, _35822_);
  not (_02569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  nor (_02570_, _02564_, _02569_);
  or (_37265_, _02570_, _02568_);
  and (_02571_, _02564_, _35826_);
  not (_02572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  nor (_02573_, _02564_, _02572_);
  or (_37266_, _02573_, _02571_);
  and (_02574_, _02564_, _35830_);
  not (_02575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  nor (_02576_, _02564_, _02575_);
  or (_37267_, _02576_, _02574_);
  and (_02577_, _02564_, _35834_);
  not (_02578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor (_02579_, _02564_, _02578_);
  or (_37268_, _02579_, _02577_);
  and (_02580_, _02564_, _35838_);
  not (_02581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  nor (_02582_, _02564_, _02581_);
  or (_37269_, _02582_, _02580_);
  and (_02583_, _02564_, _35842_);
  not (_02584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  nor (_02585_, _02564_, _02584_);
  or (_37270_, _02585_, _02583_);
  and (_02586_, _02564_, _35846_);
  not (_02587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nor (_02588_, _02564_, _02587_);
  or (_37271_, _02588_, _02586_);
  and (_02589_, _02313_, _36088_);
  and (_02590_, _02589_, _35815_);
  not (_02591_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  nor (_02592_, _02589_, _02591_);
  or (_37272_, _02592_, _02590_);
  and (_02593_, _02589_, _35822_);
  not (_02594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor (_02595_, _02589_, _02594_);
  or (_37273_, _02595_, _02593_);
  and (_02596_, _02589_, _35826_);
  not (_02597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor (_02598_, _02589_, _02597_);
  or (_37274_, _02598_, _02596_);
  and (_02599_, _02589_, _35830_);
  not (_02600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  nor (_02601_, _02589_, _02600_);
  or (_37275_, _02601_, _02599_);
  and (_02602_, _02589_, _35834_);
  not (_02603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  nor (_02604_, _02589_, _02603_);
  or (_37276_, _02604_, _02602_);
  and (_02605_, _02589_, _35838_);
  not (_02606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  nor (_02607_, _02589_, _02606_);
  or (_37277_, _02607_, _02605_);
  and (_02608_, _02589_, _35842_);
  not (_02609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nor (_02610_, _02589_, _02609_);
  or (_37278_, _02610_, _02608_);
  and (_02611_, _02589_, _35846_);
  not (_02612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nor (_02613_, _02589_, _02612_);
  or (_37279_, _02613_, _02611_);
  and (_02614_, _02313_, _36115_);
  and (_02615_, _02614_, _35815_);
  not (_02616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nor (_02617_, _02614_, _02616_);
  or (_37288_, _02617_, _02615_);
  and (_02618_, _02614_, _35822_);
  not (_02619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  nor (_02620_, _02614_, _02619_);
  or (_37289_, _02620_, _02618_);
  and (_02621_, _02614_, _35826_);
  not (_02622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  nor (_02623_, _02614_, _02622_);
  or (_37290_, _02623_, _02621_);
  and (_02624_, _02614_, _35830_);
  not (_02625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nor (_02626_, _02614_, _02625_);
  or (_37291_, _02626_, _02624_);
  and (_02627_, _02614_, _35834_);
  not (_02628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nor (_02629_, _02614_, _02628_);
  or (_37292_, _02629_, _02627_);
  and (_02630_, _02614_, _35838_);
  not (_02631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  nor (_02632_, _02614_, _02631_);
  or (_37293_, _02632_, _02630_);
  and (_02633_, _02614_, _35842_);
  not (_02634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nor (_02635_, _02614_, _02634_);
  or (_37294_, _02635_, _02633_);
  and (_02636_, _02614_, _35846_);
  not (_02637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nor (_02638_, _02614_, _02637_);
  or (_37295_, _02638_, _02636_);
  and (_02639_, _02313_, _36141_);
  and (_02640_, _02639_, _35815_);
  not (_02641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nor (_02642_, _02639_, _02641_);
  or (_37296_, _02642_, _02640_);
  and (_02643_, _02639_, _35822_);
  not (_02644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nor (_02645_, _02639_, _02644_);
  or (_37297_, _02645_, _02643_);
  and (_02646_, _02639_, _35826_);
  not (_02647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nor (_02648_, _02639_, _02647_);
  or (_37298_, _02648_, _02646_);
  and (_02649_, _02639_, _35830_);
  not (_02650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nor (_02651_, _02639_, _02650_);
  or (_37299_, _02651_, _02649_);
  and (_02652_, _02639_, _35834_);
  not (_02653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  nor (_02654_, _02639_, _02653_);
  or (_37300_, _02654_, _02652_);
  and (_02655_, _02639_, _35838_);
  not (_02656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  nor (_02657_, _02639_, _02656_);
  or (_37301_, _02657_, _02655_);
  and (_02658_, _02639_, _35842_);
  not (_02659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nor (_02660_, _02639_, _02659_);
  or (_37302_, _02660_, _02658_);
  and (_02661_, _02639_, _35846_);
  not (_02662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nor (_02663_, _02639_, _02662_);
  or (_37303_, _02663_, _02661_);
  and (_02664_, _02313_, _36167_);
  and (_02665_, _02664_, _35815_);
  not (_02666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  nor (_02667_, _02664_, _02666_);
  or (_37304_, _02667_, _02665_);
  and (_02668_, _02664_, _35822_);
  not (_02669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  nor (_02670_, _02664_, _02669_);
  or (_37305_, _02670_, _02668_);
  and (_02671_, _02664_, _35826_);
  not (_02672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  nor (_02673_, _02664_, _02672_);
  or (_37306_, _02673_, _02671_);
  and (_02674_, _02664_, _35830_);
  not (_02675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  nor (_02676_, _02664_, _02675_);
  or (_37307_, _02676_, _02674_);
  and (_02677_, _02664_, _35834_);
  not (_02678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor (_02679_, _02664_, _02678_);
  or (_37308_, _02679_, _02677_);
  and (_02680_, _02664_, _35838_);
  not (_02681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  nor (_02682_, _02664_, _02681_);
  or (_37309_, _02682_, _02680_);
  and (_02683_, _02664_, _35842_);
  not (_02684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nor (_02685_, _02664_, _02684_);
  or (_37310_, _02685_, _02683_);
  and (_02686_, _02664_, _35846_);
  not (_02687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nor (_02688_, _02664_, _02687_);
  or (_37311_, _02688_, _02686_);
  and (_02689_, _02313_, _36193_);
  and (_02690_, _02689_, _35815_);
  not (_02691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor (_02692_, _02689_, _02691_);
  or (_37312_, _02692_, _02690_);
  and (_02693_, _02689_, _35822_);
  not (_02694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor (_02695_, _02689_, _02694_);
  or (_37313_, _02695_, _02693_);
  and (_02696_, _02689_, _35826_);
  not (_02697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor (_02698_, _02689_, _02697_);
  or (_37314_, _02698_, _02696_);
  and (_02699_, _02689_, _35830_);
  not (_02700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  nor (_02701_, _02689_, _02700_);
  or (_37315_, _02701_, _02699_);
  and (_02702_, _02689_, _35834_);
  not (_02703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nor (_02704_, _02689_, _02703_);
  or (_37316_, _02704_, _02702_);
  and (_02705_, _02689_, _35838_);
  not (_02706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  nor (_02707_, _02689_, _02706_);
  or (_37317_, _02707_, _02705_);
  and (_02708_, _02689_, _35842_);
  not (_02709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor (_02710_, _02689_, _02709_);
  or (_37318_, _02710_, _02708_);
  and (_02711_, _02689_, _35846_);
  not (_02712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nor (_02713_, _02689_, _02712_);
  or (_37319_, _02713_, _02711_);
  and (_02714_, _36220_, _33632_);
  and (_02715_, _02714_, _35572_);
  and (_02716_, _02715_, _35815_);
  not (_02717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  nor (_02718_, _02715_, _02717_);
  or (_37320_, _02718_, _02716_);
  and (_02719_, _02715_, _35822_);
  not (_02720_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  nor (_02721_, _02715_, _02720_);
  or (_37321_, _02721_, _02719_);
  and (_02722_, _02715_, _35826_);
  not (_02723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  nor (_02724_, _02715_, _02723_);
  or (_37322_, _02724_, _02722_);
  and (_02725_, _02715_, _35830_);
  not (_02726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nor (_02727_, _02715_, _02726_);
  or (_37323_, _02727_, _02725_);
  and (_02728_, _02715_, _35834_);
  not (_02729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  nor (_02730_, _02715_, _02729_);
  or (_37324_, _02730_, _02728_);
  and (_02731_, _02715_, _35838_);
  not (_02732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  nor (_02733_, _02715_, _02732_);
  or (_37325_, _02733_, _02731_);
  and (_02734_, _02715_, _35842_);
  not (_02735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  nor (_02736_, _02715_, _02735_);
  or (_37326_, _02736_, _02734_);
  and (_02737_, _02715_, _35846_);
  not (_02738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  nor (_02739_, _02715_, _02738_);
  or (_37327_, _02739_, _02737_);
  and (_02740_, _02714_, _35817_);
  and (_02741_, _02740_, _35815_);
  not (_02742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nor (_02743_, _02740_, _02742_);
  or (_37328_, _02743_, _02741_);
  and (_02744_, _02740_, _35822_);
  not (_02745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nor (_02746_, _02740_, _02745_);
  or (_37329_, _02746_, _02744_);
  and (_02747_, _02740_, _35826_);
  not (_02748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nor (_02749_, _02740_, _02748_);
  or (_37330_, _02749_, _02747_);
  and (_02750_, _02740_, _35830_);
  not (_02751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nor (_02752_, _02740_, _02751_);
  or (_37331_, _02752_, _02750_);
  and (_02753_, _02740_, _35834_);
  not (_02754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nor (_02755_, _02740_, _02754_);
  or (_37332_, _02755_, _02753_);
  and (_02756_, _02740_, _35838_);
  not (_02757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  nor (_02758_, _02740_, _02757_);
  or (_37333_, _02758_, _02756_);
  and (_02759_, _02740_, _35842_);
  not (_02760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  nor (_02761_, _02740_, _02760_);
  or (_37334_, _02761_, _02759_);
  and (_02762_, _02740_, _35846_);
  not (_02763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  nor (_02764_, _02740_, _02763_);
  or (_37335_, _02764_, _02762_);
  and (_02765_, _02714_, _35851_);
  and (_02766_, _02765_, _35815_);
  not (_02767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  nor (_02768_, _02765_, _02767_);
  or (_37336_, _02768_, _02766_);
  and (_02769_, _02765_, _35822_);
  not (_02770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  nor (_02771_, _02765_, _02770_);
  or (_37337_, _02771_, _02769_);
  and (_02772_, _02765_, _35826_);
  not (_02773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  nor (_02774_, _02765_, _02773_);
  or (_37338_, _02774_, _02772_);
  and (_02775_, _02765_, _35830_);
  not (_02776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  nor (_02777_, _02765_, _02776_);
  or (_37339_, _02777_, _02775_);
  and (_02778_, _02765_, _35834_);
  not (_02779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  nor (_02780_, _02765_, _02779_);
  or (_37340_, _02780_, _02778_);
  and (_02781_, _02765_, _35838_);
  not (_02782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  nor (_02783_, _02765_, _02782_);
  or (_37341_, _02783_, _02781_);
  and (_02784_, _02765_, _35842_);
  not (_02785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nor (_02786_, _02765_, _02785_);
  or (_37342_, _02786_, _02784_);
  and (_02787_, _02765_, _35846_);
  not (_02788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  nor (_02789_, _02765_, _02788_);
  or (_37343_, _02789_, _02787_);
  and (_02790_, _02714_, _35878_);
  and (_02791_, _02790_, _35815_);
  not (_02792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nor (_02793_, _02790_, _02792_);
  or (_37344_, _02793_, _02791_);
  and (_02794_, _02790_, _35822_);
  not (_02795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nor (_02796_, _02790_, _02795_);
  or (_37345_, _02796_, _02794_);
  and (_02797_, _02790_, _35826_);
  not (_02798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  nor (_02799_, _02790_, _02798_);
  or (_37346_, _02799_, _02797_);
  and (_02800_, _02790_, _35830_);
  not (_02801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nor (_02802_, _02790_, _02801_);
  or (_37347_, _02802_, _02800_);
  and (_02803_, _02790_, _35834_);
  not (_02804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nor (_02805_, _02790_, _02804_);
  or (_37348_, _02805_, _02803_);
  and (_02806_, _02790_, _35838_);
  not (_02807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  nor (_02808_, _02790_, _02807_);
  or (_37349_, _02808_, _02806_);
  and (_02809_, _02790_, _35842_);
  not (_02810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nor (_02811_, _02790_, _02810_);
  or (_37350_, _02811_, _02809_);
  and (_02812_, _02790_, _35846_);
  not (_02813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  nor (_02814_, _02790_, _02813_);
  or (_37351_, _02814_, _02812_);
  and (_02815_, _02714_, _35905_);
  and (_02816_, _02815_, _35815_);
  not (_02817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  nor (_02818_, _02815_, _02817_);
  or (_37352_, _02818_, _02816_);
  and (_02819_, _02815_, _35822_);
  not (_02820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  nor (_02821_, _02815_, _02820_);
  or (_37353_, _02821_, _02819_);
  and (_02822_, _02815_, _35826_);
  not (_02823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nor (_02824_, _02815_, _02823_);
  or (_37354_, _02824_, _02822_);
  and (_02825_, _02815_, _35830_);
  not (_02826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  nor (_02827_, _02815_, _02826_);
  or (_37355_, _02827_, _02825_);
  and (_02828_, _02815_, _35834_);
  not (_02829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  nor (_02830_, _02815_, _02829_);
  or (_37356_, _02830_, _02828_);
  and (_02831_, _02815_, _35838_);
  not (_02832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  nor (_02833_, _02815_, _02832_);
  or (_37357_, _02833_, _02831_);
  and (_02834_, _02815_, _35842_);
  not (_02835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  nor (_02836_, _02815_, _02835_);
  or (_37358_, _02836_, _02834_);
  and (_02837_, _02815_, _35846_);
  not (_02838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  nor (_02839_, _02815_, _02838_);
  or (_37359_, _02839_, _02837_);
  and (_02840_, _02714_, _35931_);
  and (_02841_, _02840_, _35815_);
  not (_02842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nor (_02843_, _02840_, _02842_);
  or (_37360_, _02843_, _02841_);
  and (_02844_, _02840_, _35822_);
  not (_02845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  nor (_02846_, _02840_, _02845_);
  or (_37361_, _02846_, _02844_);
  and (_02847_, _02840_, _35826_);
  not (_02848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nor (_02849_, _02840_, _02848_);
  or (_37362_, _02849_, _02847_);
  and (_02850_, _02840_, _35830_);
  not (_02851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nor (_02852_, _02840_, _02851_);
  or (_37363_, _02852_, _02850_);
  and (_02853_, _02840_, _35834_);
  not (_02854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  nor (_02855_, _02840_, _02854_);
  or (_37364_, _02855_, _02853_);
  and (_02856_, _02840_, _35838_);
  not (_02857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  nor (_02858_, _02840_, _02857_);
  or (_37365_, _02858_, _02856_);
  and (_02859_, _02840_, _35842_);
  not (_02860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  nor (_02861_, _02840_, _02860_);
  or (_37366_, _02861_, _02859_);
  and (_02862_, _02840_, _35846_);
  not (_02863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  nor (_02864_, _02840_, _02863_);
  or (_37367_, _02864_, _02862_);
  and (_02865_, _02714_, _35957_);
  and (_02866_, _02865_, _35815_);
  not (_02867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  nor (_02868_, _02865_, _02867_);
  or (_37376_, _02868_, _02866_);
  and (_02869_, _02865_, _35822_);
  not (_02870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nor (_02871_, _02865_, _02870_);
  or (_37377_, _02871_, _02869_);
  and (_02872_, _02865_, _35826_);
  not (_02873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  nor (_02874_, _02865_, _02873_);
  or (_37378_, _02874_, _02872_);
  and (_02875_, _02865_, _35830_);
  not (_02876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  nor (_02877_, _02865_, _02876_);
  or (_37379_, _02877_, _02875_);
  and (_02878_, _02865_, _35834_);
  not (_02879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nor (_02880_, _02865_, _02879_);
  or (_37380_, _02880_, _02878_);
  and (_02881_, _02865_, _35838_);
  not (_02882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  nor (_02883_, _02865_, _02882_);
  or (_37381_, _02883_, _02881_);
  and (_02884_, _02865_, _35842_);
  not (_02885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nor (_02886_, _02865_, _02885_);
  or (_37382_, _02886_, _02884_);
  and (_02887_, _02865_, _35846_);
  not (_02888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  nor (_02889_, _02865_, _02888_);
  or (_37383_, _02889_, _02887_);
  and (_02890_, _02714_, _35983_);
  and (_02891_, _02890_, _35815_);
  not (_02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nor (_02893_, _02890_, _02892_);
  or (_37384_, _02893_, _02891_);
  and (_02894_, _02890_, _35822_);
  not (_02895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nor (_02896_, _02890_, _02895_);
  or (_37385_, _02896_, _02894_);
  and (_02897_, _02890_, _35826_);
  not (_02898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  nor (_02899_, _02890_, _02898_);
  or (_37386_, _02899_, _02897_);
  and (_02900_, _02890_, _35830_);
  not (_02901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nor (_02902_, _02890_, _02901_);
  or (_37387_, _02902_, _02900_);
  and (_02903_, _02890_, _35834_);
  not (_02904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nor (_02905_, _02890_, _02904_);
  or (_37388_, _02905_, _02903_);
  and (_02906_, _02890_, _35838_);
  not (_02907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  nor (_02908_, _02890_, _02907_);
  or (_37389_, _02908_, _02906_);
  and (_02909_, _02890_, _35842_);
  not (_02910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nor (_02911_, _02890_, _02910_);
  or (_37390_, _02911_, _02909_);
  and (_02912_, _02890_, _35846_);
  not (_02913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  nor (_02914_, _02890_, _02913_);
  or (_37391_, _02914_, _02912_);
  and (_02915_, _02714_, _36010_);
  and (_02916_, _02915_, _35815_);
  not (_02917_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  nor (_02918_, _02915_, _02917_);
  or (_37392_, _02918_, _02916_);
  and (_02919_, _02915_, _35822_);
  not (_02920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  nor (_02921_, _02915_, _02920_);
  or (_37393_, _02921_, _02919_);
  and (_02922_, _02915_, _35826_);
  not (_02923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor (_02924_, _02915_, _02923_);
  or (_37394_, _02924_, _02922_);
  and (_02925_, _02915_, _35830_);
  not (_02926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  nor (_02927_, _02915_, _02926_);
  or (_37395_, _02927_, _02925_);
  and (_02928_, _02915_, _35834_);
  not (_02929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  nor (_02930_, _02915_, _02929_);
  or (_37396_, _02930_, _02928_);
  and (_02931_, _02915_, _35838_);
  not (_02932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  nor (_02933_, _02915_, _02932_);
  or (_37397_, _02933_, _02931_);
  and (_02934_, _02915_, _35842_);
  not (_02935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  nor (_02936_, _02915_, _02935_);
  or (_37398_, _02936_, _02934_);
  and (_02937_, _02915_, _35846_);
  not (_02938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  nor (_02939_, _02915_, _02938_);
  or (_37399_, _02939_, _02937_);
  and (_02940_, _02714_, _36036_);
  and (_02941_, _02940_, _35815_);
  not (_02942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor (_02943_, _02940_, _02942_);
  or (_37400_, _02943_, _02941_);
  and (_02944_, _02940_, _35822_);
  not (_02945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor (_02946_, _02940_, _02945_);
  or (_37401_, _02946_, _02944_);
  and (_02947_, _02940_, _35826_);
  not (_02948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor (_02949_, _02940_, _02948_);
  or (_37402_, _02949_, _02947_);
  and (_02950_, _02940_, _35830_);
  not (_02951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  nor (_02952_, _02940_, _02951_);
  or (_37403_, _02952_, _02950_);
  and (_02953_, _02940_, _35834_);
  not (_02954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor (_02955_, _02940_, _02954_);
  or (_37404_, _02955_, _02953_);
  and (_02956_, _02940_, _35838_);
  not (_02957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  nor (_02958_, _02940_, _02957_);
  or (_37405_, _02958_, _02956_);
  and (_02959_, _02940_, _35842_);
  not (_02960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nor (_02961_, _02940_, _02960_);
  or (_37406_, _02961_, _02959_);
  and (_02962_, _02940_, _35846_);
  not (_02963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  nor (_02964_, _02940_, _02963_);
  or (_37407_, _02964_, _02962_);
  and (_02965_, _02714_, _36062_);
  and (_02966_, _02965_, _35815_);
  not (_02967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  nor (_02968_, _02965_, _02967_);
  or (_37408_, _02968_, _02966_);
  and (_02969_, _02965_, _35822_);
  not (_02970_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  nor (_02971_, _02965_, _02970_);
  or (_37409_, _02971_, _02969_);
  and (_02972_, _02965_, _35826_);
  not (_02973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  nor (_02974_, _02965_, _02973_);
  or (_37410_, _02974_, _02972_);
  and (_02975_, _02965_, _35830_);
  not (_02976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor (_02977_, _02965_, _02976_);
  or (_37411_, _02977_, _02975_);
  and (_02978_, _02965_, _35834_);
  not (_02979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  nor (_02980_, _02965_, _02979_);
  or (_37412_, _02980_, _02978_);
  and (_02981_, _02965_, _35838_);
  not (_02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  nor (_02983_, _02965_, _02982_);
  or (_37413_, _02983_, _02981_);
  and (_02984_, _02965_, _35842_);
  not (_02985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  nor (_02986_, _02965_, _02985_);
  or (_37414_, _02986_, _02984_);
  and (_02987_, _02965_, _35846_);
  not (_02988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  nor (_02989_, _02965_, _02988_);
  or (_37415_, _02989_, _02987_);
  and (_02990_, _02714_, _36088_);
  and (_02991_, _02990_, _35815_);
  not (_02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  nor (_02993_, _02990_, _02992_);
  or (_37416_, _02993_, _02991_);
  and (_02994_, _02990_, _35822_);
  not (_02995_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor (_02996_, _02990_, _02995_);
  or (_37417_, _02996_, _02994_);
  and (_02997_, _02990_, _35826_);
  not (_02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  nor (_02999_, _02990_, _02998_);
  or (_37418_, _02999_, _02997_);
  and (_03000_, _02990_, _35830_);
  not (_03001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  nor (_03002_, _02990_, _03001_);
  or (_37419_, _03002_, _03000_);
  and (_03003_, _02990_, _35834_);
  not (_03004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor (_03005_, _02990_, _03004_);
  or (_37420_, _03005_, _03003_);
  and (_03006_, _02990_, _35838_);
  not (_03007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  nor (_03008_, _02990_, _03007_);
  or (_37421_, _03008_, _03006_);
  and (_03009_, _02990_, _35842_);
  not (_03010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor (_03011_, _02990_, _03010_);
  or (_37422_, _03011_, _03009_);
  and (_03012_, _02990_, _35846_);
  not (_03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  nor (_03014_, _02990_, _03013_);
  or (_37423_, _03014_, _03012_);
  and (_03015_, _02714_, _36115_);
  and (_03016_, _03015_, _35815_);
  not (_03017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor (_03018_, _03015_, _03017_);
  or (_37424_, _03018_, _03016_);
  and (_03019_, _03015_, _35822_);
  not (_03020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  nor (_03021_, _03015_, _03020_);
  or (_37425_, _03021_, _03019_);
  and (_03022_, _03015_, _35826_);
  not (_03023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor (_03024_, _03015_, _03023_);
  or (_37426_, _03024_, _03022_);
  and (_03025_, _03015_, _35830_);
  not (_03026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor (_03027_, _03015_, _03026_);
  or (_37427_, _03027_, _03025_);
  and (_03028_, _03015_, _35834_);
  not (_03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  nor (_03030_, _03015_, _03029_);
  or (_37428_, _03030_, _03028_);
  and (_03031_, _03015_, _35838_);
  not (_03032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  nor (_03033_, _03015_, _03032_);
  or (_37429_, _03033_, _03031_);
  and (_03034_, _03015_, _35842_);
  not (_03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  nor (_03036_, _03015_, _03035_);
  or (_37430_, _03036_, _03034_);
  and (_03037_, _03015_, _35846_);
  not (_03038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  nor (_03039_, _03015_, _03038_);
  or (_37431_, _03039_, _03037_);
  and (_03040_, _02714_, _36141_);
  and (_03041_, _03040_, _35815_);
  not (_03042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor (_03043_, _03040_, _03042_);
  or (_37432_, _03043_, _03041_);
  and (_03044_, _03040_, _35822_);
  not (_03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  nor (_03046_, _03040_, _03045_);
  or (_37433_, _03046_, _03044_);
  and (_03047_, _03040_, _35826_);
  not (_03048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor (_03049_, _03040_, _03048_);
  or (_37434_, _03049_, _03047_);
  and (_03050_, _03040_, _35830_);
  not (_03051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  nor (_03052_, _03040_, _03051_);
  or (_37435_, _03052_, _03050_);
  and (_03053_, _03040_, _35834_);
  not (_03054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor (_03055_, _03040_, _03054_);
  or (_37436_, _03055_, _03053_);
  and (_03056_, _03040_, _35838_);
  not (_03057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  nor (_03058_, _03040_, _03057_);
  or (_37437_, _03058_, _03056_);
  and (_03059_, _03040_, _35842_);
  not (_03060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor (_03061_, _03040_, _03060_);
  or (_37438_, _03061_, _03059_);
  and (_03062_, _03040_, _35846_);
  not (_03063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  nor (_03064_, _03040_, _03063_);
  or (_37439_, _03064_, _03062_);
  and (_03065_, _02714_, _36167_);
  and (_03066_, _03065_, _35815_);
  not (_03067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  nor (_03068_, _03065_, _03067_);
  or (_37440_, _03068_, _03066_);
  and (_03069_, _03065_, _35822_);
  not (_03070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor (_03071_, _03065_, _03070_);
  or (_37441_, _03071_, _03069_);
  and (_03072_, _03065_, _35826_);
  not (_03073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  nor (_03074_, _03065_, _03073_);
  or (_37442_, _03074_, _03072_);
  and (_03075_, _03065_, _35830_);
  not (_03076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor (_03077_, _03065_, _03076_);
  or (_37443_, _03077_, _03075_);
  and (_03078_, _03065_, _35834_);
  not (_03079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  nor (_03080_, _03065_, _03079_);
  or (_37444_, _03080_, _03078_);
  and (_03081_, _03065_, _35838_);
  not (_03082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  nor (_03083_, _03065_, _03082_);
  or (_37445_, _03083_, _03081_);
  and (_03084_, _03065_, _35842_);
  not (_03085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  nor (_03086_, _03065_, _03085_);
  or (_37446_, _03086_, _03084_);
  and (_03087_, _03065_, _35846_);
  not (_03088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  nor (_03089_, _03065_, _03088_);
  or (_37447_, _03089_, _03087_);
  and (_03090_, _02714_, _36193_);
  and (_03091_, _03090_, _35815_);
  not (_03092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  nor (_03093_, _03090_, _03092_);
  or (_37448_, _03093_, _03091_);
  and (_03094_, _03090_, _35822_);
  not (_03095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  nor (_03096_, _03090_, _03095_);
  or (_37449_, _03096_, _03094_);
  and (_03097_, _03090_, _35826_);
  not (_03098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  nor (_03099_, _03090_, _03098_);
  or (_37450_, _03099_, _03097_);
  and (_03100_, _03090_, _35830_);
  not (_03101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor (_03102_, _03090_, _03101_);
  or (_37451_, _03102_, _03100_);
  and (_03103_, _03090_, _35834_);
  not (_03104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor (_03105_, _03090_, _03104_);
  or (_37452_, _03105_, _03103_);
  and (_03106_, _03090_, _35838_);
  not (_03107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor (_03108_, _03090_, _03107_);
  or (_37453_, _03108_, _03106_);
  and (_03109_, _03090_, _35842_);
  not (_03110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nor (_03111_, _03090_, _03110_);
  or (_37454_, _03111_, _03109_);
  and (_03112_, _03090_, _35846_);
  not (_03113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  nor (_03114_, _03090_, _03113_);
  or (_37455_, _03114_, _03112_);
  not (_03115_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and (_03116_, _02312_, _36622_);
  and (_03117_, _03116_, _35572_);
  nor (_03118_, _03117_, _03115_);
  and (_03119_, _03117_, _35815_);
  or (_37464_, _03119_, _03118_);
  not (_03120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nor (_03121_, _03117_, _03120_);
  and (_03122_, _03117_, _35822_);
  or (_37465_, _03122_, _03121_);
  not (_03123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nor (_03124_, _03117_, _03123_);
  and (_03125_, _03117_, _35826_);
  or (_37466_, _03125_, _03124_);
  not (_03126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  nor (_03127_, _03117_, _03126_);
  and (_03128_, _03117_, _35830_);
  or (_37467_, _03128_, _03127_);
  not (_03129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  nor (_03130_, _03117_, _03129_);
  and (_03131_, _03117_, _35834_);
  or (_37468_, _03131_, _03130_);
  not (_03132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  nor (_03133_, _03117_, _03132_);
  and (_03134_, _03117_, _35838_);
  or (_37469_, _03134_, _03133_);
  not (_03135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  nor (_03136_, _03117_, _03135_);
  and (_03137_, _03117_, _35842_);
  or (_37470_, _03137_, _03136_);
  not (_03138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  nor (_03139_, _03117_, _03138_);
  and (_03140_, _03117_, _35846_);
  or (_37471_, _03140_, _03139_);
  not (_03141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_03142_, _03116_, _35817_);
  nor (_03143_, _03142_, _03141_);
  and (_03144_, _03142_, _35815_);
  or (_37472_, _03144_, _03143_);
  not (_03145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nor (_03146_, _03142_, _03145_);
  and (_03147_, _03142_, _35822_);
  or (_37473_, _03147_, _03146_);
  not (_03148_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nor (_03149_, _03142_, _03148_);
  and (_03150_, _03142_, _35826_);
  or (_37474_, _03150_, _03149_);
  not (_03151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  nor (_03152_, _03142_, _03151_);
  and (_03153_, _03142_, _35830_);
  or (_37475_, _03153_, _03152_);
  not (_03154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nor (_03155_, _03142_, _03154_);
  and (_03156_, _03142_, _35834_);
  or (_37476_, _03156_, _03155_);
  not (_03157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  nor (_03158_, _03142_, _03157_);
  and (_03159_, _03142_, _35838_);
  or (_37477_, _03159_, _03158_);
  not (_03160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nor (_03161_, _03142_, _03160_);
  and (_03162_, _03142_, _35842_);
  or (_37478_, _03162_, _03161_);
  not (_03163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  nor (_03164_, _03142_, _03163_);
  and (_03165_, _03142_, _35846_);
  or (_37479_, _03165_, _03164_);
  not (_03166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_03167_, _03116_, _35851_);
  nor (_03168_, _03167_, _03166_);
  and (_03169_, _03167_, _35815_);
  or (_37480_, _03169_, _03168_);
  not (_03170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  nor (_03171_, _03167_, _03170_);
  and (_03172_, _03167_, _35822_);
  or (_37481_, _03172_, _03171_);
  not (_03173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  nor (_03174_, _03167_, _03173_);
  and (_03175_, _03167_, _35826_);
  or (_37482_, _03175_, _03174_);
  not (_03176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nor (_03177_, _03167_, _03176_);
  and (_03178_, _03167_, _35830_);
  or (_37483_, _03178_, _03177_);
  not (_03179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  nor (_03180_, _03167_, _03179_);
  and (_03181_, _03167_, _35834_);
  or (_37484_, _03181_, _03180_);
  not (_03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  nor (_03183_, _03167_, _03182_);
  and (_03184_, _03167_, _35838_);
  or (_37485_, _03184_, _03183_);
  not (_03185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  nor (_03186_, _03167_, _03185_);
  and (_03187_, _03167_, _35842_);
  or (_37486_, _03187_, _03186_);
  not (_03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  nor (_03189_, _03167_, _03188_);
  and (_03190_, _03167_, _35846_);
  or (_37487_, _03190_, _03189_);
  not (_03191_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and (_03192_, _03116_, _35878_);
  nor (_03193_, _03192_, _03191_);
  and (_03194_, _03192_, _35815_);
  or (_37488_, _03194_, _03193_);
  not (_03195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  nor (_03196_, _03192_, _03195_);
  and (_03197_, _03192_, _35822_);
  or (_37489_, _03197_, _03196_);
  not (_03198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nor (_03199_, _03192_, _03198_);
  and (_03200_, _03192_, _35826_);
  or (_37490_, _03200_, _03199_);
  not (_03201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nor (_03202_, _03192_, _03201_);
  and (_03203_, _03192_, _35830_);
  or (_37491_, _03203_, _03202_);
  not (_03204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nor (_03205_, _03192_, _03204_);
  and (_03206_, _03192_, _35834_);
  or (_37492_, _03206_, _03205_);
  not (_03207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  nor (_03208_, _03192_, _03207_);
  and (_03209_, _03192_, _35838_);
  or (_37493_, _03209_, _03208_);
  not (_03210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nor (_03211_, _03192_, _03210_);
  and (_03212_, _03192_, _35842_);
  or (_37494_, _03212_, _03211_);
  not (_03213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  nor (_03214_, _03192_, _03213_);
  and (_03215_, _03192_, _35846_);
  or (_37495_, _03215_, _03214_);
  not (_03216_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_03217_, _03116_, _35905_);
  nor (_03218_, _03217_, _03216_);
  and (_03219_, _03217_, _35815_);
  or (_37496_, _03219_, _03218_);
  not (_03220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nor (_03221_, _03217_, _03220_);
  and (_03222_, _03217_, _35822_);
  or (_37497_, _03222_, _03221_);
  not (_03223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  nor (_03224_, _03217_, _03223_);
  and (_03225_, _03217_, _35826_);
  or (_37498_, _03225_, _03224_);
  not (_03226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  nor (_03227_, _03217_, _03226_);
  and (_03228_, _03217_, _35830_);
  or (_37499_, _03228_, _03227_);
  not (_03229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  nor (_03230_, _03217_, _03229_);
  and (_03231_, _03217_, _35834_);
  or (_37500_, _03231_, _03230_);
  not (_03232_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nor (_03233_, _03217_, _03232_);
  and (_03234_, _03217_, _35838_);
  or (_37501_, _03234_, _03233_);
  not (_03235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  nor (_03236_, _03217_, _03235_);
  and (_03237_, _03217_, _35842_);
  or (_37502_, _03237_, _03236_);
  not (_03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  nor (_03239_, _03217_, _03238_);
  and (_03240_, _03217_, _35846_);
  or (_37503_, _03240_, _03239_);
  not (_03241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_03242_, _03116_, _35931_);
  nor (_03243_, _03242_, _03241_);
  and (_03244_, _03242_, _35815_);
  or (_37504_, _03244_, _03243_);
  not (_03245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  nor (_03246_, _03242_, _03245_);
  and (_03247_, _03242_, _35822_);
  or (_37505_, _03247_, _03246_);
  not (_03248_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nor (_03249_, _03242_, _03248_);
  and (_03250_, _03242_, _35826_);
  or (_37506_, _03250_, _03249_);
  not (_03251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nor (_03252_, _03242_, _03251_);
  and (_03253_, _03242_, _35830_);
  or (_37507_, _03253_, _03252_);
  not (_03254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  nor (_03255_, _03242_, _03254_);
  and (_03256_, _03242_, _35834_);
  or (_37508_, _03256_, _03255_);
  not (_03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  nor (_03258_, _03242_, _03257_);
  and (_03259_, _03242_, _35838_);
  or (_37509_, _03259_, _03258_);
  not (_03260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nor (_03261_, _03242_, _03260_);
  and (_03262_, _03242_, _35842_);
  or (_37510_, _03262_, _03261_);
  not (_03263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  nor (_03264_, _03242_, _03263_);
  and (_03265_, _03242_, _35846_);
  or (_37511_, _03265_, _03264_);
  not (_03266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_03267_, _03116_, _35957_);
  nor (_03268_, _03267_, _03266_);
  and (_03269_, _03267_, _35815_);
  or (_37512_, _03269_, _03268_);
  not (_03270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nor (_03271_, _03267_, _03270_);
  and (_03272_, _03267_, _35822_);
  or (_37513_, _03272_, _03271_);
  not (_03273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  nor (_03274_, _03267_, _03273_);
  and (_03275_, _03267_, _35826_);
  or (_37514_, _03275_, _03274_);
  not (_03276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  nor (_03277_, _03267_, _03276_);
  and (_03278_, _03267_, _35830_);
  or (_37515_, _03278_, _03277_);
  not (_03279_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nor (_03280_, _03267_, _03279_);
  and (_03281_, _03267_, _35834_);
  or (_37516_, _03281_, _03280_);
  not (_03282_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  nor (_03283_, _03267_, _03282_);
  and (_03284_, _03267_, _35838_);
  or (_37517_, _03284_, _03283_);
  not (_03285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  nor (_03286_, _03267_, _03285_);
  and (_03287_, _03267_, _35842_);
  or (_37518_, _03287_, _03286_);
  not (_03288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  nor (_03289_, _03267_, _03288_);
  and (_03290_, _03267_, _35846_);
  or (_37519_, _03290_, _03289_);
  not (_03291_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_03292_, _03116_, _35983_);
  nor (_03293_, _03292_, _03291_);
  and (_03294_, _03292_, _35815_);
  or (_37520_, _03294_, _03293_);
  not (_03295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nor (_03296_, _03292_, _03295_);
  and (_03297_, _03292_, _35822_);
  or (_37521_, _03297_, _03296_);
  not (_03298_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  nor (_03299_, _03292_, _03298_);
  and (_03300_, _03292_, _35826_);
  or (_37522_, _03300_, _03299_);
  not (_03301_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nor (_03302_, _03292_, _03301_);
  and (_03303_, _03292_, _35830_);
  or (_37523_, _03303_, _03302_);
  not (_03304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  nor (_03305_, _03292_, _03304_);
  and (_03306_, _03292_, _35834_);
  or (_37524_, _03306_, _03305_);
  not (_03307_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  nor (_03308_, _03292_, _03307_);
  and (_03309_, _03292_, _35838_);
  or (_37525_, _03309_, _03308_);
  not (_03310_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  nor (_03311_, _03292_, _03310_);
  and (_03312_, _03292_, _35842_);
  or (_37526_, _03312_, _03311_);
  not (_03313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  nor (_03314_, _03292_, _03313_);
  and (_03315_, _03292_, _35846_);
  or (_37527_, _03315_, _03314_);
  not (_03316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_03317_, _03116_, _36010_);
  nor (_03318_, _03317_, _03316_);
  and (_03319_, _03317_, _35815_);
  or (_37528_, _03319_, _03318_);
  not (_03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  nor (_03321_, _03317_, _03320_);
  and (_03322_, _03317_, _35822_);
  or (_37529_, _03322_, _03321_);
  not (_03323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nor (_03324_, _03317_, _03323_);
  and (_03325_, _03317_, _35826_);
  or (_37530_, _03325_, _03324_);
  not (_03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  nor (_03327_, _03317_, _03326_);
  and (_03328_, _03317_, _35830_);
  or (_37531_, _03328_, _03327_);
  not (_03329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nor (_03330_, _03317_, _03329_);
  and (_03331_, _03317_, _35834_);
  or (_37532_, _03331_, _03330_);
  not (_03332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  nor (_03333_, _03317_, _03332_);
  and (_03334_, _03317_, _35838_);
  or (_37533_, _03334_, _03333_);
  not (_03335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nor (_03336_, _03317_, _03335_);
  and (_03337_, _03317_, _35842_);
  or (_37534_, _03337_, _03336_);
  not (_03338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  nor (_03339_, _03317_, _03338_);
  and (_03340_, _03317_, _35846_);
  or (_37535_, _03340_, _03339_);
  not (_03341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and (_03342_, _03116_, _36036_);
  nor (_03343_, _03342_, _03341_);
  and (_03344_, _03342_, _35815_);
  or (_37536_, _03344_, _03343_);
  not (_03345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nor (_03346_, _03342_, _03345_);
  and (_03347_, _03342_, _35822_);
  or (_37537_, _03347_, _03346_);
  not (_03348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nor (_03349_, _03342_, _03348_);
  and (_03350_, _03342_, _35826_);
  or (_37538_, _03350_, _03349_);
  not (_03351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  nor (_03352_, _03342_, _03351_);
  and (_03353_, _03342_, _35830_);
  or (_37539_, _03353_, _03352_);
  not (_03354_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nor (_03355_, _03342_, _03354_);
  and (_03356_, _03342_, _35834_);
  or (_37540_, _03356_, _03355_);
  not (_03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  nor (_03358_, _03342_, _03357_);
  and (_03359_, _03342_, _35838_);
  or (_37541_, _03359_, _03358_);
  not (_03360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nor (_03361_, _03342_, _03360_);
  and (_03362_, _03342_, _35842_);
  or (_37542_, _03362_, _03361_);
  not (_03363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  nor (_03364_, _03342_, _03363_);
  and (_03365_, _03342_, _35846_);
  or (_37543_, _03365_, _03364_);
  not (_03366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_03367_, _03116_, _36062_);
  nor (_03368_, _03367_, _03366_);
  and (_03369_, _03367_, _35815_);
  or (_37552_, _03369_, _03368_);
  not (_03370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  nor (_03371_, _03367_, _03370_);
  and (_03372_, _03367_, _35822_);
  or (_37553_, _03372_, _03371_);
  not (_03373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  nor (_03374_, _03367_, _03373_);
  and (_03375_, _03367_, _35826_);
  or (_37554_, _03375_, _03374_);
  not (_03376_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor (_03377_, _03367_, _03376_);
  and (_03378_, _03367_, _35830_);
  or (_37555_, _03378_, _03377_);
  not (_03379_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  nor (_03380_, _03367_, _03379_);
  and (_03381_, _03367_, _35834_);
  or (_37556_, _03381_, _03380_);
  not (_03382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  nor (_03383_, _03367_, _03382_);
  and (_03384_, _03367_, _35838_);
  or (_37557_, _03384_, _03383_);
  not (_03385_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  nor (_03386_, _03367_, _03385_);
  and (_03387_, _03367_, _35842_);
  or (_37558_, _03387_, _03386_);
  not (_03388_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nor (_03389_, _03367_, _03388_);
  and (_03390_, _03367_, _35846_);
  or (_37559_, _03390_, _03389_);
  not (_03391_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_03392_, _03116_, _36088_);
  nor (_03393_, _03392_, _03391_);
  and (_03394_, _03392_, _35815_);
  or (_37560_, _03394_, _03393_);
  not (_03395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  nor (_03396_, _03392_, _03395_);
  and (_03397_, _03392_, _35822_);
  or (_37561_, _03397_, _03396_);
  not (_03398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  nor (_03399_, _03392_, _03398_);
  and (_03400_, _03392_, _35826_);
  or (_37562_, _03400_, _03399_);
  not (_03401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  nor (_03402_, _03392_, _03401_);
  and (_03403_, _03392_, _35830_);
  or (_37563_, _03403_, _03402_);
  not (_03404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor (_03405_, _03392_, _03404_);
  and (_03406_, _03392_, _35834_);
  or (_37564_, _03406_, _03405_);
  not (_03407_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  nor (_03408_, _03392_, _03407_);
  and (_03409_, _03392_, _35838_);
  or (_37565_, _03409_, _03408_);
  not (_03410_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  nor (_03411_, _03392_, _03410_);
  and (_03412_, _03392_, _35842_);
  or (_37566_, _03412_, _03411_);
  not (_03413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  nor (_03414_, _03392_, _03413_);
  and (_03415_, _03392_, _35846_);
  or (_37567_, _03415_, _03414_);
  not (_03416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_03417_, _03116_, _36115_);
  nor (_03418_, _03417_, _03416_);
  and (_03419_, _03417_, _35815_);
  or (_37568_, _03419_, _03418_);
  not (_03420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nor (_03421_, _03417_, _03420_);
  and (_03422_, _03417_, _35822_);
  or (_37569_, _03422_, _03421_);
  not (_03423_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nor (_03424_, _03417_, _03423_);
  and (_03425_, _03417_, _35826_);
  or (_37570_, _03425_, _03424_);
  not (_03426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nor (_03427_, _03417_, _03426_);
  and (_03428_, _03417_, _35830_);
  or (_37571_, _03428_, _03427_);
  not (_03429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  nor (_03430_, _03417_, _03429_);
  and (_03431_, _03417_, _35834_);
  or (_37572_, _03431_, _03430_);
  not (_03432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  nor (_03433_, _03417_, _03432_);
  and (_03434_, _03417_, _35838_);
  or (_37573_, _03434_, _03433_);
  not (_03435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nor (_03436_, _03417_, _03435_);
  and (_03437_, _03417_, _35842_);
  or (_37574_, _03437_, _03436_);
  not (_03438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  nor (_03439_, _03417_, _03438_);
  and (_03440_, _03417_, _35846_);
  or (_37575_, _03440_, _03439_);
  not (_03441_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_03442_, _03116_, _36141_);
  nor (_03443_, _03442_, _03441_);
  and (_03444_, _03442_, _35815_);
  or (_37576_, _03444_, _03443_);
  not (_03445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  nor (_03446_, _03442_, _03445_);
  and (_03447_, _03442_, _35822_);
  or (_37577_, _03447_, _03446_);
  not (_03448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nor (_03449_, _03442_, _03448_);
  and (_03450_, _03442_, _35826_);
  or (_37578_, _03450_, _03449_);
  not (_03451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nor (_03452_, _03442_, _03451_);
  and (_03453_, _03442_, _35830_);
  or (_37579_, _03453_, _03452_);
  not (_03454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  nor (_03455_, _03442_, _03454_);
  and (_03456_, _03442_, _35834_);
  or (_37580_, _03456_, _03455_);
  not (_03457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  nor (_03458_, _03442_, _03457_);
  and (_03459_, _03442_, _35838_);
  or (_37581_, _03459_, _03458_);
  not (_03460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nor (_03461_, _03442_, _03460_);
  and (_03462_, _03442_, _35842_);
  or (_37582_, _03462_, _03461_);
  not (_03463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  nor (_03464_, _03442_, _03463_);
  and (_03465_, _03442_, _35846_);
  or (_37583_, _03465_, _03464_);
  not (_03466_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_03467_, _03116_, _36167_);
  nor (_03468_, _03467_, _03466_);
  and (_03469_, _03467_, _35815_);
  or (_37584_, _03469_, _03468_);
  not (_03470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor (_03471_, _03467_, _03470_);
  and (_03472_, _03467_, _35822_);
  or (_37585_, _03472_, _03471_);
  not (_03473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  nor (_03474_, _03467_, _03473_);
  and (_03475_, _03467_, _35826_);
  or (_37586_, _03475_, _03474_);
  not (_03476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  nor (_03477_, _03467_, _03476_);
  and (_03478_, _03467_, _35830_);
  or (_37587_, _03478_, _03477_);
  not (_03479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor (_03480_, _03467_, _03479_);
  and (_03481_, _03467_, _35834_);
  or (_37588_, _03481_, _03480_);
  not (_03482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  nor (_03483_, _03467_, _03482_);
  and (_03484_, _03467_, _35838_);
  or (_37589_, _03484_, _03483_);
  not (_03485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  nor (_03486_, _03467_, _03485_);
  and (_03487_, _03467_, _35842_);
  or (_37590_, _03487_, _03486_);
  not (_03488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  nor (_03489_, _03467_, _03488_);
  and (_03490_, _03467_, _35846_);
  or (_37591_, _03490_, _03489_);
  not (_03491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_03492_, _03116_, _36193_);
  nor (_03493_, _03492_, _03491_);
  and (_03494_, _03492_, _35815_);
  or (_37592_, _03494_, _03493_);
  not (_03495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor (_03496_, _03492_, _03495_);
  and (_03497_, _03492_, _35822_);
  or (_37593_, _03497_, _03496_);
  not (_03498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  nor (_03499_, _03492_, _03498_);
  and (_03500_, _03492_, _35826_);
  or (_37594_, _03500_, _03499_);
  not (_03501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nor (_03502_, _03492_, _03501_);
  and (_03503_, _03492_, _35830_);
  or (_37595_, _03503_, _03502_);
  not (_03504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor (_03505_, _03492_, _03504_);
  and (_03506_, _03492_, _35834_);
  or (_37596_, _03506_, _03505_);
  not (_03507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nor (_03508_, _03492_, _03507_);
  and (_03509_, _03492_, _35838_);
  or (_37597_, _03509_, _03508_);
  not (_03510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor (_03511_, _03492_, _03510_);
  and (_03512_, _03492_, _35842_);
  or (_37598_, _03512_, _03511_);
  not (_03513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  nor (_03514_, _03492_, _03513_);
  and (_03515_, _03492_, _35846_);
  or (_37599_, _03515_, _03514_);
  and (_03516_, _00304_, _33632_);
  and (_03517_, _03516_, _35572_);
  and (_03518_, _03517_, _35815_);
  not (_03519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nor (_03520_, _03517_, _03519_);
  or (_37600_, _03520_, _03518_);
  and (_03521_, _03517_, _35822_);
  not (_03522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nor (_03523_, _03517_, _03522_);
  or (_37601_, _03523_, _03521_);
  and (_03524_, _03517_, _35826_);
  not (_03525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nor (_03526_, _03517_, _03525_);
  or (_37602_, _03526_, _03524_);
  and (_03527_, _03517_, _35830_);
  not (_03528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  nor (_03529_, _03517_, _03528_);
  or (_37603_, _03529_, _03527_);
  and (_03530_, _03517_, _35834_);
  not (_03531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  nor (_03532_, _03517_, _03531_);
  or (_37604_, _03532_, _03530_);
  and (_03533_, _03517_, _35838_);
  not (_03534_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  nor (_03535_, _03517_, _03534_);
  or (_37605_, _03535_, _03533_);
  and (_03536_, _03517_, _35842_);
  not (_03537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  nor (_03538_, _03517_, _03537_);
  or (_37606_, _03538_, _03536_);
  and (_03539_, _03517_, _35846_);
  not (_03540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  nor (_03541_, _03517_, _03540_);
  or (_37607_, _03541_, _03539_);
  and (_03542_, _03516_, _35817_);
  and (_03543_, _03542_, _35815_);
  not (_03544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nor (_03545_, _03542_, _03544_);
  or (_37608_, _03545_, _03543_);
  and (_03546_, _03542_, _35822_);
  not (_03547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  nor (_03548_, _03542_, _03547_);
  or (_37609_, _03548_, _03546_);
  and (_03549_, _03542_, _35826_);
  not (_03550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  nor (_03551_, _03542_, _03550_);
  or (_37610_, _03551_, _03549_);
  and (_03552_, _03542_, _35830_);
  not (_03553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  nor (_03554_, _03542_, _03553_);
  or (_37611_, _03554_, _03552_);
  and (_03555_, _03542_, _35834_);
  not (_03556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nor (_03557_, _03542_, _03556_);
  or (_37612_, _03557_, _03555_);
  and (_03558_, _03542_, _35838_);
  not (_03559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  nor (_03560_, _03542_, _03559_);
  or (_37613_, _03560_, _03558_);
  and (_03561_, _03542_, _35842_);
  not (_03562_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  nor (_03563_, _03542_, _03562_);
  or (_37614_, _03563_, _03561_);
  and (_03564_, _03542_, _35846_);
  not (_03565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  nor (_03566_, _03542_, _03565_);
  or (_37615_, _03566_, _03564_);
  and (_03567_, _03516_, _35851_);
  and (_03568_, _03567_, _35815_);
  not (_03569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  nor (_03570_, _03567_, _03569_);
  or (_37616_, _03570_, _03568_);
  and (_03571_, _03567_, _35822_);
  not (_03572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nor (_03573_, _03567_, _03572_);
  or (_37617_, _03573_, _03571_);
  and (_03574_, _03567_, _35826_);
  not (_03575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nor (_03576_, _03567_, _03575_);
  or (_37618_, _03576_, _03574_);
  and (_03577_, _03567_, _35830_);
  not (_03578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nor (_03579_, _03567_, _03578_);
  or (_37619_, _03579_, _03577_);
  and (_03580_, _03567_, _35834_);
  not (_03581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  nor (_03582_, _03567_, _03581_);
  or (_37620_, _03582_, _03580_);
  and (_03583_, _03567_, _35838_);
  not (_03584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  nor (_03585_, _03567_, _03584_);
  or (_37621_, _03585_, _03583_);
  and (_03586_, _03567_, _35842_);
  not (_03587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nor (_03588_, _03567_, _03587_);
  or (_37622_, _03588_, _03586_);
  and (_03589_, _03567_, _35846_);
  not (_03590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  nor (_03591_, _03567_, _03590_);
  or (_37623_, _03591_, _03589_);
  and (_03592_, _03516_, _35878_);
  and (_03593_, _03592_, _35815_);
  not (_03594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  nor (_03595_, _03592_, _03594_);
  or (_37624_, _03595_, _03593_);
  and (_03596_, _03592_, _35822_);
  not (_03597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nor (_03598_, _03592_, _03597_);
  or (_37625_, _03598_, _03596_);
  and (_03599_, _03592_, _35826_);
  not (_03600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nor (_03601_, _03592_, _03600_);
  or (_37626_, _03601_, _03599_);
  and (_03602_, _03592_, _35830_);
  not (_03603_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  nor (_03604_, _03592_, _03603_);
  or (_37627_, _03604_, _03602_);
  and (_03605_, _03592_, _35834_);
  not (_03606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nor (_03607_, _03592_, _03606_);
  or (_37628_, _03607_, _03605_);
  and (_03608_, _03592_, _35838_);
  not (_03609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  nor (_03610_, _03592_, _03609_);
  or (_37629_, _03610_, _03608_);
  and (_03611_, _03592_, _35842_);
  not (_03612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  nor (_03613_, _03592_, _03612_);
  or (_37630_, _03613_, _03611_);
  and (_03614_, _03592_, _35846_);
  not (_03615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  nor (_03616_, _03592_, _03615_);
  or (_37631_, _03616_, _03614_);
  and (_03617_, _03516_, _35905_);
  and (_03618_, _03617_, _35815_);
  not (_03619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nor (_03620_, _03617_, _03619_);
  or (_37640_, _03620_, _03618_);
  and (_03621_, _03617_, _35822_);
  not (_03622_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  nor (_03623_, _03617_, _03622_);
  or (_37641_, _03623_, _03621_);
  and (_03624_, _03617_, _35826_);
  not (_03625_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  nor (_03626_, _03617_, _03625_);
  or (_37642_, _03626_, _03624_);
  and (_03627_, _03617_, _35830_);
  not (_03628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nor (_03629_, _03617_, _03628_);
  or (_37643_, _03629_, _03627_);
  and (_03630_, _03617_, _35834_);
  not (_03631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  nor (_03632_, _03617_, _03631_);
  or (_37644_, _03632_, _03630_);
  and (_03633_, _03617_, _35838_);
  not (_03634_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  nor (_03635_, _03617_, _03634_);
  or (_37645_, _03635_, _03633_);
  and (_03636_, _03617_, _35842_);
  not (_03637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nor (_03638_, _03617_, _03637_);
  or (_37646_, _03638_, _03636_);
  and (_03639_, _03617_, _35846_);
  not (_03640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  nor (_03641_, _03617_, _03640_);
  or (_37647_, _03641_, _03639_);
  and (_03642_, _03516_, _35931_);
  and (_03643_, _03642_, _35815_);
  not (_03644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  nor (_03645_, _03642_, _03644_);
  or (_37648_, _03645_, _03643_);
  and (_03646_, _03642_, _35822_);
  not (_03647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nor (_03648_, _03642_, _03647_);
  or (_37649_, _03648_, _03646_);
  and (_03649_, _03642_, _35826_);
  not (_03650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  nor (_03651_, _03642_, _03650_);
  or (_37650_, _03651_, _03649_);
  and (_03652_, _03642_, _35830_);
  not (_03653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  nor (_03654_, _03642_, _03653_);
  or (_37651_, _03654_, _03652_);
  and (_03655_, _03642_, _35834_);
  not (_03656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nor (_03657_, _03642_, _03656_);
  or (_37652_, _03657_, _03655_);
  and (_03658_, _03642_, _35838_);
  not (_03659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  nor (_03660_, _03642_, _03659_);
  or (_37653_, _03660_, _03658_);
  and (_03661_, _03642_, _35842_);
  not (_03662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nor (_03663_, _03642_, _03662_);
  or (_37654_, _03663_, _03661_);
  and (_03664_, _03642_, _35846_);
  not (_03665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  nor (_03666_, _03642_, _03665_);
  or (_37655_, _03666_, _03664_);
  and (_03667_, _03516_, _35957_);
  and (_03668_, _03667_, _35815_);
  not (_03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nor (_03670_, _03667_, _03669_);
  or (_37656_, _03670_, _03668_);
  and (_03671_, _03667_, _35822_);
  not (_03672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  nor (_03673_, _03667_, _03672_);
  or (_37657_, _03673_, _03671_);
  and (_03674_, _03667_, _35826_);
  not (_03675_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nor (_03676_, _03667_, _03675_);
  or (_37658_, _03676_, _03674_);
  and (_03677_, _03667_, _35830_);
  not (_03678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nor (_03679_, _03667_, _03678_);
  or (_37659_, _03679_, _03677_);
  and (_03680_, _03667_, _35834_);
  not (_03681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  nor (_03682_, _03667_, _03681_);
  or (_37660_, _03682_, _03680_);
  and (_03683_, _03667_, _35838_);
  not (_03684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  nor (_03685_, _03667_, _03684_);
  or (_37661_, _03685_, _03683_);
  and (_03686_, _03667_, _35842_);
  not (_03687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  nor (_03688_, _03667_, _03687_);
  or (_37662_, _03688_, _03686_);
  and (_03689_, _03667_, _35846_);
  not (_03690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  nor (_03691_, _03667_, _03690_);
  or (_37663_, _03691_, _03689_);
  and (_03692_, _03516_, _35983_);
  and (_03693_, _03692_, _35815_);
  not (_03694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  nor (_03695_, _03692_, _03694_);
  or (_37664_, _03695_, _03693_);
  and (_03696_, _03692_, _35822_);
  not (_03697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nor (_03698_, _03692_, _03697_);
  or (_37665_, _03698_, _03696_);
  and (_03699_, _03692_, _35826_);
  not (_03700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nor (_03701_, _03692_, _03700_);
  or (_37666_, _03701_, _03699_);
  and (_03702_, _03692_, _35830_);
  not (_03703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  nor (_03704_, _03692_, _03703_);
  or (_37667_, _03704_, _03702_);
  and (_03705_, _03692_, _35834_);
  not (_03706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  nor (_03707_, _03692_, _03706_);
  or (_37668_, _03707_, _03705_);
  and (_03708_, _03692_, _35838_);
  not (_03709_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  nor (_03710_, _03692_, _03709_);
  or (_37669_, _03710_, _03708_);
  and (_03711_, _03692_, _35842_);
  not (_03712_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  nor (_03713_, _03692_, _03712_);
  or (_37670_, _03713_, _03711_);
  and (_03714_, _03692_, _35846_);
  not (_03715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  nor (_03716_, _03692_, _03715_);
  or (_37671_, _03716_, _03714_);
  and (_03717_, _03516_, _36010_);
  and (_03718_, _03717_, _35815_);
  not (_03719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor (_03720_, _03717_, _03719_);
  or (_37672_, _03720_, _03718_);
  and (_03721_, _03717_, _35822_);
  not (_03722_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  nor (_03723_, _03717_, _03722_);
  or (_37673_, _03723_, _03721_);
  and (_03724_, _03717_, _35826_);
  not (_03725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  nor (_03726_, _03717_, _03725_);
  or (_37674_, _03726_, _03724_);
  and (_03727_, _03717_, _35830_);
  not (_03728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor (_03729_, _03717_, _03728_);
  or (_37675_, _03729_, _03727_);
  and (_03730_, _03717_, _35834_);
  not (_03731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nor (_03732_, _03717_, _03731_);
  or (_37676_, _03732_, _03730_);
  and (_03733_, _03717_, _35838_);
  not (_03734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  nor (_03735_, _03717_, _03734_);
  or (_37677_, _03735_, _03733_);
  and (_03736_, _03717_, _35842_);
  not (_03737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor (_03738_, _03717_, _03737_);
  or (_37678_, _03738_, _03736_);
  and (_03739_, _03717_, _35846_);
  not (_03740_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  nor (_03741_, _03717_, _03740_);
  or (_37679_, _03741_, _03739_);
  and (_03742_, _03516_, _36036_);
  and (_03743_, _03742_, _35815_);
  not (_03744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor (_03745_, _03742_, _03744_);
  or (_37680_, _03745_, _03743_);
  and (_03746_, _03742_, _35822_);
  not (_03747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  nor (_03748_, _03742_, _03747_);
  or (_37681_, _03748_, _03746_);
  and (_03749_, _03742_, _35826_);
  not (_03750_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  nor (_03751_, _03742_, _03750_);
  or (_37682_, _03751_, _03749_);
  and (_03752_, _03742_, _35830_);
  not (_03753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nor (_03754_, _03742_, _03753_);
  or (_37683_, _03754_, _03752_);
  and (_03755_, _03742_, _35834_);
  not (_03756_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  nor (_03757_, _03742_, _03756_);
  or (_37684_, _03757_, _03755_);
  and (_03758_, _03742_, _35838_);
  not (_03759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  nor (_03760_, _03742_, _03759_);
  or (_37685_, _03760_, _03758_);
  and (_03761_, _03742_, _35842_);
  not (_03762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  nor (_03763_, _03742_, _03762_);
  or (_37686_, _03763_, _03761_);
  and (_03764_, _03742_, _35846_);
  not (_03765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  nor (_03766_, _03742_, _03765_);
  or (_37687_, _03766_, _03764_);
  and (_03767_, _03516_, _36062_);
  and (_03768_, _03767_, _35815_);
  not (_03769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  nor (_03770_, _03767_, _03769_);
  or (_37688_, _03770_, _03768_);
  and (_03771_, _03767_, _35822_);
  not (_03772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor (_03773_, _03767_, _03772_);
  or (_37689_, _03773_, _03771_);
  and (_03774_, _03767_, _35826_);
  not (_03775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor (_03776_, _03767_, _03775_);
  or (_37690_, _03776_, _03774_);
  and (_03777_, _03767_, _35830_);
  not (_03778_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  nor (_03779_, _03767_, _03778_);
  or (_37691_, _03779_, _03777_);
  and (_03780_, _03767_, _35834_);
  not (_03781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor (_03782_, _03767_, _03781_);
  or (_37692_, _03782_, _03780_);
  and (_03783_, _03767_, _35838_);
  not (_03784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  nor (_03785_, _03767_, _03784_);
  or (_37693_, _03785_, _03783_);
  and (_03786_, _03767_, _35842_);
  not (_03787_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor (_03788_, _03767_, _03787_);
  or (_37694_, _03788_, _03786_);
  and (_03789_, _03767_, _35846_);
  not (_03790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  nor (_03791_, _03767_, _03790_);
  or (_37695_, _03791_, _03789_);
  and (_03792_, _03516_, _36088_);
  and (_03793_, _03792_, _35815_);
  not (_03794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  nor (_03795_, _03792_, _03794_);
  or (_37696_, _03795_, _03793_);
  and (_03796_, _03792_, _35822_);
  not (_03797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  nor (_03798_, _03792_, _03797_);
  or (_37697_, _03798_, _03796_);
  and (_03799_, _03792_, _35826_);
  not (_03800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  nor (_03801_, _03792_, _03800_);
  or (_37698_, _03801_, _03799_);
  and (_03802_, _03792_, _35830_);
  not (_03803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor (_03804_, _03792_, _03803_);
  or (_37699_, _03804_, _03802_);
  and (_03805_, _03792_, _35834_);
  not (_03806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  nor (_03807_, _03792_, _03806_);
  or (_37700_, _03807_, _03805_);
  and (_03808_, _03792_, _35838_);
  not (_03809_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  nor (_03810_, _03792_, _03809_);
  or (_37701_, _03810_, _03808_);
  and (_03811_, _03792_, _35842_);
  not (_03812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor (_03813_, _03792_, _03812_);
  or (_37702_, _03813_, _03811_);
  and (_03814_, _03792_, _35846_);
  not (_03815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  nor (_03816_, _03792_, _03815_);
  or (_37703_, _03816_, _03814_);
  and (_03817_, _03516_, _36115_);
  and (_03818_, _03817_, _35815_);
  not (_03819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor (_03820_, _03817_, _03819_);
  or (_37704_, _03820_, _03818_);
  and (_03821_, _03817_, _35822_);
  not (_03822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor (_03823_, _03817_, _03822_);
  or (_37705_, _03823_, _03821_);
  and (_03824_, _03817_, _35826_);
  not (_03825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nor (_03826_, _03817_, _03825_);
  or (_37706_, _03826_, _03824_);
  and (_03827_, _03817_, _35830_);
  not (_03828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  nor (_03829_, _03817_, _03828_);
  or (_37707_, _03829_, _03827_);
  and (_03830_, _03817_, _35834_);
  not (_03831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor (_03832_, _03817_, _03831_);
  or (_37708_, _03832_, _03830_);
  and (_03833_, _03817_, _35838_);
  not (_03834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  nor (_03835_, _03817_, _03834_);
  or (_37709_, _03835_, _03833_);
  and (_03836_, _03817_, _35842_);
  not (_03837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  nor (_03838_, _03817_, _03837_);
  or (_37710_, _03838_, _03836_);
  and (_03839_, _03817_, _35846_);
  not (_03840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  nor (_03841_, _03817_, _03840_);
  or (_37711_, _03841_, _03839_);
  and (_03842_, _03516_, _36141_);
  and (_03843_, _03842_, _35815_);
  not (_03844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor (_03845_, _03842_, _03844_);
  or (_37712_, _03845_, _03843_);
  and (_03846_, _03842_, _35822_);
  not (_03847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  nor (_03848_, _03842_, _03847_);
  or (_37713_, _03848_, _03846_);
  and (_03849_, _03842_, _35826_);
  not (_03850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor (_03851_, _03842_, _03850_);
  or (_37714_, _03851_, _03849_);
  and (_03852_, _03842_, _35830_);
  not (_03853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  nor (_03854_, _03842_, _03853_);
  or (_37715_, _03854_, _03852_);
  and (_03855_, _03842_, _35834_);
  not (_03856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor (_03857_, _03842_, _03856_);
  or (_37716_, _03857_, _03855_);
  and (_03858_, _03842_, _35838_);
  not (_03859_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  nor (_03860_, _03842_, _03859_);
  or (_37717_, _03860_, _03858_);
  and (_03861_, _03842_, _35842_);
  not (_03862_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  nor (_03863_, _03842_, _03862_);
  or (_37718_, _03863_, _03861_);
  and (_03864_, _03842_, _35846_);
  not (_03865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  nor (_03866_, _03842_, _03865_);
  or (_37719_, _03866_, _03864_);
  and (_03867_, _03516_, _36167_);
  and (_03868_, _03867_, _35815_);
  not (_03869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  nor (_03870_, _03867_, _03869_);
  or (_37728_, _03870_, _03868_);
  and (_03871_, _03867_, _35822_);
  not (_03872_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nor (_03873_, _03867_, _03872_);
  or (_37729_, _03873_, _03871_);
  and (_03874_, _03867_, _35826_);
  not (_03875_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  nor (_03876_, _03867_, _03875_);
  or (_37730_, _03876_, _03874_);
  and (_03877_, _03867_, _35830_);
  not (_03878_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor (_03879_, _03867_, _03878_);
  or (_37731_, _03879_, _03877_);
  and (_03880_, _03867_, _35834_);
  not (_03881_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  nor (_03882_, _03867_, _03881_);
  or (_37732_, _03882_, _03880_);
  and (_03883_, _03867_, _35838_);
  not (_03884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  nor (_03885_, _03867_, _03884_);
  or (_37733_, _03885_, _03883_);
  and (_03886_, _03867_, _35842_);
  not (_03887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor (_03888_, _03867_, _03887_);
  or (_37734_, _03888_, _03886_);
  and (_03889_, _03867_, _35846_);
  not (_03890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  nor (_03891_, _03867_, _03890_);
  or (_37735_, _03891_, _03889_);
  and (_03892_, _03516_, _36193_);
  and (_03893_, _03892_, _35815_);
  not (_03894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  nor (_03895_, _03892_, _03894_);
  or (_37736_, _03895_, _03893_);
  and (_03896_, _03892_, _35822_);
  not (_03897_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor (_03898_, _03892_, _03897_);
  or (_37737_, _03898_, _03896_);
  and (_03899_, _03892_, _35826_);
  not (_03900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  nor (_03901_, _03892_, _03900_);
  or (_37738_, _03901_, _03899_);
  and (_03902_, _03892_, _35830_);
  not (_03903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  nor (_03904_, _03892_, _03903_);
  or (_37739_, _03904_, _03902_);
  and (_03905_, _03892_, _35834_);
  not (_03906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor (_03907_, _03892_, _03906_);
  or (_37740_, _03907_, _03905_);
  and (_03908_, _03892_, _35838_);
  not (_03909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  nor (_03910_, _03892_, _03909_);
  or (_37741_, _03910_, _03908_);
  and (_03911_, _03892_, _35842_);
  not (_03912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nor (_03913_, _03892_, _03912_);
  or (_37742_, _03913_, _03911_);
  and (_03914_, _03892_, _35846_);
  not (_03915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  nor (_03916_, _03892_, _03915_);
  or (_37743_, _03916_, _03914_);
  and (_03917_, _34784_, _34231_);
  and (_03918_, _03917_, _35575_);
  and (_03919_, _03918_, _35572_);
  and (_03920_, _03919_, _35815_);
  not (_03921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nor (_03922_, _03919_, _03921_);
  or (_37744_, _03922_, _03920_);
  and (_03923_, _03919_, _35822_);
  not (_03924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  nor (_03925_, _03919_, _03924_);
  or (_37745_, _03925_, _03923_);
  and (_03926_, _03919_, _35826_);
  not (_03927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nor (_03928_, _03919_, _03927_);
  or (_37746_, _03928_, _03926_);
  and (_03929_, _03919_, _35830_);
  not (_03930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nor (_03931_, _03919_, _03930_);
  or (_37747_, _03931_, _03929_);
  and (_03932_, _03919_, _35834_);
  not (_03933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  nor (_03934_, _03919_, _03933_);
  or (_37748_, _03934_, _03932_);
  and (_03935_, _03919_, _35838_);
  not (_03936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  nor (_03937_, _03919_, _03936_);
  or (_37749_, _03937_, _03935_);
  and (_03938_, _03919_, _35842_);
  not (_03939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  nor (_03940_, _03919_, _03939_);
  or (_37750_, _03940_, _03938_);
  and (_03941_, _03919_, _35846_);
  not (_03942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  nor (_03943_, _03919_, _03942_);
  or (_37751_, _03943_, _03941_);
  and (_03944_, _03918_, _35817_);
  and (_03945_, _03944_, _35815_);
  not (_03946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  nor (_03947_, _03944_, _03946_);
  or (_37752_, _03947_, _03945_);
  and (_03948_, _03944_, _35822_);
  not (_03949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nor (_03950_, _03944_, _03949_);
  or (_37753_, _03950_, _03948_);
  and (_03951_, _03944_, _35826_);
  not (_03952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  nor (_03953_, _03944_, _03952_);
  or (_37754_, _03953_, _03951_);
  and (_03954_, _03944_, _35830_);
  not (_03955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nor (_03956_, _03944_, _03955_);
  or (_37755_, _03956_, _03954_);
  and (_03957_, _03944_, _35834_);
  not (_03958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  nor (_03959_, _03944_, _03958_);
  or (_37756_, _03959_, _03957_);
  and (_03960_, _03944_, _35838_);
  not (_03961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  nor (_03962_, _03944_, _03961_);
  or (_37757_, _03962_, _03960_);
  and (_03963_, _03944_, _35842_);
  not (_03964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  nor (_03965_, _03944_, _03964_);
  or (_37758_, _03965_, _03963_);
  and (_03966_, _03944_, _35846_);
  not (_03967_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  nor (_03968_, _03944_, _03967_);
  or (_37759_, _03968_, _03966_);
  and (_03969_, _03918_, _35851_);
  and (_03970_, _03969_, _35815_);
  not (_03971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nor (_03972_, _03969_, _03971_);
  or (_37760_, _03972_, _03970_);
  and (_03973_, _03969_, _35822_);
  not (_03974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  nor (_03975_, _03969_, _03974_);
  or (_37761_, _03975_, _03973_);
  and (_03976_, _03969_, _35826_);
  not (_03977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nor (_03978_, _03969_, _03977_);
  or (_37762_, _03978_, _03976_);
  and (_03979_, _03969_, _35830_);
  not (_03980_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  nor (_03981_, _03969_, _03980_);
  or (_37763_, _03981_, _03979_);
  and (_03982_, _03969_, _35834_);
  not (_03983_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nor (_03984_, _03969_, _03983_);
  or (_37764_, _03984_, _03982_);
  and (_03985_, _03969_, _35838_);
  not (_03986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  nor (_03987_, _03969_, _03986_);
  or (_37765_, _03987_, _03985_);
  and (_03988_, _03969_, _35842_);
  not (_03989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nor (_03990_, _03969_, _03989_);
  or (_37766_, _03990_, _03988_);
  and (_03991_, _03969_, _35846_);
  not (_03992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  nor (_03993_, _03969_, _03992_);
  or (_37767_, _03993_, _03991_);
  and (_03994_, _03918_, _35878_);
  and (_03995_, _03994_, _35815_);
  not (_03996_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nor (_03997_, _03994_, _03996_);
  or (_37768_, _03997_, _03995_);
  and (_03998_, _03994_, _35822_);
  not (_03999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nor (_04000_, _03994_, _03999_);
  or (_37769_, _04000_, _03998_);
  and (_04001_, _03994_, _35826_);
  not (_04002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  nor (_04003_, _03994_, _04002_);
  or (_37770_, _04003_, _04001_);
  and (_04004_, _03994_, _35830_);
  not (_04005_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nor (_04006_, _03994_, _04005_);
  or (_37771_, _04006_, _04004_);
  and (_04007_, _03994_, _35834_);
  not (_04008_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  nor (_04009_, _03994_, _04008_);
  or (_37772_, _04009_, _04007_);
  and (_04010_, _03994_, _35838_);
  not (_04011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  nor (_04012_, _03994_, _04011_);
  or (_37773_, _04012_, _04010_);
  and (_04013_, _03994_, _35842_);
  not (_04014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nor (_04015_, _03994_, _04014_);
  or (_37774_, _04015_, _04013_);
  and (_04016_, _03994_, _35846_);
  not (_04017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  nor (_04018_, _03994_, _04017_);
  or (_37775_, _04018_, _04016_);
  and (_04019_, _03918_, _35905_);
  and (_04020_, _04019_, _35815_);
  not (_04021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  nor (_04022_, _04019_, _04021_);
  or (_37776_, _04022_, _04020_);
  and (_04023_, _04019_, _35822_);
  not (_04024_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  nor (_04025_, _04019_, _04024_);
  or (_37777_, _04025_, _04023_);
  and (_04026_, _04019_, _35826_);
  not (_04027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nor (_04028_, _04019_, _04027_);
  or (_37778_, _04028_, _04026_);
  and (_04029_, _04019_, _35830_);
  not (_04030_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  nor (_04031_, _04019_, _04030_);
  or (_37779_, _04031_, _04029_);
  and (_04032_, _04019_, _35834_);
  not (_04033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nor (_04034_, _04019_, _04033_);
  or (_37780_, _04034_, _04032_);
  and (_04035_, _04019_, _35838_);
  not (_04036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  nor (_04037_, _04019_, _04036_);
  or (_37781_, _04037_, _04035_);
  and (_04038_, _04019_, _35842_);
  not (_04039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  nor (_04040_, _04019_, _04039_);
  or (_37782_, _04040_, _04038_);
  and (_04041_, _04019_, _35846_);
  not (_04042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  nor (_04043_, _04019_, _04042_);
  or (_37783_, _04043_, _04041_);
  and (_04044_, _03918_, _35931_);
  and (_04045_, _04044_, _35815_);
  not (_04046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nor (_04047_, _04044_, _04046_);
  or (_37784_, _04047_, _04045_);
  and (_04048_, _04044_, _35822_);
  not (_04049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  nor (_04050_, _04044_, _04049_);
  or (_37785_, _04050_, _04048_);
  and (_04051_, _04044_, _35826_);
  not (_04052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nor (_04053_, _04044_, _04052_);
  or (_37786_, _04053_, _04051_);
  and (_04054_, _04044_, _35830_);
  not (_04055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  nor (_04056_, _04044_, _04055_);
  or (_37787_, _04056_, _04054_);
  and (_04057_, _04044_, _35834_);
  not (_04058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  nor (_04059_, _04044_, _04058_);
  or (_37788_, _04059_, _04057_);
  and (_04060_, _04044_, _35838_);
  not (_04061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  nor (_04062_, _04044_, _04061_);
  or (_37789_, _04062_, _04060_);
  and (_04063_, _04044_, _35842_);
  not (_04064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  nor (_04065_, _04044_, _04064_);
  or (_37790_, _04065_, _04063_);
  and (_04066_, _04044_, _35846_);
  not (_04067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  nor (_04068_, _04044_, _04067_);
  or (_37791_, _04068_, _04066_);
  and (_04069_, _03918_, _35957_);
  and (_04070_, _04069_, _35815_);
  not (_04071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  nor (_04072_, _04069_, _04071_);
  or (_37792_, _04072_, _04070_);
  and (_04073_, _04069_, _35822_);
  not (_04074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nor (_04075_, _04069_, _04074_);
  or (_37793_, _04075_, _04073_);
  and (_04076_, _04069_, _35826_);
  not (_04077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  nor (_04078_, _04069_, _04077_);
  or (_37794_, _04078_, _04076_);
  and (_04079_, _04069_, _35830_);
  not (_04080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nor (_04081_, _04069_, _04080_);
  or (_37795_, _04081_, _04079_);
  and (_04082_, _04069_, _35834_);
  not (_04083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nor (_04084_, _04069_, _04083_);
  or (_37796_, _04084_, _04082_);
  and (_04085_, _04069_, _35838_);
  not (_04086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  nor (_04087_, _04069_, _04086_);
  or (_37797_, _04087_, _04085_);
  and (_04088_, _04069_, _35842_);
  not (_04089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nor (_04090_, _04069_, _04089_);
  or (_37798_, _04090_, _04088_);
  and (_04091_, _04069_, _35846_);
  not (_04092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  nor (_04093_, _04069_, _04092_);
  or (_37799_, _04093_, _04091_);
  and (_04094_, _03918_, _35983_);
  and (_04095_, _04094_, _35815_);
  not (_04096_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nor (_04097_, _04094_, _04096_);
  or (_37800_, _04097_, _04095_);
  and (_04098_, _04094_, _35822_);
  not (_04099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  nor (_04100_, _04094_, _04099_);
  or (_37801_, _04100_, _04098_);
  and (_04101_, _04094_, _35826_);
  not (_04102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  nor (_04103_, _04094_, _04102_);
  or (_37802_, _04103_, _04101_);
  and (_04104_, _04094_, _35830_);
  not (_04105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  nor (_04106_, _04094_, _04105_);
  or (_37803_, _04106_, _04104_);
  and (_04107_, _04094_, _35834_);
  not (_04108_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  nor (_04109_, _04094_, _04108_);
  or (_37804_, _04109_, _04107_);
  and (_04110_, _04094_, _35838_);
  not (_04111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  nor (_04112_, _04094_, _04111_);
  or (_37805_, _04112_, _04110_);
  and (_04113_, _04094_, _35842_);
  not (_04114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nor (_04115_, _04094_, _04114_);
  or (_37806_, _04115_, _04113_);
  and (_04116_, _04094_, _35846_);
  not (_04117_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  nor (_04118_, _04094_, _04117_);
  or (_37807_, _04118_, _04116_);
  and (_04119_, _03918_, _36010_);
  and (_04120_, _04119_, _35815_);
  not (_04121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  nor (_04122_, _04119_, _04121_);
  or (_37824_, _04122_, _04120_);
  and (_04123_, _04119_, _35822_);
  not (_04124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nor (_04125_, _04119_, _04124_);
  or (_37825_, _04125_, _04123_);
  and (_04126_, _04119_, _35826_);
  not (_04127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor (_04128_, _04119_, _04127_);
  or (_37826_, _04128_, _04126_);
  and (_04129_, _04119_, _35830_);
  not (_04130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nor (_04131_, _04119_, _04130_);
  or (_37827_, _04131_, _04129_);
  and (_04132_, _04119_, _35834_);
  not (_04133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor (_04134_, _04119_, _04133_);
  or (_37828_, _04134_, _04132_);
  and (_04135_, _04119_, _35838_);
  not (_04136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  nor (_04137_, _04119_, _04136_);
  or (_37829_, _04137_, _04135_);
  and (_04138_, _04119_, _35842_);
  not (_04139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  nor (_04140_, _04119_, _04139_);
  or (_37830_, _04140_, _04138_);
  and (_04141_, _04119_, _35846_);
  not (_04142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  nor (_04143_, _04119_, _04142_);
  or (_37831_, _04143_, _04141_);
  and (_04144_, _03918_, _36036_);
  and (_04145_, _04144_, _35815_);
  not (_04146_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nor (_04147_, _04144_, _04146_);
  or (_37832_, _04147_, _04145_);
  and (_04148_, _04144_, _35822_);
  not (_04149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  nor (_04150_, _04144_, _04149_);
  or (_37833_, _04150_, _04148_);
  and (_04151_, _04144_, _35826_);
  not (_04152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor (_04153_, _04144_, _04152_);
  or (_37834_, _04153_, _04151_);
  and (_04154_, _04144_, _35830_);
  not (_04155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  nor (_04156_, _04144_, _04155_);
  or (_37835_, _04156_, _04154_);
  and (_04157_, _04144_, _35834_);
  not (_04158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  nor (_04159_, _04144_, _04158_);
  or (_37836_, _04159_, _04157_);
  and (_04160_, _04144_, _35838_);
  not (_04161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  nor (_04162_, _04144_, _04161_);
  or (_37837_, _04162_, _04160_);
  and (_04163_, _04144_, _35842_);
  not (_04164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nor (_04165_, _04144_, _04164_);
  or (_37838_, _04165_, _04163_);
  and (_04166_, _04144_, _35846_);
  not (_04167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  nor (_04168_, _04144_, _04167_);
  or (_37839_, _04168_, _04166_);
  and (_04169_, _03918_, _36062_);
  and (_04170_, _04169_, _35815_);
  not (_04171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  nor (_04172_, _04169_, _04171_);
  or (_37840_, _04172_, _04170_);
  and (_04173_, _04169_, _35822_);
  not (_04174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor (_04175_, _04169_, _04174_);
  or (_37841_, _04175_, _04173_);
  and (_04176_, _04169_, _35826_);
  not (_04177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  nor (_04178_, _04169_, _04177_);
  or (_37842_, _04178_, _04176_);
  and (_04179_, _04169_, _35830_);
  not (_04180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor (_04181_, _04169_, _04180_);
  or (_37843_, _04181_, _04179_);
  and (_04182_, _04169_, _35834_);
  not (_04183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nor (_04184_, _04169_, _04183_);
  or (_37844_, _04184_, _04182_);
  and (_04185_, _04169_, _35838_);
  not (_04186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  nor (_04187_, _04169_, _04186_);
  or (_37845_, _04187_, _04185_);
  and (_04188_, _04169_, _35842_);
  not (_04189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  nor (_04190_, _04169_, _04189_);
  or (_37846_, _04190_, _04188_);
  and (_04191_, _04169_, _35846_);
  not (_04192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  nor (_04193_, _04169_, _04192_);
  or (_37847_, _04193_, _04191_);
  and (_04194_, _03918_, _36088_);
  and (_04195_, _04194_, _35815_);
  not (_04196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  nor (_04197_, _04194_, _04196_);
  or (_37848_, _04197_, _04195_);
  and (_04198_, _04194_, _35822_);
  not (_04199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor (_04200_, _04194_, _04199_);
  or (_37849_, _04200_, _04198_);
  and (_04201_, _04194_, _35826_);
  not (_04202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nor (_04203_, _04194_, _04202_);
  or (_37850_, _04203_, _04201_);
  and (_04204_, _04194_, _35830_);
  not (_04205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  nor (_04206_, _04194_, _04205_);
  or (_37851_, _04206_, _04204_);
  and (_04207_, _04194_, _35834_);
  not (_04208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  nor (_04209_, _04194_, _04208_);
  or (_37852_, _04209_, _04207_);
  and (_04210_, _04194_, _35838_);
  not (_04211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  nor (_04212_, _04194_, _04211_);
  or (_37853_, _04212_, _04210_);
  and (_04213_, _04194_, _35842_);
  not (_04214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor (_04215_, _04194_, _04214_);
  or (_37854_, _04215_, _04213_);
  and (_04216_, _04194_, _35846_);
  not (_04217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor (_04218_, _04194_, _04217_);
  or (_37855_, _04218_, _04216_);
  and (_04219_, _03918_, _36115_);
  and (_04220_, _04219_, _35815_);
  not (_04221_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nor (_04222_, _04219_, _04221_);
  or (_37856_, _04222_, _04220_);
  and (_04223_, _04219_, _35822_);
  not (_04224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  nor (_04225_, _04219_, _04224_);
  or (_37857_, _04225_, _04223_);
  and (_04226_, _04219_, _35826_);
  not (_04227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  nor (_04228_, _04219_, _04227_);
  or (_37858_, _04228_, _04226_);
  and (_04229_, _04219_, _35830_);
  not (_04230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nor (_04231_, _04219_, _04230_);
  or (_37859_, _04231_, _04229_);
  and (_04232_, _04219_, _35834_);
  not (_04233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor (_04234_, _04219_, _04233_);
  or (_37860_, _04234_, _04232_);
  and (_04235_, _04219_, _35838_);
  not (_04236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  nor (_04237_, _04219_, _04236_);
  or (_37861_, _04237_, _04235_);
  and (_04238_, _04219_, _35842_);
  not (_04239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  nor (_04240_, _04219_, _04239_);
  or (_37862_, _04240_, _04238_);
  and (_04241_, _04219_, _35846_);
  not (_04242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  nor (_04243_, _04219_, _04242_);
  or (_37863_, _04243_, _04241_);
  and (_04244_, _03918_, _36141_);
  and (_04245_, _04244_, _35815_);
  not (_04246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nor (_04247_, _04244_, _04246_);
  or (_37864_, _04247_, _04245_);
  and (_04248_, _04244_, _35822_);
  not (_04249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nor (_04250_, _04244_, _04249_);
  or (_37865_, _04250_, _04248_);
  and (_04251_, _04244_, _35826_);
  not (_04252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  nor (_04253_, _04244_, _04252_);
  or (_37866_, _04253_, _04251_);
  and (_04254_, _04244_, _35830_);
  not (_04255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nor (_04256_, _04244_, _04255_);
  or (_37867_, _04256_, _04254_);
  and (_04257_, _04244_, _35834_);
  not (_04258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  nor (_04259_, _04244_, _04258_);
  or (_37868_, _04259_, _04257_);
  and (_04260_, _04244_, _35838_);
  not (_04261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  nor (_04262_, _04244_, _04261_);
  or (_37869_, _04262_, _04260_);
  and (_04263_, _04244_, _35842_);
  not (_04264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  nor (_04265_, _04244_, _04264_);
  or (_37870_, _04265_, _04263_);
  and (_04266_, _04244_, _35846_);
  not (_04267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nor (_04268_, _04244_, _04267_);
  or (_37871_, _04268_, _04266_);
  and (_04269_, _03918_, _36167_);
  and (_04270_, _04269_, _35815_);
  not (_04271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  nor (_04272_, _04269_, _04271_);
  or (_37872_, _04272_, _04270_);
  and (_04273_, _04269_, _35822_);
  not (_04274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  nor (_04275_, _04269_, _04274_);
  or (_37873_, _04275_, _04273_);
  and (_04276_, _04269_, _35826_);
  not (_04277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor (_04278_, _04269_, _04277_);
  or (_37874_, _04278_, _04276_);
  and (_04279_, _04269_, _35830_);
  not (_04280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  nor (_04281_, _04269_, _04280_);
  or (_37875_, _04281_, _04279_);
  and (_04282_, _04269_, _35834_);
  not (_04283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nor (_04284_, _04269_, _04283_);
  or (_37876_, _04284_, _04282_);
  and (_04285_, _04269_, _35838_);
  not (_04286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  nor (_04287_, _04269_, _04286_);
  or (_37877_, _04287_, _04285_);
  and (_04288_, _04269_, _35842_);
  not (_04289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor (_04290_, _04269_, _04289_);
  or (_37878_, _04290_, _04288_);
  and (_04291_, _04269_, _35846_);
  not (_04292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  nor (_04293_, _04269_, _04292_);
  or (_37879_, _04293_, _04291_);
  and (_04294_, _03918_, _36193_);
  and (_04295_, _04294_, _35815_);
  not (_04296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor (_04297_, _04294_, _04296_);
  or (_37880_, _04297_, _04295_);
  and (_04298_, _04294_, _35822_);
  not (_04299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  nor (_04300_, _04294_, _04299_);
  or (_37881_, _04300_, _04298_);
  and (_04301_, _04294_, _35826_);
  not (_04302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor (_04303_, _04294_, _04302_);
  or (_37882_, _04303_, _04301_);
  and (_04304_, _04294_, _35830_);
  not (_04305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nor (_04306_, _04294_, _04305_);
  or (_37883_, _04306_, _04304_);
  and (_04307_, _04294_, _35834_);
  not (_04308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor (_04309_, _04294_, _04308_);
  or (_37884_, _04309_, _04307_);
  and (_04310_, _04294_, _35838_);
  not (_04311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  nor (_04312_, _04294_, _04311_);
  or (_37885_, _04312_, _04310_);
  and (_04313_, _04294_, _35842_);
  not (_04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  nor (_04315_, _04294_, _04314_);
  or (_37886_, _04315_, _04313_);
  and (_04316_, _04294_, _35846_);
  not (_04317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor (_04318_, _04294_, _04317_);
  or (_37887_, _04318_, _04316_);
  not (_04319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_04320_, _36220_, _34231_);
  and (_04321_, _04320_, _35572_);
  nor (_04322_, _04321_, _04319_);
  and (_04323_, _04321_, _35815_);
  or (_37888_, _04323_, _04322_);
  not (_04324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nor (_04325_, _04321_, _04324_);
  and (_04326_, _04321_, _35822_);
  or (_37889_, _04326_, _04325_);
  not (_04327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  nor (_04328_, _04321_, _04327_);
  and (_04329_, _04321_, _35826_);
  or (_37890_, _04329_, _04328_);
  not (_04330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  nor (_04331_, _04321_, _04330_);
  and (_04332_, _04321_, _35830_);
  or (_37891_, _04332_, _04331_);
  not (_04333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  nor (_04334_, _04321_, _04333_);
  and (_04335_, _04321_, _35834_);
  or (_37892_, _04335_, _04334_);
  not (_04336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  nor (_04337_, _04321_, _04336_);
  and (_04338_, _04321_, _35838_);
  or (_37893_, _04338_, _04337_);
  not (_04339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nor (_04340_, _04321_, _04339_);
  and (_04341_, _04321_, _35842_);
  or (_37894_, _04341_, _04340_);
  not (_04342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  nor (_04343_, _04321_, _04342_);
  and (_04344_, _04321_, _35846_);
  or (_37895_, _04344_, _04343_);
  not (_04345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and (_04346_, _04320_, _35817_);
  nor (_04347_, _04346_, _04345_);
  and (_04348_, _04346_, _35815_);
  or (_37896_, _04348_, _04347_);
  not (_04349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  nor (_04350_, _04346_, _04349_);
  and (_04351_, _04346_, _35822_);
  or (_37897_, _04351_, _04350_);
  not (_04352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nor (_04353_, _04346_, _04352_);
  and (_04354_, _04346_, _35826_);
  or (_37898_, _04354_, _04353_);
  not (_04355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  nor (_04356_, _04346_, _04355_);
  and (_04357_, _04346_, _35830_);
  or (_37899_, _04357_, _04356_);
  not (_04358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  nor (_04359_, _04346_, _04358_);
  and (_04360_, _04346_, _35834_);
  or (_37900_, _04360_, _04359_);
  not (_04361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  nor (_04362_, _04346_, _04361_);
  and (_04363_, _04346_, _35838_);
  or (_37901_, _04363_, _04362_);
  not (_04364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  nor (_04365_, _04346_, _04364_);
  and (_04366_, _04346_, _35842_);
  or (_37902_, _04366_, _04365_);
  not (_04367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  nor (_04368_, _04346_, _04367_);
  and (_04369_, _04346_, _35846_);
  or (_37903_, _04369_, _04368_);
  not (_04370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and (_04371_, _04320_, _35851_);
  nor (_04372_, _04371_, _04370_);
  and (_04373_, _04371_, _35815_);
  or (_37912_, _04373_, _04372_);
  not (_04374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nor (_04375_, _04371_, _04374_);
  and (_04376_, _04371_, _35822_);
  or (_37913_, _04376_, _04375_);
  not (_04377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  nor (_04378_, _04371_, _04377_);
  and (_04379_, _04371_, _35826_);
  or (_37914_, _04379_, _04378_);
  not (_04380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nor (_04381_, _04371_, _04380_);
  and (_04382_, _04371_, _35830_);
  or (_37915_, _04382_, _04381_);
  not (_04383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nor (_04384_, _04371_, _04383_);
  and (_04385_, _04371_, _35834_);
  or (_37916_, _04385_, _04384_);
  not (_04386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  nor (_04387_, _04371_, _04386_);
  and (_04388_, _04371_, _35838_);
  or (_37917_, _04388_, _04387_);
  not (_04389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nor (_04390_, _04371_, _04389_);
  and (_04391_, _04371_, _35842_);
  or (_37918_, _04391_, _04390_);
  not (_04392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  nor (_04393_, _04371_, _04392_);
  and (_04394_, _04371_, _35846_);
  or (_37919_, _04394_, _04393_);
  not (_04395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_04396_, _04320_, _35878_);
  nor (_04397_, _04396_, _04395_);
  and (_04398_, _04396_, _35815_);
  or (_37920_, _04398_, _04397_);
  not (_04399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nor (_04400_, _04396_, _04399_);
  and (_04401_, _04396_, _35822_);
  or (_37921_, _04401_, _04400_);
  not (_04402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nor (_04403_, _04396_, _04402_);
  and (_04404_, _04396_, _35826_);
  or (_37922_, _04404_, _04403_);
  not (_04405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  nor (_04406_, _04396_, _04405_);
  and (_04407_, _04396_, _35830_);
  or (_37923_, _04407_, _04406_);
  not (_04408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nor (_04409_, _04396_, _04408_);
  and (_04410_, _04396_, _35834_);
  or (_37924_, _04410_, _04409_);
  not (_04411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nor (_04412_, _04396_, _04411_);
  and (_04413_, _04396_, _35838_);
  or (_37925_, _04413_, _04412_);
  not (_04414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  nor (_04415_, _04396_, _04414_);
  and (_04416_, _04396_, _35842_);
  or (_37926_, _04416_, _04415_);
  not (_04417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  nor (_04418_, _04396_, _04417_);
  and (_04419_, _04396_, _35846_);
  or (_37927_, _04419_, _04418_);
  not (_04420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_04421_, _04320_, _35905_);
  nor (_04422_, _04421_, _04420_);
  and (_04423_, _04421_, _35815_);
  or (_37928_, _04423_, _04422_);
  not (_04424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  nor (_04425_, _04421_, _04424_);
  and (_04426_, _04421_, _35822_);
  or (_37929_, _04426_, _04425_);
  not (_04427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  nor (_04428_, _04421_, _04427_);
  and (_04429_, _04421_, _35826_);
  or (_37930_, _04429_, _04428_);
  not (_04430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nor (_04431_, _04421_, _04430_);
  and (_04432_, _04421_, _35830_);
  or (_37931_, _04432_, _04431_);
  not (_04433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  nor (_04434_, _04421_, _04433_);
  and (_04435_, _04421_, _35834_);
  or (_37932_, _04435_, _04434_);
  not (_04436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  nor (_04437_, _04421_, _04436_);
  and (_04438_, _04421_, _35838_);
  or (_37933_, _04438_, _04437_);
  not (_04439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nor (_04440_, _04421_, _04439_);
  and (_04441_, _04421_, _35842_);
  or (_37934_, _04441_, _04440_);
  not (_04442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  nor (_04443_, _04421_, _04442_);
  and (_04444_, _04421_, _35846_);
  or (_37935_, _04444_, _04443_);
  not (_04445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and (_04446_, _04320_, _35931_);
  nor (_04447_, _04446_, _04445_);
  and (_04448_, _04446_, _35815_);
  or (_37936_, _04448_, _04447_);
  not (_04449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  nor (_04450_, _04446_, _04449_);
  and (_04451_, _04446_, _35822_);
  or (_37937_, _04451_, _04450_);
  not (_04452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nor (_04453_, _04446_, _04452_);
  and (_04454_, _04446_, _35826_);
  or (_37938_, _04454_, _04453_);
  not (_04455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nor (_04456_, _04446_, _04455_);
  and (_04457_, _04446_, _35830_);
  or (_37939_, _04457_, _04456_);
  not (_04458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nor (_04459_, _04446_, _04458_);
  and (_04460_, _04446_, _35834_);
  or (_37940_, _04460_, _04459_);
  not (_04461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  nor (_04462_, _04446_, _04461_);
  and (_04463_, _04446_, _35838_);
  or (_37941_, _04463_, _04462_);
  not (_04464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  nor (_04465_, _04446_, _04464_);
  and (_04466_, _04446_, _35842_);
  or (_37942_, _04466_, _04465_);
  not (_04467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  nor (_04468_, _04446_, _04467_);
  and (_04469_, _04446_, _35846_);
  or (_37943_, _04469_, _04468_);
  not (_04470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and (_04471_, _04320_, _35957_);
  nor (_04472_, _04471_, _04470_);
  and (_04473_, _04471_, _35815_);
  or (_37944_, _04473_, _04472_);
  not (_04474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nor (_04475_, _04471_, _04474_);
  and (_04476_, _04471_, _35822_);
  or (_37945_, _04476_, _04475_);
  not (_04477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  nor (_04478_, _04471_, _04477_);
  and (_04479_, _04471_, _35826_);
  or (_37946_, _04479_, _04478_);
  not (_04480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  nor (_04481_, _04471_, _04480_);
  and (_04482_, _04471_, _35830_);
  or (_37947_, _04482_, _04481_);
  not (_04483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  nor (_04484_, _04471_, _04483_);
  and (_04485_, _04471_, _35834_);
  or (_37948_, _04485_, _04484_);
  not (_04486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  nor (_04487_, _04471_, _04486_);
  and (_04488_, _04471_, _35838_);
  or (_37949_, _04488_, _04487_);
  not (_04489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nor (_04490_, _04471_, _04489_);
  and (_04491_, _04471_, _35842_);
  or (_37950_, _04491_, _04490_);
  not (_04492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  nor (_04493_, _04471_, _04492_);
  and (_04494_, _04471_, _35846_);
  or (_37951_, _04494_, _04493_);
  not (_04495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_04496_, _04320_, _35983_);
  nor (_04497_, _04496_, _04495_);
  and (_04498_, _04496_, _35815_);
  or (_37952_, _04498_, _04497_);
  not (_04499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nor (_04500_, _04496_, _04499_);
  and (_04501_, _04496_, _35822_);
  or (_37953_, _04501_, _04500_);
  not (_04502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nor (_04503_, _04496_, _04502_);
  and (_04504_, _04496_, _35826_);
  or (_37954_, _04504_, _04503_);
  not (_04505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  nor (_04506_, _04496_, _04505_);
  and (_04507_, _04496_, _35830_);
  or (_37955_, _04507_, _04506_);
  not (_04508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  nor (_04509_, _04496_, _04508_);
  and (_04510_, _04496_, _35834_);
  or (_37956_, _04510_, _04509_);
  not (_04511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  nor (_04512_, _04496_, _04511_);
  and (_04513_, _04496_, _35838_);
  or (_37957_, _04513_, _04512_);
  not (_04514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nor (_04515_, _04496_, _04514_);
  and (_04516_, _04496_, _35842_);
  or (_37958_, _04516_, _04515_);
  not (_04517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  nor (_04518_, _04496_, _04517_);
  and (_04519_, _04496_, _35846_);
  or (_37959_, _04519_, _04518_);
  not (_04520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and (_04521_, _04320_, _36010_);
  nor (_04522_, _04521_, _04520_);
  and (_04523_, _04521_, _35815_);
  or (_37960_, _04523_, _04522_);
  not (_04524_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  nor (_04525_, _04521_, _04524_);
  and (_04526_, _04521_, _35822_);
  or (_37961_, _04526_, _04525_);
  not (_04527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  nor (_04528_, _04521_, _04527_);
  and (_04529_, _04521_, _35826_);
  or (_37962_, _04529_, _04528_);
  not (_04530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor (_04531_, _04521_, _04530_);
  and (_04532_, _04521_, _35830_);
  or (_37963_, _04532_, _04531_);
  not (_04533_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nor (_04534_, _04521_, _04533_);
  and (_04535_, _04521_, _35834_);
  or (_37964_, _04535_, _04534_);
  not (_04536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  nor (_04537_, _04521_, _04536_);
  and (_04538_, _04521_, _35838_);
  or (_37965_, _04538_, _04537_);
  not (_04539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  nor (_04540_, _04521_, _04539_);
  and (_04541_, _04521_, _35842_);
  or (_37966_, _04541_, _04540_);
  not (_04542_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  nor (_04543_, _04521_, _04542_);
  and (_04544_, _04521_, _35846_);
  or (_37967_, _04544_, _04543_);
  not (_04545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_04546_, _04320_, _36036_);
  nor (_04547_, _04546_, _04545_);
  and (_04548_, _04546_, _35815_);
  or (_37968_, _04548_, _04547_);
  not (_04549_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  nor (_04550_, _04546_, _04549_);
  and (_04551_, _04546_, _35822_);
  or (_37969_, _04551_, _04550_);
  not (_04552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  nor (_04553_, _04546_, _04552_);
  and (_04554_, _04546_, _35826_);
  or (_37970_, _04554_, _04553_);
  not (_04555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nor (_04556_, _04546_, _04555_);
  and (_04557_, _04546_, _35830_);
  or (_37971_, _04557_, _04556_);
  not (_04558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor (_04559_, _04546_, _04558_);
  and (_04560_, _04546_, _35834_);
  or (_37972_, _04560_, _04559_);
  not (_04561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  nor (_04562_, _04546_, _04561_);
  and (_04563_, _04546_, _35838_);
  or (_37973_, _04563_, _04562_);
  not (_04564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor (_04565_, _04546_, _04564_);
  and (_04566_, _04546_, _35842_);
  or (_37974_, _04566_, _04565_);
  not (_04567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  nor (_04568_, _04546_, _04567_);
  and (_04569_, _04546_, _35846_);
  or (_37975_, _04569_, _04568_);
  not (_04570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_04571_, _04320_, _36062_);
  nor (_04572_, _04571_, _04570_);
  and (_04573_, _04571_, _35815_);
  or (_37976_, _04573_, _04572_);
  not (_04574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor (_04575_, _04571_, _04574_);
  and (_04576_, _04571_, _35822_);
  or (_37977_, _04576_, _04575_);
  not (_04577_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor (_04578_, _04571_, _04577_);
  and (_04579_, _04571_, _35826_);
  or (_37978_, _04579_, _04578_);
  not (_04580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  nor (_04581_, _04571_, _04580_);
  and (_04582_, _04571_, _35830_);
  or (_37979_, _04582_, _04581_);
  not (_04583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  nor (_04584_, _04571_, _04583_);
  and (_04585_, _04571_, _35834_);
  or (_37980_, _04585_, _04584_);
  not (_04586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  nor (_04587_, _04571_, _04586_);
  and (_04588_, _04571_, _35838_);
  or (_37981_, _04588_, _04587_);
  not (_04589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  nor (_04590_, _04571_, _04589_);
  and (_04591_, _04571_, _35842_);
  or (_37982_, _04591_, _04590_);
  not (_04592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  nor (_04593_, _04571_, _04592_);
  and (_04594_, _04571_, _35846_);
  or (_37983_, _04594_, _04593_);
  not (_04595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and (_04596_, _04320_, _36088_);
  nor (_04597_, _04596_, _04595_);
  and (_04598_, _04596_, _35815_);
  or (_37984_, _04598_, _04597_);
  not (_04599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor (_04600_, _04596_, _04599_);
  and (_04601_, _04596_, _35822_);
  or (_37985_, _04601_, _04600_);
  not (_04602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  nor (_04603_, _04596_, _04602_);
  and (_04604_, _04596_, _35826_);
  or (_37986_, _04604_, _04603_);
  not (_04605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor (_04606_, _04596_, _04605_);
  and (_04607_, _04596_, _35830_);
  or (_37987_, _04607_, _04606_);
  not (_04608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor (_04609_, _04596_, _04608_);
  and (_04610_, _04596_, _35834_);
  or (_37988_, _04610_, _04609_);
  not (_04611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  nor (_04612_, _04596_, _04611_);
  and (_04613_, _04596_, _35838_);
  or (_37989_, _04613_, _04612_);
  not (_04614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nor (_04615_, _04596_, _04614_);
  and (_04616_, _04596_, _35842_);
  or (_37990_, _04616_, _04615_);
  not (_04617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  nor (_04618_, _04596_, _04617_);
  and (_04619_, _04596_, _35846_);
  or (_37991_, _04619_, _04618_);
  not (_04620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and (_04621_, _04320_, _36115_);
  nor (_04622_, _04621_, _04620_);
  and (_04623_, _04621_, _35815_);
  or (_38000_, _04623_, _04622_);
  not (_04624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  nor (_04625_, _04621_, _04624_);
  and (_04626_, _04621_, _35822_);
  or (_38001_, _04626_, _04625_);
  not (_04627_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor (_04628_, _04621_, _04627_);
  and (_04629_, _04621_, _35826_);
  or (_38002_, _04629_, _04628_);
  not (_04630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  nor (_04631_, _04621_, _04630_);
  and (_04632_, _04621_, _35830_);
  or (_38003_, _04632_, _04631_);
  not (_04633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  nor (_04634_, _04621_, _04633_);
  and (_04635_, _04621_, _35834_);
  or (_38004_, _04635_, _04634_);
  not (_04636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  nor (_04637_, _04621_, _04636_);
  and (_04638_, _04621_, _35838_);
  or (_38005_, _04638_, _04637_);
  not (_04639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  nor (_04640_, _04621_, _04639_);
  and (_04641_, _04621_, _35842_);
  or (_38006_, _04641_, _04640_);
  not (_04642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  nor (_04643_, _04621_, _04642_);
  and (_04644_, _04621_, _35846_);
  or (_38007_, _04644_, _04643_);
  not (_04645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_04646_, _04320_, _36141_);
  nor (_04647_, _04646_, _04645_);
  and (_04648_, _04646_, _35815_);
  or (_38008_, _04648_, _04647_);
  not (_04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor (_04650_, _04646_, _04649_);
  and (_04651_, _04646_, _35822_);
  or (_38009_, _04651_, _04650_);
  not (_04652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  nor (_04653_, _04646_, _04652_);
  and (_04654_, _04646_, _35826_);
  or (_38010_, _04654_, _04653_);
  not (_04655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nor (_04656_, _04646_, _04655_);
  and (_04657_, _04646_, _35830_);
  or (_38011_, _04657_, _04656_);
  not (_04658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  nor (_04659_, _04646_, _04658_);
  and (_04660_, _04646_, _35834_);
  or (_38012_, _04660_, _04659_);
  not (_04661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  nor (_04662_, _04646_, _04661_);
  and (_04663_, _04646_, _35838_);
  or (_38013_, _04663_, _04662_);
  not (_04664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor (_04665_, _04646_, _04664_);
  and (_04666_, _04646_, _35842_);
  or (_38014_, _04666_, _04665_);
  not (_04667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  nor (_04668_, _04646_, _04667_);
  and (_04669_, _04646_, _35846_);
  or (_38015_, _04669_, _04668_);
  not (_04670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_04671_, _04320_, _36167_);
  nor (_04672_, _04671_, _04670_);
  and (_04673_, _04671_, _35815_);
  or (_38016_, _04673_, _04672_);
  not (_04674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  nor (_04675_, _04671_, _04674_);
  and (_04676_, _04671_, _35822_);
  or (_38017_, _04676_, _04675_);
  not (_04677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nor (_04678_, _04671_, _04677_);
  and (_04679_, _04671_, _35826_);
  or (_38018_, _04679_, _04678_);
  not (_04680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  nor (_04681_, _04671_, _04680_);
  and (_04682_, _04671_, _35830_);
  or (_38019_, _04682_, _04681_);
  not (_04683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor (_04684_, _04671_, _04683_);
  and (_04685_, _04671_, _35834_);
  or (_38020_, _04685_, _04684_);
  not (_04686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  nor (_04687_, _04671_, _04686_);
  and (_04688_, _04671_, _35838_);
  or (_38021_, _04688_, _04687_);
  not (_04689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  nor (_04690_, _04671_, _04689_);
  and (_04691_, _04671_, _35842_);
  or (_38022_, _04691_, _04690_);
  not (_04692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor (_04693_, _04671_, _04692_);
  and (_04694_, _04671_, _35846_);
  or (_38023_, _04694_, _04693_);
  not (_04695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and (_04696_, _04320_, _36193_);
  nor (_04697_, _04696_, _04695_);
  and (_04698_, _04696_, _35815_);
  or (_38024_, _04698_, _04697_);
  not (_04699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  nor (_04700_, _04696_, _04699_);
  and (_04701_, _04696_, _35822_);
  or (_38025_, _04701_, _04700_);
  not (_04702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor (_04703_, _04696_, _04702_);
  and (_04704_, _04696_, _35826_);
  or (_38026_, _04704_, _04703_);
  not (_04705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  nor (_04706_, _04696_, _04705_);
  and (_04707_, _04696_, _35830_);
  or (_38027_, _04707_, _04706_);
  not (_04708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  nor (_04709_, _04696_, _04708_);
  and (_04710_, _04696_, _35834_);
  or (_38028_, _04710_, _04709_);
  not (_04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  nor (_04712_, _04696_, _04711_);
  and (_04713_, _04696_, _35838_);
  or (_38029_, _04713_, _04712_);
  not (_04714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  nor (_04715_, _04696_, _04714_);
  and (_04716_, _04696_, _35842_);
  or (_38030_, _04716_, _04715_);
  not (_04717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  nor (_04718_, _04696_, _04717_);
  and (_04719_, _04696_, _35846_);
  or (_38031_, _04719_, _04718_);
  and (_04720_, _36622_, _34231_);
  and (_04721_, _04720_, _35572_);
  and (_04722_, _04721_, _35815_);
  not (_04723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nor (_04724_, _04721_, _04723_);
  or (_38032_, _04724_, _04722_);
  and (_04725_, _04721_, _35822_);
  not (_04726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nor (_04727_, _04721_, _04726_);
  or (_38033_, _04727_, _04725_);
  and (_04728_, _04721_, _35826_);
  not (_04729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  nor (_04730_, _04721_, _04729_);
  or (_38034_, _04730_, _04728_);
  and (_04731_, _04721_, _35830_);
  not (_04732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nor (_04733_, _04721_, _04732_);
  or (_38035_, _04733_, _04731_);
  and (_04734_, _04721_, _35834_);
  not (_04735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nor (_04736_, _04721_, _04735_);
  or (_38036_, _04736_, _04734_);
  and (_04737_, _04721_, _35838_);
  not (_04738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  nor (_04739_, _04721_, _04738_);
  or (_38037_, _04739_, _04737_);
  and (_04740_, _04721_, _35842_);
  not (_04741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nor (_04742_, _04721_, _04741_);
  or (_38038_, _04742_, _04740_);
  and (_04743_, _04721_, _35846_);
  not (_04744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  nor (_04745_, _04721_, _04744_);
  or (_38039_, _04745_, _04743_);
  and (_04746_, _04720_, _35817_);
  and (_04747_, _04746_, _35815_);
  not (_04748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nor (_04749_, _04746_, _04748_);
  or (_38040_, _04749_, _04747_);
  and (_04750_, _04746_, _35822_);
  not (_04751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nor (_04752_, _04746_, _04751_);
  or (_38041_, _04752_, _04750_);
  and (_04753_, _04746_, _35826_);
  not (_04754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  nor (_04755_, _04746_, _04754_);
  or (_38042_, _04755_, _04753_);
  and (_04756_, _04746_, _35830_);
  not (_04757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  nor (_04758_, _04746_, _04757_);
  or (_38043_, _04758_, _04756_);
  and (_04759_, _04746_, _35834_);
  not (_04760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  nor (_04761_, _04746_, _04760_);
  or (_38044_, _04761_, _04759_);
  and (_04762_, _04746_, _35838_);
  not (_04763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nor (_04764_, _04746_, _04763_);
  or (_38045_, _04764_, _04762_);
  and (_04765_, _04746_, _35842_);
  not (_04766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  nor (_04767_, _04746_, _04766_);
  or (_38046_, _04767_, _04765_);
  and (_04768_, _04746_, _35846_);
  not (_04769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  nor (_04770_, _04746_, _04769_);
  or (_38047_, _04770_, _04768_);
  and (_04771_, _04720_, _35851_);
  and (_04772_, _04771_, _35815_);
  not (_04773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  nor (_04774_, _04771_, _04773_);
  or (_38048_, _04774_, _04772_);
  and (_04775_, _04771_, _35822_);
  not (_04776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  nor (_04777_, _04771_, _04776_);
  or (_38049_, _04777_, _04775_);
  and (_04778_, _04771_, _35826_);
  not (_04779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nor (_04780_, _04771_, _04779_);
  or (_38050_, _04780_, _04778_);
  and (_04781_, _04771_, _35830_);
  not (_04782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nor (_04783_, _04771_, _04782_);
  or (_38051_, _04783_, _04781_);
  and (_04784_, _04771_, _35834_);
  not (_04785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nor (_04786_, _04771_, _04785_);
  or (_38052_, _04786_, _04784_);
  and (_04787_, _04771_, _35838_);
  not (_04788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  nor (_04789_, _04771_, _04788_);
  or (_38053_, _04789_, _04787_);
  and (_04790_, _04771_, _35842_);
  not (_04791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nor (_04792_, _04771_, _04791_);
  or (_38054_, _04792_, _04790_);
  and (_04793_, _04771_, _35846_);
  not (_04794_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  nor (_04795_, _04771_, _04794_);
  or (_38055_, _04795_, _04793_);
  and (_04796_, _04720_, _35878_);
  and (_04797_, _04796_, _35815_);
  not (_04798_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nor (_04799_, _04796_, _04798_);
  or (_38056_, _04799_, _04797_);
  and (_04800_, _04796_, _35822_);
  not (_04801_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nor (_04802_, _04796_, _04801_);
  or (_38057_, _04802_, _04800_);
  and (_04803_, _04796_, _35826_);
  not (_04804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nor (_04805_, _04796_, _04804_);
  or (_38058_, _04805_, _04803_);
  and (_04806_, _04796_, _35830_);
  not (_04807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  nor (_04808_, _04796_, _04807_);
  or (_38059_, _04808_, _04806_);
  and (_04809_, _04796_, _35834_);
  not (_04810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  nor (_04811_, _04796_, _04810_);
  or (_38060_, _04811_, _04809_);
  and (_04812_, _04796_, _35838_);
  not (_04813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  nor (_04814_, _04796_, _04813_);
  or (_38061_, _04814_, _04812_);
  and (_04815_, _04796_, _35842_);
  not (_04816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nor (_04817_, _04796_, _04816_);
  or (_38062_, _04817_, _04815_);
  and (_04818_, _04796_, _35846_);
  not (_04819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  nor (_04820_, _04796_, _04819_);
  or (_38063_, _04820_, _04818_);
  and (_04821_, _04720_, _35905_);
  and (_04822_, _04821_, _35815_);
  not (_04823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  nor (_04824_, _04821_, _04823_);
  or (_38064_, _04824_, _04822_);
  and (_04825_, _04821_, _35822_);
  not (_04826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  nor (_04827_, _04821_, _04826_);
  or (_38065_, _04827_, _04825_);
  and (_04828_, _04821_, _35826_);
  not (_04829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  nor (_04830_, _04821_, _04829_);
  or (_38066_, _04830_, _04828_);
  and (_04831_, _04821_, _35830_);
  not (_04832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nor (_04833_, _04821_, _04832_);
  or (_38067_, _04833_, _04831_);
  and (_04834_, _04821_, _35834_);
  not (_04835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nor (_04836_, _04821_, _04835_);
  or (_38068_, _04836_, _04834_);
  and (_04837_, _04821_, _35838_);
  not (_04838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  nor (_04839_, _04821_, _04838_);
  or (_38069_, _04839_, _04837_);
  and (_04840_, _04821_, _35842_);
  not (_04841_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  nor (_04842_, _04821_, _04841_);
  or (_38070_, _04842_, _04840_);
  and (_04843_, _04821_, _35846_);
  not (_04844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  nor (_04845_, _04821_, _04844_);
  or (_38071_, _04845_, _04843_);
  and (_04846_, _04720_, _35931_);
  and (_04847_, _04846_, _35815_);
  not (_04848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nor (_04849_, _04846_, _04848_);
  or (_38072_, _04849_, _04847_);
  and (_04850_, _04846_, _35822_);
  not (_04851_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  nor (_04852_, _04846_, _04851_);
  or (_38073_, _04852_, _04850_);
  and (_04853_, _04846_, _35826_);
  not (_04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nor (_04855_, _04846_, _04854_);
  or (_38074_, _04855_, _04853_);
  and (_04856_, _04846_, _35830_);
  not (_04857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  nor (_04858_, _04846_, _04857_);
  or (_38075_, _04858_, _04856_);
  and (_04859_, _04846_, _35834_);
  not (_04860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  nor (_04861_, _04846_, _04860_);
  or (_38076_, _04861_, _04859_);
  and (_04862_, _04846_, _35838_);
  not (_04863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  nor (_04864_, _04846_, _04863_);
  or (_38077_, _04864_, _04862_);
  and (_04865_, _04846_, _35842_);
  not (_04866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  nor (_04867_, _04846_, _04866_);
  or (_38078_, _04867_, _04865_);
  and (_04868_, _04846_, _35846_);
  not (_04869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  nor (_04870_, _04846_, _04869_);
  or (_38079_, _04870_, _04868_);
  and (_04871_, _04720_, _35957_);
  and (_04872_, _04871_, _35815_);
  not (_04873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  nor (_04874_, _04871_, _04873_);
  or (_38088_, _04874_, _04872_);
  and (_04875_, _04871_, _35822_);
  not (_04876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nor (_04877_, _04871_, _04876_);
  or (_38089_, _04877_, _04875_);
  and (_04878_, _04871_, _35826_);
  not (_04879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  nor (_04880_, _04871_, _04879_);
  or (_38090_, _04880_, _04878_);
  and (_04881_, _04871_, _35830_);
  not (_04882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nor (_04883_, _04871_, _04882_);
  or (_38091_, _04883_, _04881_);
  and (_04884_, _04871_, _35834_);
  not (_04885_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nor (_04886_, _04871_, _04885_);
  or (_38092_, _04886_, _04884_);
  and (_04887_, _04871_, _35838_);
  not (_04888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  nor (_04889_, _04871_, _04888_);
  or (_38093_, _04889_, _04887_);
  and (_04890_, _04871_, _35842_);
  not (_04891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nor (_04892_, _04871_, _04891_);
  or (_38094_, _04892_, _04890_);
  and (_04893_, _04871_, _35846_);
  not (_04894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  nor (_04895_, _04871_, _04894_);
  or (_38095_, _04895_, _04893_);
  and (_04896_, _04720_, _35983_);
  and (_04897_, _04896_, _35815_);
  not (_04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  nor (_04899_, _04896_, _04898_);
  or (_38096_, _04899_, _04897_);
  and (_04900_, _04896_, _35822_);
  not (_04901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nor (_04902_, _04896_, _04901_);
  or (_38097_, _04902_, _04900_);
  and (_04903_, _04896_, _35826_);
  not (_04904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nor (_04905_, _04896_, _04904_);
  or (_38098_, _04905_, _04903_);
  and (_04906_, _04896_, _35830_);
  not (_04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  nor (_04908_, _04896_, _04907_);
  or (_38099_, _04908_, _04906_);
  and (_04909_, _04896_, _35834_);
  not (_04910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  nor (_04911_, _04896_, _04910_);
  or (_38100_, _04911_, _04909_);
  and (_04912_, _04896_, _35838_);
  not (_04913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  nor (_04914_, _04896_, _04913_);
  or (_38101_, _04914_, _04912_);
  and (_04915_, _04896_, _35842_);
  not (_04916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  nor (_04917_, _04896_, _04916_);
  or (_38102_, _04917_, _04915_);
  and (_04918_, _04896_, _35846_);
  not (_04919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  nor (_04920_, _04896_, _04919_);
  or (_38103_, _04920_, _04918_);
  and (_04921_, _04720_, _36010_);
  and (_04922_, _04921_, _35815_);
  not (_04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nor (_04924_, _04921_, _04923_);
  or (_38104_, _04924_, _04922_);
  and (_04925_, _04921_, _35822_);
  not (_04926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  nor (_04927_, _04921_, _04926_);
  or (_38105_, _04927_, _04925_);
  and (_04928_, _04921_, _35826_);
  not (_04929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  nor (_04930_, _04921_, _04929_);
  or (_38106_, _04930_, _04928_);
  and (_04931_, _04921_, _35830_);
  not (_04932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nor (_04933_, _04921_, _04932_);
  or (_38107_, _04933_, _04931_);
  and (_04934_, _04921_, _35834_);
  not (_04935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nor (_04936_, _04921_, _04935_);
  or (_38108_, _04936_, _04934_);
  and (_04937_, _04921_, _35838_);
  not (_04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  nor (_04939_, _04921_, _04938_);
  or (_38109_, _04939_, _04937_);
  and (_04940_, _04921_, _35842_);
  not (_04941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nor (_04942_, _04921_, _04941_);
  or (_38110_, _04942_, _04940_);
  and (_04943_, _04921_, _35846_);
  not (_04944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  nor (_04945_, _04921_, _04944_);
  or (_38111_, _04945_, _04943_);
  and (_04946_, _04720_, _36036_);
  and (_04947_, _04946_, _35815_);
  not (_04948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  nor (_04949_, _04946_, _04948_);
  or (_38112_, _04949_, _04947_);
  and (_04950_, _04946_, _35822_);
  not (_04951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nor (_04952_, _04946_, _04951_);
  or (_38113_, _04952_, _04950_);
  and (_04953_, _04946_, _35826_);
  not (_04954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nor (_04955_, _04946_, _04954_);
  or (_38114_, _04955_, _04953_);
  and (_04956_, _04946_, _35830_);
  not (_04957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  nor (_04958_, _04946_, _04957_);
  or (_38115_, _04958_, _04956_);
  and (_04959_, _04946_, _35834_);
  not (_04960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  nor (_04961_, _04946_, _04960_);
  or (_38116_, _04961_, _04959_);
  and (_04962_, _04946_, _35838_);
  not (_04963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  nor (_04964_, _04946_, _04963_);
  or (_38117_, _04964_, _04962_);
  and (_04965_, _04946_, _35842_);
  not (_04966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nor (_04967_, _04946_, _04966_);
  or (_38118_, _04967_, _04965_);
  and (_04968_, _04946_, _35846_);
  not (_04969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nor (_04970_, _04946_, _04969_);
  or (_38119_, _04970_, _04968_);
  and (_04971_, _04720_, _36062_);
  and (_04972_, _04971_, _35815_);
  not (_04973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor (_04974_, _04971_, _04973_);
  or (_38120_, _04974_, _04972_);
  and (_04975_, _04971_, _35822_);
  not (_04976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  nor (_04977_, _04971_, _04976_);
  or (_38121_, _04977_, _04975_);
  and (_04978_, _04971_, _35826_);
  not (_04979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  nor (_04980_, _04971_, _04979_);
  or (_38122_, _04980_, _04978_);
  and (_04981_, _04971_, _35830_);
  not (_04982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor (_04983_, _04971_, _04982_);
  or (_38123_, _04983_, _04981_);
  and (_04984_, _04971_, _35834_);
  not (_04985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nor (_04986_, _04971_, _04985_);
  or (_38124_, _04986_, _04984_);
  and (_04987_, _04971_, _35838_);
  not (_04988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  nor (_04989_, _04971_, _04988_);
  or (_38125_, _04989_, _04987_);
  and (_04990_, _04971_, _35842_);
  not (_04991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  nor (_04992_, _04971_, _04991_);
  or (_38126_, _04992_, _04990_);
  and (_04993_, _04971_, _35846_);
  not (_04994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  nor (_04995_, _04971_, _04994_);
  or (_38127_, _04995_, _04993_);
  and (_04996_, _04720_, _36088_);
  and (_04997_, _04996_, _35815_);
  not (_04998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor (_04999_, _04996_, _04998_);
  or (_38128_, _04999_, _04997_);
  and (_05000_, _04996_, _35822_);
  not (_05001_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  nor (_05002_, _04996_, _05001_);
  or (_38129_, _05002_, _05000_);
  and (_05003_, _04996_, _35826_);
  not (_05004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor (_05005_, _04996_, _05004_);
  or (_38130_, _05005_, _05003_);
  and (_05006_, _04996_, _35830_);
  not (_05007_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor (_05008_, _04996_, _05007_);
  or (_38131_, _05008_, _05006_);
  and (_05009_, _04996_, _35834_);
  not (_05010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  nor (_05011_, _04996_, _05010_);
  or (_38132_, _05011_, _05009_);
  and (_05012_, _04996_, _35838_);
  not (_05013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  nor (_05014_, _04996_, _05013_);
  or (_38133_, _05014_, _05012_);
  and (_05015_, _04996_, _35842_);
  not (_05016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor (_05017_, _04996_, _05016_);
  or (_38134_, _05017_, _05015_);
  and (_05018_, _04996_, _35846_);
  not (_05019_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nor (_05020_, _04996_, _05019_);
  or (_38135_, _05020_, _05018_);
  and (_05021_, _04720_, _36115_);
  and (_05022_, _05021_, _35815_);
  not (_05023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  nor (_05024_, _05021_, _05023_);
  or (_38136_, _05024_, _05022_);
  and (_05025_, _05021_, _35822_);
  not (_05026_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nor (_05027_, _05021_, _05026_);
  or (_38137_, _05027_, _05025_);
  and (_05028_, _05021_, _35826_);
  not (_05029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  nor (_05030_, _05021_, _05029_);
  or (_38138_, _05030_, _05028_);
  and (_05031_, _05021_, _35830_);
  not (_05032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  nor (_05033_, _05021_, _05032_);
  or (_38139_, _05033_, _05031_);
  and (_05034_, _05021_, _35834_);
  not (_05035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nor (_05036_, _05021_, _05035_);
  or (_38140_, _05036_, _05034_);
  and (_05037_, _05021_, _35838_);
  not (_05038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  nor (_05039_, _05021_, _05038_);
  or (_38141_, _05039_, _05037_);
  and (_05040_, _05021_, _35842_);
  not (_05041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  nor (_05042_, _05021_, _05041_);
  or (_38142_, _05042_, _05040_);
  and (_05043_, _05021_, _35846_);
  not (_05044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  nor (_05045_, _05021_, _05044_);
  or (_38143_, _05045_, _05043_);
  and (_05046_, _04720_, _36141_);
  and (_05047_, _05046_, _35815_);
  not (_05048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  nor (_05049_, _05046_, _05048_);
  or (_38144_, _05049_, _05047_);
  and (_05050_, _05046_, _35822_);
  not (_05051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nor (_05052_, _05046_, _05051_);
  or (_38145_, _05052_, _05050_);
  and (_05053_, _05046_, _35826_);
  not (_05054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nor (_05055_, _05046_, _05054_);
  or (_38146_, _05055_, _05053_);
  and (_05056_, _05046_, _35830_);
  not (_05057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  nor (_05058_, _05046_, _05057_);
  or (_38147_, _05058_, _05056_);
  and (_05059_, _05046_, _35834_);
  not (_05060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nor (_05061_, _05046_, _05060_);
  or (_38148_, _05061_, _05059_);
  and (_05062_, _05046_, _35838_);
  not (_05063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  nor (_05064_, _05046_, _05063_);
  or (_38149_, _05064_, _05062_);
  and (_05065_, _05046_, _35842_);
  not (_05066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nor (_05067_, _05046_, _05066_);
  or (_38150_, _05067_, _05065_);
  and (_05068_, _05046_, _35846_);
  not (_05069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  nor (_05070_, _05046_, _05069_);
  or (_38151_, _05070_, _05068_);
  and (_05071_, _04720_, _36167_);
  and (_05072_, _05071_, _35815_);
  not (_05073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor (_05074_, _05071_, _05073_);
  or (_38152_, _05074_, _05072_);
  and (_05075_, _05071_, _35822_);
  not (_05076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  nor (_05077_, _05071_, _05076_);
  or (_38153_, _05077_, _05075_);
  and (_05078_, _05071_, _35826_);
  not (_05079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  nor (_05080_, _05071_, _05079_);
  or (_38154_, _05080_, _05078_);
  and (_05081_, _05071_, _35830_);
  not (_05082_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor (_05083_, _05071_, _05082_);
  or (_38155_, _05083_, _05081_);
  and (_05084_, _05071_, _35834_);
  not (_05085_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  nor (_05086_, _05071_, _05085_);
  or (_38156_, _05086_, _05084_);
  and (_05087_, _05071_, _35838_);
  not (_05088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  nor (_05089_, _05071_, _05088_);
  or (_38157_, _05089_, _05087_);
  and (_05090_, _05071_, _35842_);
  not (_05091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  nor (_05092_, _05071_, _05091_);
  or (_38158_, _05092_, _05090_);
  and (_05093_, _05071_, _35846_);
  not (_05094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  nor (_05095_, _05071_, _05094_);
  or (_38159_, _05095_, _05093_);
  and (_05096_, _04720_, _36193_);
  and (_05097_, _05096_, _35815_);
  not (_05098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nor (_05099_, _05096_, _05098_);
  or (_38160_, _05099_, _05097_);
  and (_05100_, _05096_, _35822_);
  not (_05101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  nor (_05102_, _05096_, _05101_);
  or (_38161_, _05102_, _05100_);
  and (_05103_, _05096_, _35826_);
  not (_05104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor (_05105_, _05096_, _05104_);
  or (_38162_, _05105_, _05103_);
  and (_05106_, _05096_, _35830_);
  not (_05107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  nor (_05108_, _05096_, _05107_);
  or (_38163_, _05108_, _05106_);
  and (_05109_, _05096_, _35834_);
  not (_05110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor (_05111_, _05096_, _05110_);
  or (_38164_, _05111_, _05109_);
  and (_05112_, _05096_, _35838_);
  not (_05113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  nor (_05114_, _05096_, _05113_);
  or (_38165_, _05114_, _05112_);
  and (_05115_, _05096_, _35842_);
  not (_05116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  nor (_05117_, _05096_, _05116_);
  or (_38166_, _05117_, _05115_);
  and (_05118_, _05096_, _35846_);
  not (_05119_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  nor (_05120_, _05096_, _05119_);
  or (_38167_, _05120_, _05118_);
  and (_05121_, _00304_, _34231_);
  and (_05122_, _05121_, _35572_);
  and (_05123_, _05122_, _35815_);
  not (_05124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  nor (_05125_, _05122_, _05124_);
  or (_38176_, _05125_, _05123_);
  and (_05126_, _05122_, _35822_);
  not (_05127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nor (_05128_, _05122_, _05127_);
  or (_38177_, _05128_, _05126_);
  and (_05129_, _05122_, _35826_);
  not (_05130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  nor (_05131_, _05122_, _05130_);
  or (_38178_, _05131_, _05129_);
  and (_05132_, _05122_, _35830_);
  not (_05133_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nor (_05134_, _05122_, _05133_);
  or (_38179_, _05134_, _05132_);
  and (_05135_, _05122_, _35834_);
  not (_05136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  nor (_05137_, _05122_, _05136_);
  or (_38180_, _05137_, _05135_);
  and (_05138_, _05122_, _35838_);
  not (_05139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  nor (_05140_, _05122_, _05139_);
  or (_38181_, _05140_, _05138_);
  and (_05141_, _05122_, _35842_);
  not (_05142_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nor (_05143_, _05122_, _05142_);
  or (_38182_, _05143_, _05141_);
  and (_05144_, _05122_, _35846_);
  not (_05145_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  nor (_05146_, _05122_, _05145_);
  or (_38183_, _05146_, _05144_);
  and (_05147_, _05121_, _35817_);
  and (_05148_, _05147_, _35815_);
  not (_05149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nor (_05150_, _05147_, _05149_);
  or (_38184_, _05150_, _05148_);
  and (_05151_, _05147_, _35822_);
  not (_05152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nor (_05153_, _05147_, _05152_);
  or (_38185_, _05153_, _05151_);
  and (_05154_, _05147_, _35826_);
  not (_05155_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  nor (_05156_, _05147_, _05155_);
  or (_38186_, _05156_, _05154_);
  and (_05157_, _05147_, _35830_);
  not (_05158_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  nor (_05159_, _05147_, _05158_);
  or (_38187_, _05159_, _05157_);
  and (_05160_, _05147_, _35834_);
  not (_05161_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nor (_05162_, _05147_, _05161_);
  or (_38188_, _05162_, _05160_);
  and (_05163_, _05147_, _35838_);
  not (_05164_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  nor (_05165_, _05147_, _05164_);
  or (_38189_, _05165_, _05163_);
  and (_05166_, _05147_, _35842_);
  not (_05167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nor (_05168_, _05147_, _05167_);
  or (_38190_, _05168_, _05166_);
  and (_05169_, _05147_, _35846_);
  not (_05170_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  nor (_05171_, _05147_, _05170_);
  or (_38191_, _05171_, _05169_);
  and (_05172_, _05121_, _35851_);
  and (_05173_, _05172_, _35815_);
  not (_05174_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  nor (_05175_, _05172_, _05174_);
  or (_38192_, _05175_, _05173_);
  and (_05176_, _05172_, _35822_);
  not (_05177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  nor (_05178_, _05172_, _05177_);
  or (_38193_, _05178_, _05176_);
  and (_05179_, _05172_, _35826_);
  not (_05180_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nor (_05181_, _05172_, _05180_);
  or (_38194_, _05181_, _05179_);
  and (_05182_, _05172_, _35830_);
  not (_05183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nor (_05184_, _05172_, _05183_);
  or (_38195_, _05184_, _05182_);
  and (_05185_, _05172_, _35834_);
  not (_05186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  nor (_05187_, _05172_, _05186_);
  or (_38196_, _05187_, _05185_);
  and (_05188_, _05172_, _35838_);
  not (_05189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nor (_05190_, _05172_, _05189_);
  or (_38197_, _05190_, _05188_);
  and (_05191_, _05172_, _35842_);
  not (_05192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  nor (_05193_, _05172_, _05192_);
  or (_38198_, _05193_, _05191_);
  and (_05194_, _05172_, _35846_);
  not (_05195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  nor (_05196_, _05172_, _05195_);
  or (_38199_, _05196_, _05194_);
  and (_05197_, _05121_, _35878_);
  and (_05198_, _05197_, _35815_);
  not (_05199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  nor (_05200_, _05197_, _05199_);
  or (_38200_, _05200_, _05198_);
  and (_05201_, _05197_, _35822_);
  not (_05202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  nor (_05203_, _05197_, _05202_);
  or (_38201_, _05203_, _05201_);
  and (_05204_, _05197_, _35826_);
  not (_05205_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  nor (_05206_, _05197_, _05205_);
  or (_38202_, _05206_, _05204_);
  and (_05207_, _05197_, _35830_);
  not (_05208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nor (_05209_, _05197_, _05208_);
  or (_38203_, _05209_, _05207_);
  and (_05210_, _05197_, _35834_);
  not (_05211_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nor (_05212_, _05197_, _05211_);
  or (_38204_, _05212_, _05210_);
  and (_05213_, _05197_, _35838_);
  not (_05214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  nor (_05215_, _05197_, _05214_);
  or (_38205_, _05215_, _05213_);
  and (_05216_, _05197_, _35842_);
  not (_05217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nor (_05218_, _05197_, _05217_);
  or (_38206_, _05218_, _05216_);
  and (_05219_, _05197_, _35846_);
  not (_05220_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  nor (_05221_, _05197_, _05220_);
  or (_38207_, _05221_, _05219_);
  and (_05222_, _05121_, _35905_);
  and (_05223_, _05222_, _35815_);
  not (_05224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nor (_05225_, _05222_, _05224_);
  or (_38208_, _05225_, _05223_);
  and (_05226_, _05222_, _35822_);
  not (_05227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nor (_05228_, _05222_, _05227_);
  or (_38209_, _05228_, _05226_);
  and (_05229_, _05222_, _35826_);
  not (_05230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nor (_05231_, _05222_, _05230_);
  or (_38210_, _05231_, _05229_);
  and (_05232_, _05222_, _35830_);
  not (_05233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  nor (_05234_, _05222_, _05233_);
  or (_38211_, _05234_, _05232_);
  and (_05235_, _05222_, _35834_);
  not (_05236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  nor (_05237_, _05222_, _05236_);
  or (_38212_, _05237_, _05235_);
  and (_05238_, _05222_, _35838_);
  not (_05239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  nor (_05240_, _05222_, _05239_);
  or (_38213_, _05240_, _05238_);
  and (_05241_, _05222_, _35842_);
  not (_05242_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  nor (_05243_, _05222_, _05242_);
  or (_38214_, _05243_, _05241_);
  and (_05244_, _05222_, _35846_);
  not (_05245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  nor (_05246_, _05222_, _05245_);
  or (_38215_, _05246_, _05244_);
  and (_05247_, _05121_, _35931_);
  and (_05248_, _05247_, _35815_);
  not (_05249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nor (_05250_, _05247_, _05249_);
  or (_38216_, _05250_, _05248_);
  and (_05251_, _05247_, _35822_);
  not (_05252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  nor (_05253_, _05247_, _05252_);
  or (_38217_, _05253_, _05251_);
  and (_05254_, _05247_, _35826_);
  not (_05255_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nor (_05256_, _05247_, _05255_);
  or (_38218_, _05256_, _05254_);
  and (_05257_, _05247_, _35830_);
  not (_05258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  nor (_05259_, _05247_, _05258_);
  or (_38219_, _05259_, _05257_);
  and (_05260_, _05247_, _35834_);
  not (_05261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  nor (_05262_, _05247_, _05261_);
  or (_38220_, _05262_, _05260_);
  and (_05263_, _05247_, _35838_);
  not (_05264_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  nor (_05265_, _05247_, _05264_);
  or (_38221_, _05265_, _05263_);
  and (_05266_, _05247_, _35842_);
  not (_05267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  nor (_05268_, _05247_, _05267_);
  or (_38222_, _05268_, _05266_);
  and (_05269_, _05247_, _35846_);
  not (_05270_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  nor (_05271_, _05247_, _05270_);
  or (_38223_, _05271_, _05269_);
  and (_05272_, _05121_, _35957_);
  and (_05273_, _05272_, _35815_);
  not (_05274_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  nor (_05275_, _05272_, _05274_);
  or (_38224_, _05275_, _05273_);
  and (_05276_, _05272_, _35822_);
  not (_05277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nor (_05278_, _05272_, _05277_);
  or (_38225_, _05278_, _05276_);
  and (_05279_, _05272_, _35826_);
  not (_05280_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  nor (_05281_, _05272_, _05280_);
  or (_38226_, _05281_, _05279_);
  and (_05282_, _05272_, _35830_);
  not (_05283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nor (_05284_, _05272_, _05283_);
  or (_38227_, _05284_, _05282_);
  and (_05285_, _05272_, _35834_);
  not (_05286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nor (_05287_, _05272_, _05286_);
  or (_38228_, _05287_, _05285_);
  and (_05288_, _05272_, _35838_);
  not (_05289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  nor (_05290_, _05272_, _05289_);
  or (_38229_, _05290_, _05288_);
  and (_05291_, _05272_, _35842_);
  not (_05292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nor (_05293_, _05272_, _05292_);
  or (_38230_, _05293_, _05291_);
  and (_05294_, _05272_, _35846_);
  not (_05295_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  nor (_05296_, _05272_, _05295_);
  or (_38231_, _05296_, _05294_);
  and (_05297_, _05121_, _35983_);
  and (_05298_, _05297_, _35815_);
  not (_05299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  nor (_05300_, _05297_, _05299_);
  or (_38232_, _05300_, _05298_);
  and (_05301_, _05297_, _35822_);
  not (_05302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nor (_05303_, _05297_, _05302_);
  or (_38233_, _05303_, _05301_);
  and (_05304_, _05297_, _35826_);
  not (_05305_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nor (_05306_, _05297_, _05305_);
  or (_38234_, _05306_, _05304_);
  and (_05307_, _05297_, _35830_);
  not (_05308_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nor (_05309_, _05297_, _05308_);
  or (_38235_, _05309_, _05307_);
  and (_05310_, _05297_, _35834_);
  not (_05311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  nor (_05312_, _05297_, _05311_);
  or (_38236_, _05312_, _05310_);
  and (_05313_, _05297_, _35838_);
  not (_05314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  nor (_05315_, _05297_, _05314_);
  or (_38237_, _05315_, _05313_);
  and (_05316_, _05297_, _35842_);
  not (_05317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  nor (_05318_, _05297_, _05317_);
  or (_38238_, _05318_, _05316_);
  and (_05319_, _05297_, _35846_);
  not (_05320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  nor (_05321_, _05297_, _05320_);
  or (_38239_, _05321_, _05319_);
  and (_05322_, _05121_, _36010_);
  and (_05323_, _05322_, _35815_);
  not (_05324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor (_05325_, _05322_, _05324_);
  or (_38240_, _05325_, _05323_);
  and (_05326_, _05322_, _35822_);
  not (_05327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  nor (_05328_, _05322_, _05327_);
  or (_38241_, _05328_, _05326_);
  and (_05329_, _05322_, _35826_);
  not (_05330_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  nor (_05331_, _05322_, _05330_);
  or (_38242_, _05331_, _05329_);
  and (_05332_, _05322_, _35830_);
  not (_05333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  nor (_05334_, _05322_, _05333_);
  or (_38243_, _05334_, _05332_);
  and (_05335_, _05322_, _35834_);
  not (_05336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor (_05337_, _05322_, _05336_);
  or (_38244_, _05337_, _05335_);
  and (_05338_, _05322_, _35838_);
  not (_05339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  nor (_05340_, _05322_, _05339_);
  or (_38245_, _05340_, _05338_);
  and (_05341_, _05322_, _35842_);
  not (_05342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor (_05343_, _05322_, _05342_);
  or (_38246_, _05343_, _05341_);
  and (_05344_, _05322_, _35846_);
  not (_05345_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  nor (_05346_, _05322_, _05345_);
  or (_38247_, _05346_, _05344_);
  and (_05347_, _05121_, _36036_);
  and (_05348_, _05347_, _35815_);
  not (_05349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  nor (_05350_, _05347_, _05349_);
  or (_38248_, _05350_, _05348_);
  and (_05351_, _05347_, _35822_);
  not (_05352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  nor (_05353_, _05347_, _05352_);
  or (_38249_, _05353_, _05351_);
  and (_05354_, _05347_, _35826_);
  not (_05355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  nor (_05356_, _05347_, _05355_);
  or (_38250_, _05356_, _05354_);
  and (_05357_, _05347_, _35830_);
  not (_05358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  nor (_05359_, _05347_, _05358_);
  or (_38251_, _05359_, _05357_);
  and (_05360_, _05347_, _35834_);
  not (_05361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  nor (_05362_, _05347_, _05361_);
  or (_38252_, _05362_, _05360_);
  and (_05363_, _05347_, _35838_);
  not (_05364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  nor (_05365_, _05347_, _05364_);
  or (_38253_, _05365_, _05363_);
  and (_05366_, _05347_, _35842_);
  not (_05367_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nor (_05368_, _05347_, _05367_);
  or (_38254_, _05368_, _05366_);
  and (_05369_, _05347_, _35846_);
  not (_05370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  nor (_05371_, _05347_, _05370_);
  or (_38255_, _05371_, _05369_);
  and (_05372_, _05121_, _36062_);
  and (_05373_, _05372_, _35815_);
  not (_05374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor (_05375_, _05372_, _05374_);
  or (_38264_, _05375_, _05373_);
  and (_05376_, _05372_, _35822_);
  not (_05377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor (_05378_, _05372_, _05377_);
  or (_38265_, _05378_, _05376_);
  and (_05379_, _05372_, _35826_);
  not (_05380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor (_05381_, _05372_, _05380_);
  or (_38266_, _05381_, _05379_);
  and (_05382_, _05372_, _35830_);
  not (_05383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor (_05384_, _05372_, _05383_);
  or (_38267_, _05384_, _05382_);
  and (_05385_, _05372_, _35834_);
  not (_05386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor (_05387_, _05372_, _05386_);
  or (_38268_, _05387_, _05385_);
  and (_05388_, _05372_, _35838_);
  not (_05389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nor (_05390_, _05372_, _05389_);
  or (_38269_, _05390_, _05388_);
  and (_05391_, _05372_, _35842_);
  not (_05392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  nor (_05393_, _05372_, _05392_);
  or (_38270_, _05393_, _05391_);
  and (_05394_, _05372_, _35846_);
  not (_05395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  nor (_05396_, _05372_, _05395_);
  or (_38271_, _05396_, _05394_);
  and (_05397_, _05121_, _36088_);
  and (_05398_, _05397_, _35815_);
  not (_05399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor (_05400_, _05397_, _05399_);
  or (_38272_, _05400_, _05398_);
  and (_05401_, _05397_, _35822_);
  not (_05402_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  nor (_05403_, _05397_, _05402_);
  or (_38273_, _05403_, _05401_);
  and (_05404_, _05397_, _35826_);
  not (_05405_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  nor (_05406_, _05397_, _05405_);
  or (_38274_, _05406_, _05404_);
  and (_05407_, _05397_, _35830_);
  not (_05408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  nor (_05409_, _05397_, _05408_);
  or (_38275_, _05409_, _05407_);
  and (_05410_, _05397_, _35834_);
  not (_05411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  nor (_05412_, _05397_, _05411_);
  or (_38276_, _05412_, _05410_);
  and (_05413_, _05397_, _35838_);
  not (_05414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  nor (_05415_, _05397_, _05414_);
  or (_38277_, _05415_, _05413_);
  and (_05416_, _05397_, _35842_);
  not (_05417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor (_05418_, _05397_, _05417_);
  or (_38278_, _05418_, _05416_);
  and (_05419_, _05397_, _35846_);
  not (_05420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  nor (_05421_, _05397_, _05420_);
  or (_38279_, _05421_, _05419_);
  and (_05422_, _05121_, _36115_);
  and (_05423_, _05422_, _35815_);
  not (_05424_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  nor (_05425_, _05422_, _05424_);
  or (_38280_, _05425_, _05423_);
  and (_05426_, _05422_, _35822_);
  not (_05427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor (_05428_, _05422_, _05427_);
  or (_38281_, _05428_, _05426_);
  and (_05429_, _05422_, _35826_);
  not (_05430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor (_05431_, _05422_, _05430_);
  or (_38282_, _05431_, _05429_);
  and (_05432_, _05422_, _35830_);
  not (_05433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor (_05434_, _05422_, _05433_);
  or (_38283_, _05434_, _05432_);
  and (_05435_, _05422_, _35834_);
  not (_05436_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor (_05437_, _05422_, _05436_);
  or (_38284_, _05437_, _05435_);
  and (_05438_, _05422_, _35838_);
  not (_05439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor (_05440_, _05422_, _05439_);
  or (_38285_, _05440_, _05438_);
  and (_05441_, _05422_, _35842_);
  not (_05442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor (_05443_, _05422_, _05442_);
  or (_38286_, _05443_, _05441_);
  and (_05444_, _05422_, _35846_);
  not (_05445_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  nor (_05446_, _05422_, _05445_);
  or (_38287_, _05446_, _05444_);
  and (_05447_, _05121_, _36141_);
  and (_05448_, _05447_, _35815_);
  not (_05449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  nor (_05450_, _05447_, _05449_);
  or (_38288_, _05450_, _05448_);
  and (_05451_, _05447_, _35822_);
  not (_05452_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor (_05453_, _05447_, _05452_);
  or (_38289_, _05453_, _05451_);
  and (_05454_, _05447_, _35826_);
  not (_05455_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  nor (_05456_, _05447_, _05455_);
  or (_38290_, _05456_, _05454_);
  and (_05457_, _05447_, _35830_);
  not (_05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor (_05459_, _05447_, _05458_);
  or (_38291_, _05459_, _05457_);
  and (_05460_, _05447_, _35834_);
  not (_05461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  nor (_05462_, _05447_, _05461_);
  or (_38292_, _05462_, _05460_);
  and (_05463_, _05447_, _35838_);
  not (_05464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  nor (_05465_, _05447_, _05464_);
  or (_38293_, _05465_, _05463_);
  and (_05466_, _05447_, _35842_);
  not (_05467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  nor (_05468_, _05447_, _05467_);
  or (_38294_, _05468_, _05466_);
  and (_05469_, _05447_, _35846_);
  not (_05470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  nor (_05471_, _05447_, _05470_);
  or (_38295_, _05471_, _05469_);
  and (_05472_, _05121_, _36167_);
  and (_05473_, _05472_, _35815_);
  not (_05474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor (_05475_, _05472_, _05474_);
  or (_38296_, _05475_, _05473_);
  and (_05476_, _05472_, _35822_);
  not (_05477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  nor (_05478_, _05472_, _05477_);
  or (_38297_, _05478_, _05476_);
  and (_05479_, _05472_, _35826_);
  not (_05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor (_05481_, _05472_, _05480_);
  or (_38298_, _05481_, _05479_);
  and (_05482_, _05472_, _35830_);
  not (_05483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  nor (_05484_, _05472_, _05483_);
  or (_38299_, _05484_, _05482_);
  and (_05485_, _05472_, _35834_);
  not (_05486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nor (_05487_, _05472_, _05486_);
  or (_38300_, _05487_, _05485_);
  and (_05488_, _05472_, _35838_);
  not (_05489_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  nor (_05490_, _05472_, _05489_);
  or (_38301_, _05490_, _05488_);
  and (_05491_, _05472_, _35842_);
  not (_05492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor (_05493_, _05472_, _05492_);
  or (_38302_, _05493_, _05491_);
  and (_05494_, _05472_, _35846_);
  not (_05495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  nor (_05496_, _05472_, _05495_);
  or (_38303_, _05496_, _05494_);
  and (_05497_, _05121_, _36193_);
  and (_05498_, _05497_, _35815_);
  not (_05499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  nor (_05500_, _05497_, _05499_);
  or (_38304_, _05500_, _05498_);
  and (_05501_, _05497_, _35822_);
  not (_05502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  nor (_05503_, _05497_, _05502_);
  or (_38305_, _05503_, _05501_);
  and (_05504_, _05497_, _35826_);
  not (_05505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  nor (_05506_, _05497_, _05505_);
  or (_38306_, _05506_, _05504_);
  and (_05507_, _05497_, _35830_);
  not (_05508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  nor (_05509_, _05497_, _05508_);
  or (_38307_, _05509_, _05507_);
  and (_05510_, _05497_, _35834_);
  not (_05511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  nor (_05512_, _05497_, _05511_);
  or (_38308_, _05512_, _05510_);
  and (_05513_, _05497_, _35838_);
  not (_05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  nor (_05515_, _05497_, _05514_);
  or (_38309_, _05515_, _05513_);
  and (_05516_, _05497_, _35842_);
  not (_05517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  nor (_05518_, _05497_, _05517_);
  or (_38310_, _05518_, _05516_);
  and (_05519_, _05497_, _35846_);
  not (_05520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  nor (_05521_, _05497_, _05520_);
  or (_38311_, _05521_, _05519_);
  and (_05522_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_05523_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_05524_, _05523_, _05522_);
  and (_05525_, _05524_, _34581_);
  and (_05526_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_05527_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_05528_, _05527_, _05526_);
  and (_05529_, _05528_, _34796_);
  or (_05530_, _05529_, _05525_);
  and (_05531_, _05530_, _34772_);
  and (_05532_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_05533_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_05534_, _05533_, _05532_);
  and (_05535_, _05534_, _34581_);
  and (_05536_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_05537_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_05538_, _05537_, _05536_);
  and (_05539_, _05538_, _34796_);
  or (_05540_, _05539_, _05535_);
  and (_05541_, _05540_, _34790_);
  or (_05542_, _05541_, _34719_);
  or (_05543_, _05542_, _05531_);
  or (_05544_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_05545_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_05546_, _05545_, _34796_);
  and (_05547_, _05546_, _05544_);
  or (_05548_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_05549_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_05550_, _05549_, _34581_);
  and (_05551_, _05550_, _05548_);
  or (_05552_, _05551_, _05547_);
  and (_05553_, _05552_, _34772_);
  or (_05554_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_05555_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_05556_, _05555_, _34796_);
  and (_05557_, _05556_, _05554_);
  or (_05558_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_05559_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_05560_, _05559_, _34581_);
  and (_05561_, _05560_, _05558_);
  or (_05562_, _05561_, _05557_);
  and (_05563_, _05562_, _34790_);
  or (_05564_, _05563_, _34803_);
  or (_05565_, _05564_, _05553_);
  and (_05566_, _05565_, _05543_);
  or (_05567_, _05566_, _34700_);
  and (_05568_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_05569_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_05570_, _05569_, _05568_);
  and (_05571_, _05570_, _34581_);
  and (_05572_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_05573_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_05574_, _05573_, _05572_);
  and (_05575_, _05574_, _34796_);
  or (_05576_, _05575_, _05571_);
  and (_05577_, _05576_, _34772_);
  and (_05578_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_05579_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_05580_, _05579_, _05578_);
  and (_05581_, _05580_, _34581_);
  and (_05582_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_05583_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_05584_, _05583_, _05582_);
  and (_05585_, _05584_, _34796_);
  or (_05586_, _05585_, _05581_);
  and (_05587_, _05586_, _34790_);
  or (_05588_, _05587_, _34719_);
  or (_05589_, _05588_, _05577_);
  or (_05590_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_05591_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_05592_, _05591_, _05590_);
  and (_05593_, _05592_, _34581_);
  or (_05594_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_05595_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_05596_, _05595_, _05594_);
  and (_05597_, _05596_, _34796_);
  or (_05598_, _05597_, _05593_);
  and (_05599_, _05598_, _34772_);
  or (_05600_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_05601_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_05602_, _05601_, _05600_);
  and (_05603_, _05602_, _34581_);
  or (_05604_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_05605_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_05606_, _05605_, _05604_);
  and (_05607_, _05606_, _34796_);
  or (_05608_, _05607_, _05603_);
  and (_05609_, _05608_, _34790_);
  or (_05610_, _05609_, _34803_);
  or (_05611_, _05610_, _05599_);
  and (_05612_, _05611_, _05589_);
  or (_05613_, _05612_, _34789_);
  and (_05614_, _05613_, _34638_);
  and (_05615_, _05614_, _05567_);
  and (_05616_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_05617_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_05618_, _05617_, _05616_);
  and (_05619_, _05618_, _34581_);
  and (_05620_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_05621_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_05622_, _05621_, _05620_);
  and (_05623_, _05622_, _34796_);
  or (_05624_, _05623_, _05619_);
  or (_05625_, _05624_, _34790_);
  and (_05626_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_05627_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_05628_, _05627_, _05626_);
  and (_05629_, _05628_, _34581_);
  and (_05630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_05631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_05632_, _05631_, _05630_);
  and (_05633_, _05632_, _34796_);
  or (_05634_, _05633_, _05629_);
  or (_05635_, _05634_, _34772_);
  and (_05636_, _05635_, _34803_);
  and (_05637_, _05636_, _05625_);
  or (_05638_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_05639_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_05640_, _05639_, _05638_);
  and (_05641_, _05640_, _34581_);
  or (_05642_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_05643_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_05644_, _05643_, _05642_);
  and (_05645_, _05644_, _34796_);
  or (_05646_, _05645_, _05641_);
  or (_05647_, _05646_, _34790_);
  or (_05648_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_05649_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_05650_, _05649_, _05648_);
  and (_05651_, _05650_, _34581_);
  or (_05652_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_05653_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_05654_, _05653_, _05652_);
  and (_05655_, _05654_, _34796_);
  or (_05656_, _05655_, _05651_);
  or (_05657_, _05656_, _34772_);
  and (_05658_, _05657_, _34719_);
  and (_05659_, _05658_, _05647_);
  or (_05660_, _05659_, _05637_);
  or (_05661_, _05660_, _34789_);
  and (_05662_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_05663_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_05664_, _05663_, _05662_);
  and (_05665_, _05664_, _34581_);
  and (_05666_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_05667_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_05668_, _05667_, _05666_);
  and (_05669_, _05668_, _34796_);
  or (_05670_, _05669_, _05665_);
  or (_05671_, _05670_, _34790_);
  and (_05672_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_05673_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_05674_, _05673_, _05672_);
  and (_05675_, _05674_, _34581_);
  and (_05676_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_05677_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_05678_, _05677_, _05676_);
  and (_05679_, _05678_, _34796_);
  or (_05680_, _05679_, _05675_);
  or (_05681_, _05680_, _34772_);
  and (_05682_, _05681_, _34803_);
  and (_05683_, _05682_, _05671_);
  or (_05684_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_05685_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_05686_, _05685_, _34796_);
  and (_05687_, _05686_, _05684_);
  or (_05688_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_05689_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_05690_, _05689_, _34581_);
  and (_05691_, _05690_, _05688_);
  or (_05692_, _05691_, _05687_);
  or (_05693_, _05692_, _34790_);
  or (_05694_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_05695_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_05696_, _05695_, _34796_);
  and (_05697_, _05696_, _05694_);
  or (_05698_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_05699_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_05700_, _05699_, _34581_);
  and (_05701_, _05700_, _05698_);
  or (_05702_, _05701_, _05697_);
  or (_05703_, _05702_, _34772_);
  and (_05704_, _05703_, _34719_);
  and (_05705_, _05704_, _05693_);
  or (_05706_, _05705_, _05683_);
  or (_05707_, _05706_, _34700_);
  and (_05708_, _05707_, _34840_);
  and (_05709_, _05708_, _05661_);
  or (_05710_, _05709_, _05615_);
  or (_05711_, _05710_, _34692_);
  and (_05712_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_05713_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_05714_, _05713_, _05712_);
  and (_05715_, _05714_, _34581_);
  and (_05716_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_05717_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_05718_, _05717_, _05716_);
  and (_05719_, _05718_, _34796_);
  or (_05720_, _05719_, _05715_);
  and (_05721_, _05720_, _34790_);
  and (_05722_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_05723_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_05724_, _05723_, _05722_);
  and (_05725_, _05724_, _34581_);
  and (_05726_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_05727_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_05728_, _05727_, _05726_);
  and (_05729_, _05728_, _34796_);
  or (_05730_, _05729_, _05725_);
  and (_05731_, _05730_, _34772_);
  or (_05732_, _05731_, _05721_);
  and (_05733_, _05732_, _34803_);
  or (_05734_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_05735_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_05736_, _05735_, _05734_);
  and (_05737_, _05736_, _34581_);
  or (_05738_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_05739_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_05740_, _05739_, _05738_);
  and (_05741_, _05740_, _34796_);
  or (_05742_, _05741_, _05737_);
  and (_05743_, _05742_, _34790_);
  or (_05744_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_05745_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_05746_, _05745_, _05744_);
  and (_05747_, _05746_, _34581_);
  or (_05748_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_05749_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_05750_, _05749_, _05748_);
  and (_05751_, _05750_, _34796_);
  or (_05752_, _05751_, _05747_);
  and (_05753_, _05752_, _34772_);
  or (_05754_, _05753_, _05743_);
  and (_05755_, _05754_, _34719_);
  or (_05756_, _05755_, _05733_);
  or (_05757_, _05756_, _34789_);
  and (_05758_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_05759_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_05760_, _05759_, _05758_);
  and (_05761_, _05760_, _34581_);
  and (_05762_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_05763_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_05764_, _05763_, _05762_);
  and (_05765_, _05764_, _34796_);
  or (_05766_, _05765_, _05761_);
  and (_05767_, _05766_, _34790_);
  and (_05768_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_05769_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_05770_, _05769_, _05768_);
  and (_05771_, _05770_, _34581_);
  and (_05772_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and (_05773_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_05774_, _05773_, _05772_);
  and (_05775_, _05774_, _34796_);
  or (_05776_, _05775_, _05771_);
  and (_05777_, _05776_, _34772_);
  or (_05778_, _05777_, _05767_);
  and (_05779_, _05778_, _34803_);
  or (_05780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_05781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and (_05782_, _05781_, _34796_);
  and (_05783_, _05782_, _05780_);
  or (_05784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_05785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and (_05786_, _05785_, _34581_);
  and (_05787_, _05786_, _05784_);
  or (_05788_, _05787_, _05783_);
  and (_05789_, _05788_, _34790_);
  or (_05790_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_05791_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_05792_, _05791_, _34796_);
  and (_05793_, _05792_, _05790_);
  or (_05794_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_05795_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_05796_, _05795_, _34581_);
  and (_05797_, _05796_, _05794_);
  or (_05798_, _05797_, _05793_);
  and (_05799_, _05798_, _34772_);
  or (_05800_, _05799_, _05789_);
  and (_05801_, _05800_, _34719_);
  or (_05802_, _05801_, _05779_);
  or (_05803_, _05802_, _34700_);
  and (_05804_, _05803_, _34638_);
  and (_05805_, _05804_, _05757_);
  and (_05806_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_05807_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_05808_, _05807_, _05806_);
  and (_05809_, _05808_, _34581_);
  and (_05810_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_05811_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_05812_, _05811_, _05810_);
  and (_05813_, _05812_, _34796_);
  or (_05814_, _05813_, _05809_);
  or (_05815_, _05814_, _34790_);
  and (_05816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_05817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_05818_, _05817_, _05816_);
  and (_05819_, _05818_, _34581_);
  and (_05820_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_05821_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_05822_, _05821_, _05820_);
  and (_05823_, _05822_, _34796_);
  or (_05824_, _05823_, _05819_);
  or (_05825_, _05824_, _34772_);
  and (_05826_, _05825_, _34803_);
  and (_05827_, _05826_, _05815_);
  or (_05828_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_05829_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_05830_, _05829_, _34796_);
  and (_05831_, _05830_, _05828_);
  or (_05832_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_05833_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_05834_, _05833_, _34581_);
  and (_05835_, _05834_, _05832_);
  or (_05836_, _05835_, _05831_);
  or (_05837_, _05836_, _34790_);
  or (_05838_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_05839_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_05840_, _05839_, _34796_);
  and (_05841_, _05840_, _05838_);
  or (_05842_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_05843_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_05844_, _05843_, _34581_);
  and (_05845_, _05844_, _05842_);
  or (_05846_, _05845_, _05841_);
  or (_05847_, _05846_, _34772_);
  and (_05848_, _05847_, _34719_);
  and (_05849_, _05848_, _05837_);
  or (_05850_, _05849_, _05827_);
  or (_05851_, _05850_, _34700_);
  and (_05852_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_05853_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_05854_, _05853_, _05852_);
  and (_05855_, _05854_, _34581_);
  and (_05856_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_05857_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_05858_, _05857_, _05856_);
  and (_05859_, _05858_, _34796_);
  or (_05860_, _05859_, _05855_);
  or (_05861_, _05860_, _34790_);
  and (_05862_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_05863_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_05864_, _05863_, _05862_);
  and (_05865_, _05864_, _34581_);
  and (_05866_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_05867_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_05868_, _05867_, _05866_);
  and (_05869_, _05868_, _34796_);
  or (_05870_, _05869_, _05865_);
  or (_05871_, _05870_, _34772_);
  and (_05872_, _05871_, _34803_);
  and (_05873_, _05872_, _05861_);
  or (_05874_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_05875_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_05876_, _05875_, _05874_);
  and (_05877_, _05876_, _34581_);
  or (_05878_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_05879_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_05880_, _05879_, _05878_);
  and (_05881_, _05880_, _34796_);
  or (_05882_, _05881_, _05877_);
  or (_05883_, _05882_, _34790_);
  or (_05884_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_05885_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_05886_, _05885_, _05884_);
  and (_05887_, _05886_, _34581_);
  or (_05888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_05889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_05890_, _05889_, _05888_);
  and (_05891_, _05890_, _34796_);
  or (_05892_, _05891_, _05887_);
  or (_05893_, _05892_, _34772_);
  and (_05894_, _05893_, _34719_);
  and (_05895_, _05894_, _05883_);
  or (_05896_, _05895_, _05873_);
  or (_05897_, _05896_, _34789_);
  and (_05898_, _05897_, _34840_);
  and (_05899_, _05898_, _05851_);
  or (_05900_, _05899_, _05805_);
  or (_05901_, _05900_, _34985_);
  and (_05902_, _05901_, _34346_);
  and (_05903_, _05902_, _05711_);
  and (_05904_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_05905_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_05906_, _05905_, _05904_);
  and (_05907_, _05906_, _34581_);
  and (_05908_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_05909_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_05910_, _05909_, _05908_);
  and (_05911_, _05910_, _34796_);
  or (_05912_, _05911_, _05907_);
  or (_05913_, _05912_, _34790_);
  and (_05914_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_05915_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_05916_, _05915_, _05914_);
  and (_05917_, _05916_, _34581_);
  and (_05918_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_05919_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_05920_, _05919_, _05918_);
  and (_05921_, _05920_, _34796_);
  or (_05922_, _05921_, _05917_);
  or (_05923_, _05922_, _34772_);
  and (_05924_, _05923_, _34803_);
  and (_05925_, _05924_, _05913_);
  or (_05926_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_05927_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_05928_, _05927_, _05926_);
  and (_05929_, _05928_, _34581_);
  or (_05930_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_05931_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_05932_, _05931_, _05930_);
  and (_05933_, _05932_, _34796_);
  or (_05934_, _05933_, _05929_);
  or (_05935_, _05934_, _34790_);
  or (_05936_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_05937_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_05938_, _05937_, _05936_);
  and (_05939_, _05938_, _34581_);
  or (_05940_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_05941_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_05942_, _05941_, _05940_);
  and (_05943_, _05942_, _34796_);
  or (_05944_, _05943_, _05939_);
  or (_05945_, _05944_, _34772_);
  and (_05946_, _05945_, _34719_);
  and (_05947_, _05946_, _05935_);
  or (_05948_, _05947_, _05925_);
  and (_05949_, _05948_, _34700_);
  and (_05950_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_05951_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_05952_, _05951_, _05950_);
  and (_05953_, _05952_, _34581_);
  and (_05954_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_05955_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_05956_, _05955_, _05954_);
  and (_05957_, _05956_, _34796_);
  or (_05958_, _05957_, _05953_);
  or (_05959_, _05958_, _34790_);
  and (_05960_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_05961_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_05962_, _05961_, _05960_);
  and (_05963_, _05962_, _34581_);
  and (_05964_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_05965_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_05966_, _05965_, _05964_);
  and (_05967_, _05966_, _34796_);
  or (_05968_, _05967_, _05963_);
  or (_05969_, _05968_, _34772_);
  and (_05970_, _05969_, _34803_);
  and (_05971_, _05970_, _05959_);
  or (_05972_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_05973_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_05974_, _05973_, _34796_);
  and (_05975_, _05974_, _05972_);
  or (_05976_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_05977_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_05978_, _05977_, _34581_);
  and (_05979_, _05978_, _05976_);
  or (_05980_, _05979_, _05975_);
  or (_05981_, _05980_, _34790_);
  or (_05982_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_05983_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_05984_, _05983_, _34796_);
  and (_05985_, _05984_, _05982_);
  or (_05986_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_05987_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_05988_, _05987_, _34581_);
  and (_05989_, _05988_, _05986_);
  or (_05990_, _05989_, _05985_);
  or (_05991_, _05990_, _34772_);
  and (_05992_, _05991_, _34719_);
  and (_05993_, _05992_, _05981_);
  or (_05994_, _05993_, _05971_);
  and (_05995_, _05994_, _34789_);
  or (_05996_, _05995_, _05949_);
  and (_05997_, _05996_, _34840_);
  and (_05998_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and (_05999_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_06000_, _05999_, _05998_);
  and (_06001_, _06000_, _34581_);
  and (_06002_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_06003_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_06004_, _06003_, _06002_);
  and (_06005_, _06004_, _34796_);
  or (_06006_, _06005_, _06001_);
  and (_06007_, _06006_, _34772_);
  and (_06008_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_06009_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_06010_, _06009_, _06008_);
  and (_06011_, _06010_, _34581_);
  and (_06012_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_06013_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_06014_, _06013_, _06012_);
  and (_06015_, _06014_, _34796_);
  or (_06016_, _06015_, _06011_);
  and (_06017_, _06016_, _34790_);
  or (_06018_, _06017_, _06007_);
  and (_06019_, _06018_, _34803_);
  or (_06020_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_06021_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_06022_, _06021_, _34796_);
  and (_06023_, _06022_, _06020_);
  or (_06024_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_06025_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and (_06026_, _06025_, _34581_);
  and (_06027_, _06026_, _06024_);
  or (_06028_, _06027_, _06023_);
  and (_06029_, _06028_, _34772_);
  or (_06030_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_06031_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_06032_, _06031_, _34796_);
  and (_06033_, _06032_, _06030_);
  or (_06034_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_06035_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_06036_, _06035_, _34581_);
  and (_06037_, _06036_, _06034_);
  or (_06038_, _06037_, _06033_);
  and (_06039_, _06038_, _34790_);
  or (_06040_, _06039_, _06029_);
  and (_06041_, _06040_, _34719_);
  or (_06042_, _06041_, _06019_);
  and (_06043_, _06042_, _34789_);
  and (_06044_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_06045_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_06046_, _06045_, _06044_);
  and (_06047_, _06046_, _34581_);
  and (_06048_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_06049_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_06050_, _06049_, _06048_);
  and (_06051_, _06050_, _34796_);
  or (_06052_, _06051_, _06047_);
  and (_06053_, _06052_, _34772_);
  and (_06054_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_06055_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_06056_, _06055_, _06054_);
  and (_06057_, _06056_, _34581_);
  and (_06058_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_06059_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_06060_, _06059_, _06058_);
  and (_06061_, _06060_, _34796_);
  or (_06062_, _06061_, _06057_);
  and (_06063_, _06062_, _34790_);
  or (_06064_, _06063_, _06053_);
  and (_06065_, _06064_, _34803_);
  or (_06066_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_06067_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_06068_, _06067_, _06066_);
  and (_06069_, _06068_, _34581_);
  or (_06070_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_06071_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_06072_, _06071_, _06070_);
  and (_06073_, _06072_, _34796_);
  or (_06074_, _06073_, _06069_);
  and (_06075_, _06074_, _34772_);
  or (_06076_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_06077_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_06078_, _06077_, _06076_);
  and (_06079_, _06078_, _34581_);
  or (_06080_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_06081_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_06082_, _06081_, _06080_);
  and (_06083_, _06082_, _34796_);
  or (_06084_, _06083_, _06079_);
  and (_06085_, _06084_, _34790_);
  or (_06086_, _06085_, _06075_);
  and (_06087_, _06086_, _34719_);
  or (_06088_, _06087_, _06065_);
  and (_06089_, _06088_, _34700_);
  or (_06090_, _06089_, _06043_);
  and (_06091_, _06090_, _34638_);
  or (_06092_, _06091_, _05997_);
  or (_06093_, _06092_, _34985_);
  or (_06094_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_06095_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_06096_, _06095_, _06094_);
  and (_06097_, _06096_, _34581_);
  or (_06098_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_06099_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_06100_, _06099_, _06098_);
  and (_06101_, _06100_, _34796_);
  or (_06102_, _06101_, _06097_);
  and (_06103_, _06102_, _34790_);
  or (_06104_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_06105_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_06106_, _06105_, _06104_);
  and (_06107_, _06106_, _34581_);
  or (_06108_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_06109_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_06110_, _06109_, _06108_);
  and (_06111_, _06110_, _34796_);
  or (_06112_, _06111_, _06107_);
  and (_06113_, _06112_, _34772_);
  or (_06114_, _06113_, _06103_);
  and (_06115_, _06114_, _34719_);
  and (_06116_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_06117_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_06118_, _06117_, _06116_);
  and (_06119_, _06118_, _34581_);
  and (_06120_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_06121_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_06122_, _06121_, _06120_);
  and (_06123_, _06122_, _34796_);
  or (_06124_, _06123_, _06119_);
  and (_06125_, _06124_, _34790_);
  and (_06126_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_06127_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_06128_, _06127_, _06126_);
  and (_06129_, _06128_, _34581_);
  and (_06130_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_06131_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_06132_, _06131_, _06130_);
  and (_06133_, _06132_, _34796_);
  or (_06134_, _06133_, _06129_);
  and (_06135_, _06134_, _34772_);
  or (_06136_, _06135_, _06125_);
  and (_06137_, _06136_, _34803_);
  or (_06138_, _06137_, _06115_);
  and (_06139_, _06138_, _34700_);
  or (_06140_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_06141_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_06142_, _06141_, _34796_);
  and (_06143_, _06142_, _06140_);
  or (_06144_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_06145_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_06146_, _06145_, _34581_);
  and (_06147_, _06146_, _06144_);
  or (_06148_, _06147_, _06143_);
  and (_06149_, _06148_, _34790_);
  or (_06150_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_06151_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_06152_, _06151_, _34796_);
  and (_06153_, _06152_, _06150_);
  or (_06154_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_06155_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_06156_, _06155_, _34581_);
  and (_06157_, _06156_, _06154_);
  or (_06158_, _06157_, _06153_);
  and (_06159_, _06158_, _34772_);
  or (_06160_, _06159_, _06149_);
  and (_06161_, _06160_, _34719_);
  and (_06162_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_06163_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_06164_, _06163_, _06162_);
  and (_06165_, _06164_, _34581_);
  and (_06166_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_06167_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_06168_, _06167_, _06166_);
  and (_06169_, _06168_, _34796_);
  or (_06170_, _06169_, _06165_);
  and (_06171_, _06170_, _34790_);
  and (_06172_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_06173_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_06174_, _06173_, _06172_);
  and (_06175_, _06174_, _34581_);
  and (_06176_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_06177_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_06178_, _06177_, _06176_);
  and (_06179_, _06178_, _34796_);
  or (_06180_, _06179_, _06175_);
  and (_06181_, _06180_, _34772_);
  or (_06182_, _06181_, _06171_);
  and (_06183_, _06182_, _34803_);
  or (_06184_, _06183_, _06161_);
  and (_06185_, _06184_, _34789_);
  or (_06186_, _06185_, _06139_);
  and (_06187_, _06186_, _34638_);
  and (_06188_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_06189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_06190_, _06189_, _06188_);
  and (_06191_, _06190_, _34581_);
  and (_06192_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_06193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_06194_, _06193_, _06192_);
  and (_06195_, _06194_, _34796_);
  or (_06196_, _06195_, _06191_);
  or (_06197_, _06196_, _34790_);
  and (_06198_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_06199_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_06200_, _06199_, _06198_);
  and (_06201_, _06200_, _34581_);
  and (_06202_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_06203_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_06204_, _06203_, _06202_);
  and (_06205_, _06204_, _34796_);
  or (_06206_, _06205_, _06201_);
  or (_06207_, _06206_, _34772_);
  and (_06208_, _06207_, _34803_);
  and (_06209_, _06208_, _06197_);
  or (_06210_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_06211_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_06212_, _06211_, _34796_);
  and (_06213_, _06212_, _06210_);
  or (_06214_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_06215_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_06216_, _06215_, _34581_);
  and (_06217_, _06216_, _06214_);
  or (_06218_, _06217_, _06213_);
  or (_06219_, _06218_, _34790_);
  or (_06220_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_06221_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_06222_, _06221_, _34796_);
  and (_06223_, _06222_, _06220_);
  or (_06224_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_06225_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_06226_, _06225_, _34581_);
  and (_06227_, _06226_, _06224_);
  or (_06228_, _06227_, _06223_);
  or (_06229_, _06228_, _34772_);
  and (_06230_, _06229_, _34719_);
  and (_06231_, _06230_, _06219_);
  or (_06232_, _06231_, _06209_);
  and (_06233_, _06232_, _34789_);
  and (_06234_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_06235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_06236_, _06235_, _06234_);
  and (_06237_, _06236_, _34581_);
  and (_06238_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_06239_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_06240_, _06239_, _06238_);
  and (_06241_, _06240_, _34796_);
  or (_06242_, _06241_, _06237_);
  or (_06243_, _06242_, _34790_);
  and (_06244_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_06245_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_06246_, _06245_, _06244_);
  and (_06247_, _06246_, _34581_);
  and (_06248_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_06249_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_06250_, _06249_, _06248_);
  and (_06251_, _06250_, _34796_);
  or (_06252_, _06251_, _06247_);
  or (_06253_, _06252_, _34772_);
  and (_06254_, _06253_, _34803_);
  and (_06255_, _06254_, _06243_);
  or (_06256_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_06257_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_06258_, _06257_, _06256_);
  and (_06259_, _06258_, _34581_);
  or (_06260_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_06261_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_06262_, _06261_, _06260_);
  and (_06263_, _06262_, _34796_);
  or (_06264_, _06263_, _06259_);
  or (_06265_, _06264_, _34790_);
  or (_06266_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_06267_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_06268_, _06267_, _06266_);
  and (_06269_, _06268_, _34581_);
  or (_06270_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_06271_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_06272_, _06271_, _06270_);
  and (_06273_, _06272_, _34796_);
  or (_06274_, _06273_, _06269_);
  or (_06275_, _06274_, _34772_);
  and (_06276_, _06275_, _34719_);
  and (_06277_, _06276_, _06265_);
  or (_06278_, _06277_, _06255_);
  and (_06279_, _06278_, _34700_);
  or (_06280_, _06279_, _06233_);
  and (_06281_, _06280_, _34840_);
  or (_06282_, _06281_, _06187_);
  or (_06283_, _06282_, _34692_);
  and (_06284_, _06283_, _35178_);
  and (_06285_, _06284_, _06093_);
  or (_06286_, _06285_, _05903_);
  or (_06287_, _06286_, _34788_);
  or (_06288_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_06289_, _06288_, _38997_);
  and (_38984_[0], _06289_, _06287_);
  and (_06290_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_06291_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_06292_, _06291_, _06290_);
  and (_06293_, _06292_, _34796_);
  and (_06294_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_06295_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_06296_, _06295_, _06294_);
  and (_06297_, _06296_, _34581_);
  or (_06298_, _06297_, _06293_);
  or (_06299_, _06298_, _34790_);
  and (_06300_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_06301_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_06302_, _06301_, _06300_);
  and (_06303_, _06302_, _34796_);
  and (_06304_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_06305_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_06306_, _06305_, _06304_);
  and (_06307_, _06306_, _34581_);
  or (_06308_, _06307_, _06303_);
  or (_06309_, _06308_, _34772_);
  and (_06310_, _06309_, _34803_);
  and (_06311_, _06310_, _06299_);
  or (_06312_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_06313_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_06314_, _06313_, _34581_);
  and (_06315_, _06314_, _06312_);
  or (_06316_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_06317_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_06318_, _06317_, _34796_);
  and (_06319_, _06318_, _06316_);
  or (_06320_, _06319_, _06315_);
  or (_06321_, _06320_, _34790_);
  or (_06322_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_06323_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_06324_, _06323_, _34581_);
  and (_06325_, _06324_, _06322_);
  or (_06326_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_06327_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_06328_, _06327_, _34796_);
  and (_06329_, _06328_, _06326_);
  or (_06330_, _06329_, _06325_);
  or (_06331_, _06330_, _34772_);
  and (_06332_, _06331_, _34719_);
  and (_06333_, _06332_, _06321_);
  or (_06334_, _06333_, _06311_);
  or (_06335_, _06334_, _34700_);
  and (_06336_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_06337_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_06338_, _06337_, _34581_);
  or (_06339_, _06338_, _06336_);
  and (_06340_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_06341_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_06342_, _06341_, _34796_);
  or (_06343_, _06342_, _06340_);
  and (_06344_, _06343_, _06339_);
  or (_06345_, _06344_, _34790_);
  and (_06346_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_06347_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_06348_, _06347_, _34581_);
  or (_06349_, _06348_, _06346_);
  and (_06350_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_06351_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_06352_, _06351_, _34796_);
  or (_06353_, _06352_, _06350_);
  and (_06354_, _06353_, _06349_);
  or (_06355_, _06354_, _34772_);
  and (_06356_, _06355_, _34803_);
  and (_06357_, _06356_, _06345_);
  or (_06358_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_06359_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_06360_, _06359_, _06358_);
  or (_06361_, _06360_, _34796_);
  or (_06362_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_06363_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_06364_, _06363_, _06362_);
  or (_06365_, _06364_, _34581_);
  and (_06366_, _06365_, _06361_);
  or (_06367_, _06366_, _34790_);
  or (_06368_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_06369_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_06370_, _06369_, _06368_);
  or (_06371_, _06370_, _34796_);
  or (_06372_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_06373_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_06374_, _06373_, _06372_);
  or (_06375_, _06374_, _34581_);
  and (_06376_, _06375_, _06371_);
  or (_06377_, _06376_, _34772_);
  and (_06378_, _06377_, _34719_);
  and (_06379_, _06378_, _06367_);
  or (_06380_, _06379_, _06357_);
  or (_06381_, _06380_, _34789_);
  and (_06382_, _06381_, _34840_);
  and (_06383_, _06382_, _06335_);
  and (_06384_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_06385_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_06386_, _06385_, _06384_);
  and (_06387_, _06386_, _34581_);
  and (_06388_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_06389_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_06390_, _06389_, _06388_);
  and (_06391_, _06390_, _34796_);
  or (_06392_, _06391_, _06387_);
  and (_06393_, _06392_, _34772_);
  and (_06394_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_06395_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_06396_, _06395_, _06394_);
  and (_06397_, _06396_, _34581_);
  and (_06398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_06399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_06400_, _06399_, _06398_);
  and (_06401_, _06400_, _34796_);
  or (_06402_, _06401_, _06397_);
  and (_06403_, _06402_, _34790_);
  or (_06404_, _06403_, _06393_);
  and (_06405_, _06404_, _34803_);
  or (_06406_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_06407_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_06408_, _06407_, _06406_);
  and (_06409_, _06408_, _34581_);
  or (_06410_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_06411_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_06412_, _06411_, _06410_);
  and (_06413_, _06412_, _34796_);
  or (_06414_, _06413_, _06409_);
  and (_06415_, _06414_, _34772_);
  or (_06416_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_06417_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_06418_, _06417_, _06416_);
  and (_06419_, _06418_, _34581_);
  or (_06420_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_06421_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_06422_, _06421_, _06420_);
  and (_06423_, _06422_, _34796_);
  or (_06424_, _06423_, _06419_);
  and (_06425_, _06424_, _34790_);
  or (_06426_, _06425_, _06415_);
  and (_06427_, _06426_, _34719_);
  or (_06428_, _06427_, _06405_);
  and (_06429_, _06428_, _34789_);
  and (_06430_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_06431_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_06432_, _06431_, _06430_);
  and (_06433_, _06432_, _34581_);
  and (_06434_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_06435_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_06436_, _06435_, _06434_);
  and (_06437_, _06436_, _34796_);
  or (_06438_, _06437_, _06433_);
  and (_06439_, _06438_, _34772_);
  and (_06440_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_06441_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_06442_, _06441_, _06440_);
  and (_06443_, _06442_, _34581_);
  and (_06444_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_06445_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_06446_, _06445_, _06444_);
  and (_06447_, _06446_, _34796_);
  or (_06448_, _06447_, _06443_);
  and (_06449_, _06448_, _34790_);
  or (_06450_, _06449_, _06439_);
  and (_06451_, _06450_, _34803_);
  or (_06452_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_06453_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_06454_, _06453_, _06452_);
  and (_06455_, _06454_, _34581_);
  or (_06456_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_06457_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_06458_, _06457_, _06456_);
  and (_06459_, _06458_, _34796_);
  or (_06460_, _06459_, _06455_);
  and (_06461_, _06460_, _34772_);
  or (_06462_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_06463_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_06464_, _06463_, _06462_);
  and (_06465_, _06464_, _34581_);
  or (_06466_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_06467_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_06468_, _06467_, _06466_);
  and (_06469_, _06468_, _34796_);
  or (_06470_, _06469_, _06465_);
  and (_06471_, _06470_, _34790_);
  or (_06472_, _06471_, _06461_);
  and (_06473_, _06472_, _34719_);
  or (_06474_, _06473_, _06451_);
  and (_06475_, _06474_, _34700_);
  or (_06476_, _06475_, _06429_);
  and (_06477_, _06476_, _34638_);
  or (_06478_, _06477_, _06383_);
  or (_06479_, _06478_, _34692_);
  and (_06480_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_06481_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_06482_, _06481_, _06480_);
  and (_06483_, _06482_, _34581_);
  and (_06484_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_06485_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_06486_, _06485_, _06484_);
  and (_06487_, _06486_, _34796_);
  or (_06488_, _06487_, _06483_);
  or (_06489_, _06488_, _34790_);
  and (_06490_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_06491_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_06492_, _06491_, _06490_);
  and (_06493_, _06492_, _34581_);
  and (_06494_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_06495_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_06496_, _06495_, _06494_);
  and (_06497_, _06496_, _34796_);
  or (_06498_, _06497_, _06493_);
  or (_06499_, _06498_, _34772_);
  and (_06500_, _06499_, _34803_);
  and (_06501_, _06500_, _06489_);
  or (_06502_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_06503_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_06504_, _06503_, _34796_);
  and (_06505_, _06504_, _06502_);
  or (_06506_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_06507_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_06508_, _06507_, _34581_);
  and (_06509_, _06508_, _06506_);
  or (_06510_, _06509_, _06505_);
  or (_06511_, _06510_, _34790_);
  or (_06512_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_06513_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_06514_, _06513_, _34796_);
  and (_06515_, _06514_, _06512_);
  or (_06516_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_06517_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_06518_, _06517_, _34581_);
  and (_06519_, _06518_, _06516_);
  or (_06520_, _06519_, _06515_);
  or (_06521_, _06520_, _34772_);
  and (_06522_, _06521_, _34719_);
  and (_06523_, _06522_, _06511_);
  or (_06524_, _06523_, _06501_);
  and (_06525_, _06524_, _34789_);
  and (_06526_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_06527_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_06528_, _06527_, _06526_);
  and (_06529_, _06528_, _34581_);
  and (_06530_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_06531_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_06532_, _06531_, _06530_);
  and (_06533_, _06532_, _34796_);
  or (_06534_, _06533_, _06529_);
  or (_06535_, _06534_, _34790_);
  and (_06536_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_06537_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_06538_, _06537_, _06536_);
  and (_06539_, _06538_, _34581_);
  and (_06540_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_06541_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_06542_, _06541_, _06540_);
  and (_06543_, _06542_, _34796_);
  or (_06544_, _06543_, _06539_);
  or (_06545_, _06544_, _34772_);
  and (_06546_, _06545_, _34803_);
  and (_06547_, _06546_, _06535_);
  or (_06548_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_06549_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_06550_, _06549_, _06548_);
  and (_06551_, _06550_, _34581_);
  or (_06552_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_06553_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_06554_, _06553_, _06552_);
  and (_06555_, _06554_, _34796_);
  or (_06556_, _06555_, _06551_);
  or (_06557_, _06556_, _34790_);
  or (_06558_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_06559_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_06560_, _06559_, _06558_);
  and (_06561_, _06560_, _34581_);
  or (_06562_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_06563_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_06564_, _06563_, _06562_);
  and (_06565_, _06564_, _34796_);
  or (_06566_, _06565_, _06561_);
  or (_06567_, _06566_, _34772_);
  and (_06568_, _06567_, _34719_);
  and (_06569_, _06568_, _06557_);
  or (_06570_, _06569_, _06547_);
  and (_06571_, _06570_, _34700_);
  or (_06572_, _06571_, _06525_);
  and (_06573_, _06572_, _34840_);
  or (_06574_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_06575_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_06576_, _06575_, _06574_);
  and (_06577_, _06576_, _34581_);
  or (_06578_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_06579_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_06580_, _06579_, _06578_);
  and (_06581_, _06580_, _34796_);
  or (_06582_, _06581_, _06577_);
  and (_06583_, _06582_, _34790_);
  or (_06584_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_06585_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_06586_, _06585_, _06584_);
  and (_06587_, _06586_, _34581_);
  or (_06588_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_06589_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_06590_, _06589_, _06588_);
  and (_06591_, _06590_, _34796_);
  or (_06592_, _06591_, _06587_);
  and (_06593_, _06592_, _34772_);
  or (_06594_, _06593_, _06583_);
  and (_06595_, _06594_, _34719_);
  and (_06596_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_06597_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_06598_, _06597_, _06596_);
  and (_06599_, _06598_, _34581_);
  and (_06600_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_06601_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_06602_, _06601_, _06600_);
  and (_06603_, _06602_, _34796_);
  or (_06604_, _06603_, _06599_);
  and (_06605_, _06604_, _34790_);
  and (_06606_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_06607_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_06608_, _06607_, _06606_);
  and (_06609_, _06608_, _34581_);
  and (_06610_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_06611_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_06612_, _06611_, _06610_);
  and (_06613_, _06612_, _34796_);
  or (_06614_, _06613_, _06609_);
  and (_06615_, _06614_, _34772_);
  or (_06616_, _06615_, _06605_);
  and (_06617_, _06616_, _34803_);
  or (_06618_, _06617_, _06595_);
  and (_06619_, _06618_, _34700_);
  or (_06620_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_06621_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and (_06622_, _06621_, _34796_);
  and (_06623_, _06622_, _06620_);
  or (_06624_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_06625_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_06626_, _06625_, _34581_);
  and (_06627_, _06626_, _06624_);
  or (_06628_, _06627_, _06623_);
  and (_06629_, _06628_, _34790_);
  or (_06630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_06631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and (_06632_, _06631_, _34796_);
  and (_06633_, _06632_, _06630_);
  or (_06634_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_06635_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and (_06636_, _06635_, _34581_);
  and (_06637_, _06636_, _06634_);
  or (_06638_, _06637_, _06633_);
  and (_06639_, _06638_, _34772_);
  or (_06640_, _06639_, _06629_);
  and (_06641_, _06640_, _34719_);
  and (_06642_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and (_06643_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_06644_, _06643_, _06642_);
  and (_06645_, _06644_, _34581_);
  and (_06646_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and (_06647_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_06648_, _06647_, _06646_);
  and (_06649_, _06648_, _34796_);
  or (_06650_, _06649_, _06645_);
  and (_06651_, _06650_, _34790_);
  and (_06652_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_06653_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_06654_, _06653_, _06652_);
  and (_06655_, _06654_, _34581_);
  and (_06656_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and (_06657_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_06658_, _06657_, _06656_);
  and (_06659_, _06658_, _34796_);
  or (_06660_, _06659_, _06655_);
  and (_06661_, _06660_, _34772_);
  or (_06662_, _06661_, _06651_);
  and (_06663_, _06662_, _34803_);
  or (_06664_, _06663_, _06641_);
  and (_06665_, _06664_, _34789_);
  or (_06666_, _06665_, _06619_);
  and (_06667_, _06666_, _34638_);
  or (_06668_, _06667_, _06573_);
  or (_06669_, _06668_, _34985_);
  and (_06670_, _06669_, _06479_);
  or (_06671_, _06670_, _34346_);
  and (_06672_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_06673_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_06674_, _06673_, _06672_);
  and (_06675_, _06674_, _34796_);
  and (_06676_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_06677_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_06678_, _06677_, _06676_);
  and (_06679_, _06678_, _34581_);
  or (_06680_, _06679_, _06675_);
  or (_06681_, _06680_, _34790_);
  and (_06682_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_06683_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_06684_, _06683_, _06682_);
  and (_06685_, _06684_, _34796_);
  and (_06686_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_06687_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_06688_, _06687_, _06686_);
  and (_06689_, _06688_, _34581_);
  or (_06690_, _06689_, _06685_);
  or (_06691_, _06690_, _34772_);
  and (_06692_, _06691_, _34803_);
  and (_06693_, _06692_, _06681_);
  or (_06694_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_06695_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_06696_, _06695_, _34581_);
  and (_06697_, _06696_, _06694_);
  or (_06698_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_06699_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_06700_, _06699_, _34796_);
  and (_06701_, _06700_, _06698_);
  or (_06702_, _06701_, _06697_);
  or (_06703_, _06702_, _34790_);
  or (_06704_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_06705_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_06706_, _06705_, _34581_);
  and (_06707_, _06706_, _06704_);
  or (_06708_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_06709_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_06710_, _06709_, _34796_);
  and (_06711_, _06710_, _06708_);
  or (_06712_, _06711_, _06707_);
  or (_06713_, _06712_, _34772_);
  and (_06714_, _06713_, _34719_);
  and (_06715_, _06714_, _06703_);
  or (_06716_, _06715_, _06693_);
  and (_06717_, _06716_, _34789_);
  and (_06718_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_06719_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_06720_, _06719_, _34581_);
  or (_06721_, _06720_, _06718_);
  and (_06722_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_06723_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_06724_, _06723_, _34796_);
  or (_06725_, _06724_, _06722_);
  and (_06726_, _06725_, _06721_);
  or (_06727_, _06726_, _34790_);
  and (_06728_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_06729_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_06730_, _06729_, _34581_);
  or (_06731_, _06730_, _06728_);
  and (_06732_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_06733_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_06734_, _06733_, _34796_);
  or (_06735_, _06734_, _06732_);
  and (_06736_, _06735_, _06731_);
  or (_06737_, _06736_, _34772_);
  and (_06738_, _06737_, _34803_);
  and (_06739_, _06738_, _06727_);
  or (_06740_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_06741_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_06742_, _06741_, _06740_);
  or (_06743_, _06742_, _34796_);
  or (_06744_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_06745_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_06746_, _06745_, _06744_);
  or (_06747_, _06746_, _34581_);
  and (_06748_, _06747_, _06743_);
  or (_06749_, _06748_, _34790_);
  or (_06750_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_06751_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_06752_, _06751_, _06750_);
  or (_06753_, _06752_, _34796_);
  or (_06754_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_06755_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_06756_, _06755_, _06754_);
  or (_06757_, _06756_, _34581_);
  and (_06758_, _06757_, _06753_);
  or (_06759_, _06758_, _34772_);
  and (_06760_, _06759_, _34719_);
  and (_06761_, _06760_, _06749_);
  or (_06762_, _06761_, _06739_);
  and (_06763_, _06762_, _34700_);
  or (_06764_, _06763_, _06717_);
  and (_06765_, _06764_, _34840_);
  and (_06766_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and (_06767_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_06768_, _06767_, _06766_);
  and (_06769_, _06768_, _34581_);
  and (_06770_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  and (_06771_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or (_06772_, _06771_, _06770_);
  and (_06773_, _06772_, _34796_);
  or (_06774_, _06773_, _06769_);
  and (_06775_, _06774_, _34772_);
  and (_06776_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and (_06777_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_06778_, _06777_, _06776_);
  and (_06779_, _06778_, _34581_);
  and (_06780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and (_06781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or (_06782_, _06781_, _06780_);
  and (_06783_, _06782_, _34796_);
  or (_06784_, _06783_, _06779_);
  and (_06785_, _06784_, _34790_);
  or (_06786_, _06785_, _06775_);
  and (_06787_, _06786_, _34803_);
  or (_06788_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or (_06789_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  and (_06790_, _06789_, _06788_);
  and (_06791_, _06790_, _34581_);
  or (_06792_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or (_06793_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and (_06794_, _06793_, _06792_);
  and (_06795_, _06794_, _34796_);
  or (_06796_, _06795_, _06791_);
  and (_06797_, _06796_, _34772_);
  or (_06798_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_06799_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and (_06800_, _06799_, _06798_);
  and (_06801_, _06800_, _34581_);
  or (_06802_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_06803_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and (_06804_, _06803_, _06802_);
  and (_06805_, _06804_, _34796_);
  or (_06806_, _06805_, _06801_);
  and (_06807_, _06806_, _34790_);
  or (_06808_, _06807_, _06797_);
  and (_06809_, _06808_, _34719_);
  or (_06810_, _06809_, _06787_);
  and (_06811_, _06810_, _34789_);
  and (_06812_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_06813_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_06814_, _06813_, _06812_);
  and (_06815_, _06814_, _34581_);
  and (_06816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_06817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_06818_, _06817_, _06816_);
  and (_06819_, _06818_, _34796_);
  or (_06820_, _06819_, _06815_);
  and (_06821_, _06820_, _34772_);
  and (_06822_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_06823_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_06824_, _06823_, _06822_);
  and (_06825_, _06824_, _34581_);
  and (_06826_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_06827_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_06828_, _06827_, _06826_);
  and (_06829_, _06828_, _34796_);
  or (_06830_, _06829_, _06825_);
  and (_06831_, _06830_, _34790_);
  or (_06832_, _06831_, _06821_);
  and (_06833_, _06832_, _34803_);
  or (_06834_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_06835_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_06836_, _06835_, _06834_);
  and (_06837_, _06836_, _34581_);
  or (_06838_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_06839_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_06840_, _06839_, _06838_);
  and (_06841_, _06840_, _34796_);
  or (_06842_, _06841_, _06837_);
  and (_06843_, _06842_, _34772_);
  or (_06844_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_06845_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_06846_, _06845_, _06844_);
  and (_06847_, _06846_, _34581_);
  or (_06848_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_06849_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_06850_, _06849_, _06848_);
  and (_06851_, _06850_, _34796_);
  or (_06852_, _06851_, _06847_);
  and (_06853_, _06852_, _34790_);
  or (_06854_, _06853_, _06843_);
  and (_06855_, _06854_, _34719_);
  or (_06856_, _06855_, _06833_);
  and (_06857_, _06856_, _34700_);
  or (_06858_, _06857_, _06811_);
  and (_06859_, _06858_, _34638_);
  or (_06860_, _06859_, _06765_);
  or (_06861_, _06860_, _34692_);
  and (_06862_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_06863_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_06864_, _06863_, _06862_);
  and (_06865_, _06864_, _34581_);
  and (_06866_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_06867_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_06868_, _06867_, _06866_);
  and (_06869_, _06868_, _34796_);
  or (_06870_, _06869_, _06865_);
  or (_06871_, _06870_, _34790_);
  and (_06872_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_06873_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_06874_, _06873_, _06872_);
  and (_06875_, _06874_, _34581_);
  and (_06876_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_06877_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_06878_, _06877_, _06876_);
  and (_06879_, _06878_, _34796_);
  or (_06880_, _06879_, _06875_);
  or (_06881_, _06880_, _34772_);
  and (_06882_, _06881_, _34803_);
  and (_06883_, _06882_, _06871_);
  or (_06884_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_06885_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_06886_, _06885_, _34796_);
  and (_06887_, _06886_, _06884_);
  or (_06888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_06889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_06890_, _06889_, _34581_);
  and (_06891_, _06890_, _06888_);
  or (_06892_, _06891_, _06887_);
  or (_06893_, _06892_, _34790_);
  or (_06894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_06895_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_06896_, _06895_, _34796_);
  and (_06897_, _06896_, _06894_);
  or (_06898_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_06899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_06900_, _06899_, _34581_);
  and (_06901_, _06900_, _06898_);
  or (_06902_, _06901_, _06897_);
  or (_06903_, _06902_, _34772_);
  and (_06904_, _06903_, _34719_);
  and (_06905_, _06904_, _06893_);
  or (_06906_, _06905_, _06883_);
  and (_06907_, _06906_, _34789_);
  and (_06908_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_06909_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_06910_, _06909_, _06908_);
  and (_06911_, _06910_, _34581_);
  and (_06912_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_06913_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_06914_, _06913_, _06912_);
  and (_06915_, _06914_, _34796_);
  or (_06916_, _06915_, _06911_);
  or (_06917_, _06916_, _34790_);
  and (_06918_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_06919_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_06920_, _06919_, _06918_);
  and (_06921_, _06920_, _34581_);
  and (_06922_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_06923_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_06924_, _06923_, _06922_);
  and (_06925_, _06924_, _34796_);
  or (_06926_, _06925_, _06921_);
  or (_06927_, _06926_, _34772_);
  and (_06928_, _06927_, _34803_);
  and (_06929_, _06928_, _06917_);
  or (_06930_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_06931_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_06932_, _06931_, _06930_);
  and (_06933_, _06932_, _34581_);
  or (_06934_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_06935_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_06936_, _06935_, _06934_);
  and (_06937_, _06936_, _34796_);
  or (_06938_, _06937_, _06933_);
  or (_06939_, _06938_, _34790_);
  or (_06940_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_06941_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_06942_, _06941_, _06940_);
  and (_06943_, _06942_, _34581_);
  or (_06944_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_06945_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_06946_, _06945_, _06944_);
  and (_06947_, _06946_, _34796_);
  or (_06948_, _06947_, _06943_);
  or (_06949_, _06948_, _34772_);
  and (_06950_, _06949_, _34719_);
  and (_06951_, _06950_, _06939_);
  or (_06952_, _06951_, _06929_);
  and (_06953_, _06952_, _34700_);
  or (_06954_, _06953_, _06907_);
  and (_06955_, _06954_, _34840_);
  or (_06956_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_06957_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_06958_, _06957_, _06956_);
  and (_06959_, _06958_, _34581_);
  or (_06960_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_06961_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_06962_, _06961_, _06960_);
  and (_06963_, _06962_, _34796_);
  or (_06964_, _06963_, _06959_);
  and (_06965_, _06964_, _34790_);
  or (_06966_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_06967_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_06968_, _06967_, _06966_);
  and (_06969_, _06968_, _34581_);
  or (_06970_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_06971_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_06972_, _06971_, _06970_);
  and (_06973_, _06972_, _34796_);
  or (_06974_, _06973_, _06969_);
  and (_06975_, _06974_, _34772_);
  or (_06976_, _06975_, _06965_);
  and (_06977_, _06976_, _34719_);
  and (_06978_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_06979_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_06980_, _06979_, _06978_);
  and (_06981_, _06980_, _34581_);
  and (_06982_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_06983_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_06984_, _06983_, _06982_);
  and (_06985_, _06984_, _34796_);
  or (_06986_, _06985_, _06981_);
  and (_06987_, _06986_, _34790_);
  and (_06988_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_06989_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_06990_, _06989_, _06988_);
  and (_06991_, _06990_, _34581_);
  and (_06992_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_06993_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_06994_, _06993_, _06992_);
  and (_06995_, _06994_, _34796_);
  or (_06996_, _06995_, _06991_);
  and (_06997_, _06996_, _34772_);
  or (_06998_, _06997_, _06987_);
  and (_06999_, _06998_, _34803_);
  or (_07000_, _06999_, _06977_);
  and (_07001_, _07000_, _34700_);
  or (_07002_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_07003_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_07004_, _07003_, _34796_);
  and (_07005_, _07004_, _07002_);
  or (_07006_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_07007_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_07008_, _07007_, _34581_);
  and (_07009_, _07008_, _07006_);
  or (_07010_, _07009_, _07005_);
  and (_07011_, _07010_, _34790_);
  or (_07012_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_07013_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_07014_, _07013_, _34796_);
  and (_07015_, _07014_, _07012_);
  or (_07016_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_07017_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_07018_, _07017_, _34581_);
  and (_07019_, _07018_, _07016_);
  or (_07020_, _07019_, _07015_);
  and (_07021_, _07020_, _34772_);
  or (_07022_, _07021_, _07011_);
  and (_07023_, _07022_, _34719_);
  and (_07024_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_07025_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_07026_, _07025_, _07024_);
  and (_07027_, _07026_, _34581_);
  and (_07028_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_07029_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_07030_, _07029_, _07028_);
  and (_07031_, _07030_, _34796_);
  or (_07032_, _07031_, _07027_);
  and (_07033_, _07032_, _34790_);
  and (_07034_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_07035_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_07036_, _07035_, _07034_);
  and (_07037_, _07036_, _34581_);
  and (_07038_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_07039_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_07040_, _07039_, _07038_);
  and (_07041_, _07040_, _34796_);
  or (_07042_, _07041_, _07037_);
  and (_07043_, _07042_, _34772_);
  or (_07044_, _07043_, _07033_);
  and (_07045_, _07044_, _34803_);
  or (_07046_, _07045_, _07023_);
  and (_07047_, _07046_, _34789_);
  or (_07048_, _07047_, _07001_);
  and (_07049_, _07048_, _34638_);
  or (_07050_, _07049_, _06955_);
  or (_07051_, _07050_, _34985_);
  and (_07052_, _07051_, _06861_);
  or (_07053_, _07052_, _35178_);
  and (_07054_, _07053_, _06671_);
  or (_07055_, _07054_, _34788_);
  or (_07056_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_07057_, _07056_, _38997_);
  and (_38984_[1], _07057_, _07055_);
  and (_07058_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_07059_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_07060_, _07059_, _07058_);
  and (_07061_, _07060_, _34581_);
  and (_07062_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_07063_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_07064_, _07063_, _07062_);
  and (_07065_, _07064_, _34796_);
  or (_07066_, _07065_, _07061_);
  or (_07067_, _07066_, _34790_);
  and (_07068_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_07069_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_07070_, _07069_, _07068_);
  and (_07071_, _07070_, _34581_);
  and (_07072_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_07073_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_07074_, _07073_, _07072_);
  and (_07075_, _07074_, _34796_);
  or (_07076_, _07075_, _07071_);
  or (_07077_, _07076_, _34772_);
  and (_07078_, _07077_, _34803_);
  and (_07079_, _07078_, _07067_);
  or (_07080_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_07081_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_07082_, _07081_, _07080_);
  and (_07083_, _07082_, _34581_);
  or (_07084_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_07085_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_07086_, _07085_, _07084_);
  and (_07087_, _07086_, _34796_);
  or (_07088_, _07087_, _07083_);
  or (_07089_, _07088_, _34790_);
  or (_07090_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_07091_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_07092_, _07091_, _07090_);
  and (_07093_, _07092_, _34581_);
  or (_07094_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_07095_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_07096_, _07095_, _07094_);
  and (_07097_, _07096_, _34796_);
  or (_07098_, _07097_, _07093_);
  or (_07099_, _07098_, _34772_);
  and (_07100_, _07099_, _34719_);
  and (_07101_, _07100_, _07089_);
  or (_07102_, _07101_, _07079_);
  and (_07103_, _07102_, _34700_);
  and (_07104_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_07105_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_07106_, _07105_, _07104_);
  and (_07107_, _07106_, _34581_);
  and (_07108_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_07109_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_07110_, _07109_, _07108_);
  and (_07111_, _07110_, _34796_);
  or (_07112_, _07111_, _07107_);
  or (_07113_, _07112_, _34790_);
  and (_07114_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_07115_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_07116_, _07115_, _07114_);
  and (_07117_, _07116_, _34581_);
  and (_07118_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_07119_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_07120_, _07119_, _07118_);
  and (_07121_, _07120_, _34796_);
  or (_07122_, _07121_, _07117_);
  or (_07123_, _07122_, _34772_);
  and (_07124_, _07123_, _34803_);
  and (_07125_, _07124_, _07113_);
  or (_07126_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_07127_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_07128_, _07127_, _34796_);
  and (_07129_, _07128_, _07126_);
  or (_07130_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_07131_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_07132_, _07131_, _34581_);
  and (_07133_, _07132_, _07130_);
  or (_07134_, _07133_, _07129_);
  or (_07135_, _07134_, _34790_);
  or (_07136_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_07137_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_07138_, _07137_, _34796_);
  and (_07139_, _07138_, _07136_);
  or (_07140_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_07141_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_07142_, _07141_, _34581_);
  and (_07143_, _07142_, _07140_);
  or (_07144_, _07143_, _07139_);
  or (_07145_, _07144_, _34772_);
  and (_07146_, _07145_, _34719_);
  and (_07147_, _07146_, _07135_);
  or (_07148_, _07147_, _07125_);
  and (_07149_, _07148_, _34789_);
  or (_07150_, _07149_, _07103_);
  and (_07151_, _07150_, _34840_);
  and (_07152_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_07153_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_07154_, _07153_, _07152_);
  and (_07155_, _07154_, _34581_);
  and (_07156_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_07157_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_07158_, _07157_, _07156_);
  and (_07159_, _07158_, _34796_);
  or (_07160_, _07159_, _07155_);
  and (_07161_, _07160_, _34772_);
  and (_07162_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_07163_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_07164_, _07163_, _07162_);
  and (_07165_, _07164_, _34581_);
  and (_07166_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_07167_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_07168_, _07167_, _07166_);
  and (_07169_, _07168_, _34796_);
  or (_07170_, _07169_, _07165_);
  and (_07171_, _07170_, _34790_);
  or (_07172_, _07171_, _07161_);
  and (_07173_, _07172_, _34803_);
  or (_07174_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_07175_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_07176_, _07175_, _34796_);
  and (_07177_, _07176_, _07174_);
  or (_07178_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_07179_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_07180_, _07179_, _34581_);
  and (_07181_, _07180_, _07178_);
  or (_07182_, _07181_, _07177_);
  and (_07183_, _07182_, _34772_);
  or (_07184_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_07185_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_07186_, _07185_, _34796_);
  and (_07187_, _07186_, _07184_);
  or (_07188_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_07189_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_07190_, _07189_, _34581_);
  and (_07191_, _07190_, _07188_);
  or (_07192_, _07191_, _07187_);
  and (_07193_, _07192_, _34790_);
  or (_07194_, _07193_, _07183_);
  and (_07195_, _07194_, _34719_);
  or (_07196_, _07195_, _07173_);
  and (_07197_, _07196_, _34789_);
  and (_07198_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_07199_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_07200_, _07199_, _07198_);
  and (_07201_, _07200_, _34581_);
  and (_07202_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_07203_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_07204_, _07203_, _07202_);
  and (_07205_, _07204_, _34796_);
  or (_07206_, _07205_, _07201_);
  and (_07207_, _07206_, _34772_);
  and (_07208_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_07209_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_07210_, _07209_, _07208_);
  and (_07211_, _07210_, _34581_);
  and (_07212_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_07213_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_07214_, _07213_, _07212_);
  and (_07215_, _07214_, _34796_);
  or (_07216_, _07215_, _07211_);
  and (_07217_, _07216_, _34790_);
  or (_07218_, _07217_, _07207_);
  and (_07219_, _07218_, _34803_);
  or (_07220_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_07221_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_07222_, _07221_, _07220_);
  and (_07223_, _07222_, _34581_);
  or (_07224_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_07225_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_07226_, _07225_, _07224_);
  and (_07227_, _07226_, _34796_);
  or (_07228_, _07227_, _07223_);
  and (_07229_, _07228_, _34772_);
  or (_07230_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_07231_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_07232_, _07231_, _07230_);
  and (_07233_, _07232_, _34581_);
  or (_07234_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_07235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_07236_, _07235_, _07234_);
  and (_07237_, _07236_, _34796_);
  or (_07238_, _07237_, _07233_);
  and (_07239_, _07238_, _34790_);
  or (_07240_, _07239_, _07229_);
  and (_07241_, _07240_, _34719_);
  or (_07242_, _07241_, _07219_);
  and (_07243_, _07242_, _34700_);
  or (_07244_, _07243_, _07197_);
  and (_07245_, _07244_, _34638_);
  or (_07246_, _07245_, _07151_);
  or (_07247_, _07246_, _34692_);
  and (_07248_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_07249_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_07250_, _07249_, _07248_);
  and (_07251_, _07250_, _34581_);
  and (_07252_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_07253_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_07254_, _07253_, _07252_);
  and (_07255_, _07254_, _34796_);
  or (_07256_, _07255_, _07251_);
  or (_07257_, _07256_, _34790_);
  and (_07258_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_07259_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_07260_, _07259_, _07258_);
  and (_07261_, _07260_, _34581_);
  and (_07262_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_07263_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_07264_, _07263_, _07262_);
  and (_07265_, _07264_, _34796_);
  or (_07266_, _07265_, _07261_);
  or (_07267_, _07266_, _34772_);
  and (_07268_, _07267_, _34803_);
  and (_07269_, _07268_, _07257_);
  or (_07270_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_07271_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_07272_, _07271_, _34796_);
  and (_07273_, _07272_, _07270_);
  or (_07274_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_07275_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_07276_, _07275_, _34581_);
  and (_07277_, _07276_, _07274_);
  or (_07278_, _07277_, _07273_);
  or (_07279_, _07278_, _34790_);
  or (_07280_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_07281_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_07282_, _07281_, _34796_);
  and (_07283_, _07282_, _07280_);
  or (_07284_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_07285_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_07286_, _07285_, _34581_);
  and (_07287_, _07286_, _07284_);
  or (_07288_, _07287_, _07283_);
  or (_07289_, _07288_, _34772_);
  and (_07290_, _07289_, _34719_);
  and (_07291_, _07290_, _07279_);
  or (_07292_, _07291_, _07269_);
  and (_07293_, _07292_, _34789_);
  and (_07294_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_07295_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_07296_, _07295_, _07294_);
  and (_07297_, _07296_, _34581_);
  and (_07298_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_07299_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_07300_, _07299_, _07298_);
  and (_07301_, _07300_, _34796_);
  or (_07302_, _07301_, _07297_);
  or (_07303_, _07302_, _34790_);
  and (_07304_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_07305_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_07306_, _07305_, _07304_);
  and (_07307_, _07306_, _34581_);
  and (_07308_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_07309_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_07310_, _07309_, _07308_);
  and (_07311_, _07310_, _34796_);
  or (_07312_, _07311_, _07307_);
  or (_07313_, _07312_, _34772_);
  and (_07314_, _07313_, _34803_);
  and (_07315_, _07314_, _07303_);
  or (_07316_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_07317_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_07318_, _07317_, _07316_);
  and (_07319_, _07318_, _34581_);
  or (_07320_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_07321_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_07322_, _07321_, _07320_);
  and (_07323_, _07322_, _34796_);
  or (_07324_, _07323_, _07319_);
  or (_07325_, _07324_, _34790_);
  or (_07326_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_07327_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_07328_, _07327_, _07326_);
  and (_07329_, _07328_, _34581_);
  or (_07330_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_07331_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_07332_, _07331_, _07330_);
  and (_07333_, _07332_, _34796_);
  or (_07334_, _07333_, _07329_);
  or (_07335_, _07334_, _34772_);
  and (_07336_, _07335_, _34719_);
  and (_07337_, _07336_, _07325_);
  or (_07338_, _07337_, _07315_);
  and (_07339_, _07338_, _34700_);
  or (_07340_, _07339_, _07293_);
  and (_07341_, _07340_, _34840_);
  or (_07342_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_07343_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_07344_, _07343_, _07342_);
  and (_07345_, _07344_, _34581_);
  or (_07346_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_07347_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_07348_, _07347_, _07346_);
  and (_07349_, _07348_, _34796_);
  or (_07350_, _07349_, _07345_);
  and (_07351_, _07350_, _34790_);
  or (_07352_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_07353_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_07354_, _07353_, _07352_);
  and (_07355_, _07354_, _34581_);
  or (_07356_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_07357_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_07358_, _07357_, _07356_);
  and (_07359_, _07358_, _34796_);
  or (_07360_, _07359_, _07355_);
  and (_07361_, _07360_, _34772_);
  or (_07362_, _07361_, _07351_);
  and (_07363_, _07362_, _34719_);
  and (_07364_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_07365_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_07366_, _07365_, _07364_);
  and (_07367_, _07366_, _34581_);
  and (_07368_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_07369_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_07370_, _07369_, _07368_);
  and (_07371_, _07370_, _34796_);
  or (_07372_, _07371_, _07367_);
  and (_07373_, _07372_, _34790_);
  and (_07374_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_07375_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_07376_, _07375_, _07374_);
  and (_07377_, _07376_, _34581_);
  and (_07378_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_07379_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_07380_, _07379_, _07378_);
  and (_07381_, _07380_, _34796_);
  or (_07382_, _07381_, _07377_);
  and (_07383_, _07382_, _34772_);
  or (_07384_, _07383_, _07373_);
  and (_07385_, _07384_, _34803_);
  or (_07386_, _07385_, _07363_);
  and (_07387_, _07386_, _34700_);
  or (_07388_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_07389_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_07390_, _07389_, _34796_);
  and (_07391_, _07390_, _07388_);
  or (_07392_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_07393_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_07394_, _07393_, _34581_);
  and (_07395_, _07394_, _07392_);
  or (_07396_, _07395_, _07391_);
  and (_07397_, _07396_, _34790_);
  or (_07398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_07399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  and (_07400_, _07399_, _34796_);
  and (_07401_, _07400_, _07398_);
  or (_07402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_07403_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_07404_, _07403_, _34581_);
  and (_07405_, _07404_, _07402_);
  or (_07406_, _07405_, _07401_);
  and (_07407_, _07406_, _34772_);
  or (_07408_, _07407_, _07397_);
  and (_07409_, _07408_, _34719_);
  and (_07410_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_07411_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_07412_, _07411_, _07410_);
  and (_07413_, _07412_, _34581_);
  and (_07414_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  and (_07415_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_07416_, _07415_, _07414_);
  and (_07417_, _07416_, _34796_);
  or (_07418_, _07417_, _07413_);
  and (_07419_, _07418_, _34790_);
  and (_07420_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  and (_07421_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_07422_, _07421_, _07420_);
  and (_07423_, _07422_, _34581_);
  and (_07424_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_07425_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_07426_, _07425_, _07424_);
  and (_07427_, _07426_, _34796_);
  or (_07428_, _07427_, _07423_);
  and (_07429_, _07428_, _34772_);
  or (_07430_, _07429_, _07419_);
  and (_07431_, _07430_, _34803_);
  or (_07432_, _07431_, _07409_);
  and (_07433_, _07432_, _34789_);
  or (_07434_, _07433_, _07387_);
  and (_07435_, _07434_, _34638_);
  or (_07436_, _07435_, _07341_);
  or (_07437_, _07436_, _34985_);
  and (_07438_, _07437_, _07247_);
  or (_07439_, _07438_, _34346_);
  and (_07440_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_07441_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_07442_, _07441_, _07440_);
  and (_07443_, _07442_, _34796_);
  and (_07444_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_07445_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_07446_, _07445_, _07444_);
  and (_07447_, _07446_, _34581_);
  or (_07448_, _07447_, _07443_);
  or (_07449_, _07448_, _34790_);
  and (_07450_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_07451_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_07452_, _07451_, _07450_);
  and (_07453_, _07452_, _34796_);
  and (_07454_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_07455_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_07456_, _07455_, _07454_);
  and (_07457_, _07456_, _34581_);
  or (_07458_, _07457_, _07453_);
  or (_07459_, _07458_, _34772_);
  and (_07460_, _07459_, _34803_);
  and (_07461_, _07460_, _07449_);
  or (_07462_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_07463_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_07464_, _07463_, _34581_);
  and (_07465_, _07464_, _07462_);
  or (_07466_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_07467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_07468_, _07467_, _34796_);
  and (_07469_, _07468_, _07466_);
  or (_07470_, _07469_, _07465_);
  or (_07471_, _07470_, _34790_);
  or (_07472_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_07473_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_07474_, _07473_, _34581_);
  and (_07475_, _07474_, _07472_);
  or (_07476_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_07477_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_07478_, _07477_, _34796_);
  and (_07479_, _07478_, _07476_);
  or (_07480_, _07479_, _07475_);
  or (_07481_, _07480_, _34772_);
  and (_07482_, _07481_, _34719_);
  and (_07483_, _07482_, _07471_);
  or (_07484_, _07483_, _07461_);
  and (_07485_, _07484_, _34789_);
  and (_07486_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_07487_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_07488_, _07487_, _34581_);
  or (_07489_, _07488_, _07486_);
  and (_07490_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_07491_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_07492_, _07491_, _34796_);
  or (_07493_, _07492_, _07490_);
  and (_07494_, _07493_, _07489_);
  or (_07495_, _07494_, _34790_);
  and (_07496_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_07497_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_07498_, _07497_, _34581_);
  or (_07499_, _07498_, _07496_);
  and (_07500_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_07501_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_07502_, _07501_, _34796_);
  or (_07503_, _07502_, _07500_);
  and (_07504_, _07503_, _07499_);
  or (_07505_, _07504_, _34772_);
  and (_07506_, _07505_, _34803_);
  and (_07507_, _07506_, _07495_);
  or (_07508_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_07509_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_07510_, _07509_, _07508_);
  or (_07511_, _07510_, _34796_);
  or (_07512_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_07513_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_07514_, _07513_, _07512_);
  or (_07515_, _07514_, _34581_);
  and (_07516_, _07515_, _07511_);
  or (_07517_, _07516_, _34790_);
  or (_07518_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_07519_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_07520_, _07519_, _07518_);
  or (_07521_, _07520_, _34796_);
  or (_07522_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_07523_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_07524_, _07523_, _07522_);
  or (_07525_, _07524_, _34581_);
  and (_07526_, _07525_, _07521_);
  or (_07527_, _07526_, _34772_);
  and (_07528_, _07527_, _34719_);
  and (_07529_, _07528_, _07517_);
  or (_07530_, _07529_, _07507_);
  and (_07531_, _07530_, _34700_);
  or (_07532_, _07531_, _07485_);
  and (_07533_, _07532_, _34840_);
  and (_07534_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and (_07535_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_07536_, _07535_, _07534_);
  and (_07537_, _07536_, _34581_);
  and (_07538_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and (_07539_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or (_07540_, _07539_, _07538_);
  and (_07541_, _07540_, _34796_);
  or (_07542_, _07541_, _07537_);
  and (_07543_, _07542_, _34772_);
  and (_07544_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and (_07545_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_07546_, _07545_, _07544_);
  and (_07547_, _07546_, _34581_);
  and (_07548_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and (_07549_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or (_07550_, _07549_, _07548_);
  and (_07551_, _07550_, _34796_);
  or (_07552_, _07551_, _07547_);
  and (_07553_, _07552_, _34790_);
  or (_07554_, _07553_, _07543_);
  and (_07555_, _07554_, _34803_);
  or (_07556_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_07557_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  and (_07558_, _07557_, _07556_);
  and (_07559_, _07558_, _34581_);
  or (_07560_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_07561_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and (_07562_, _07561_, _07560_);
  and (_07563_, _07562_, _34796_);
  or (_07564_, _07563_, _07559_);
  and (_07565_, _07564_, _34772_);
  or (_07566_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or (_07567_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and (_07568_, _07567_, _07566_);
  and (_07569_, _07568_, _34581_);
  or (_07570_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_07571_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and (_07572_, _07571_, _07570_);
  and (_07573_, _07572_, _34796_);
  or (_07574_, _07573_, _07569_);
  and (_07575_, _07574_, _34790_);
  or (_07576_, _07575_, _07565_);
  and (_07577_, _07576_, _34719_);
  or (_07578_, _07577_, _07555_);
  and (_07579_, _07578_, _34789_);
  and (_07580_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_07581_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_07582_, _07581_, _07580_);
  and (_07583_, _07582_, _34581_);
  and (_07584_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_07585_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_07586_, _07585_, _07584_);
  and (_07587_, _07586_, _34796_);
  or (_07588_, _07587_, _07583_);
  and (_07589_, _07588_, _34772_);
  and (_07590_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_07591_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_07592_, _07591_, _07590_);
  and (_07593_, _07592_, _34581_);
  and (_07594_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_07595_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_07596_, _07595_, _07594_);
  and (_07597_, _07596_, _34796_);
  or (_07598_, _07597_, _07593_);
  and (_07599_, _07598_, _34790_);
  or (_07600_, _07599_, _07589_);
  and (_07601_, _07600_, _34803_);
  or (_07602_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_07603_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_07604_, _07603_, _07602_);
  and (_07605_, _07604_, _34581_);
  or (_07606_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_07607_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_07608_, _07607_, _07606_);
  and (_07609_, _07608_, _34796_);
  or (_07610_, _07609_, _07605_);
  and (_07611_, _07610_, _34772_);
  or (_07612_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_07613_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_07614_, _07613_, _07612_);
  and (_07615_, _07614_, _34581_);
  or (_07616_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_07617_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_07618_, _07617_, _07616_);
  and (_07619_, _07618_, _34796_);
  or (_07620_, _07619_, _07615_);
  and (_07621_, _07620_, _34790_);
  or (_07622_, _07621_, _07611_);
  and (_07623_, _07622_, _34719_);
  or (_07624_, _07623_, _07601_);
  and (_07625_, _07624_, _34700_);
  or (_07626_, _07625_, _07579_);
  and (_07627_, _07626_, _34638_);
  or (_07628_, _07627_, _07533_);
  or (_07629_, _07628_, _34692_);
  and (_07630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_07631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_07632_, _07631_, _07630_);
  and (_07633_, _07632_, _34581_);
  and (_07634_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_07635_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_07636_, _07635_, _07634_);
  and (_07637_, _07636_, _34796_);
  or (_07638_, _07637_, _07633_);
  or (_07639_, _07638_, _34790_);
  and (_07640_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_07641_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_07642_, _07641_, _07640_);
  and (_07643_, _07642_, _34581_);
  and (_07644_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_07645_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_07646_, _07645_, _07644_);
  and (_07647_, _07646_, _34796_);
  or (_07648_, _07647_, _07643_);
  or (_07649_, _07648_, _34772_);
  and (_07650_, _07649_, _34803_);
  and (_07651_, _07650_, _07639_);
  or (_07652_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_07653_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_07654_, _07653_, _34796_);
  and (_07655_, _07654_, _07652_);
  or (_07656_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_07657_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_07658_, _07657_, _34581_);
  and (_07659_, _07658_, _07656_);
  or (_07660_, _07659_, _07655_);
  or (_07661_, _07660_, _34790_);
  or (_07662_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_07663_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_07664_, _07663_, _34796_);
  and (_07665_, _07664_, _07662_);
  or (_07666_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_07667_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_07668_, _07667_, _34581_);
  and (_07669_, _07668_, _07666_);
  or (_07670_, _07669_, _07665_);
  or (_07671_, _07670_, _34772_);
  and (_07672_, _07671_, _34719_);
  and (_07673_, _07672_, _07661_);
  or (_07674_, _07673_, _07651_);
  and (_07675_, _07674_, _34789_);
  and (_07676_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_07677_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_07678_, _07677_, _07676_);
  and (_07679_, _07678_, _34581_);
  and (_07680_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_07681_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_07682_, _07681_, _07680_);
  and (_07683_, _07682_, _34796_);
  or (_07684_, _07683_, _07679_);
  or (_07685_, _07684_, _34790_);
  and (_07686_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_07687_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_07688_, _07687_, _07686_);
  and (_07689_, _07688_, _34581_);
  and (_07690_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_07691_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_07692_, _07691_, _07690_);
  and (_07693_, _07692_, _34796_);
  or (_07694_, _07693_, _07689_);
  or (_07695_, _07694_, _34772_);
  and (_07696_, _07695_, _34803_);
  and (_07697_, _07696_, _07685_);
  or (_07698_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_07699_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_07700_, _07699_, _07698_);
  and (_07701_, _07700_, _34581_);
  or (_07702_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_07703_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_07704_, _07703_, _07702_);
  and (_07705_, _07704_, _34796_);
  or (_07706_, _07705_, _07701_);
  or (_07707_, _07706_, _34790_);
  or (_07708_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_07709_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_07710_, _07709_, _07708_);
  and (_07711_, _07710_, _34581_);
  or (_07712_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_07713_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_07714_, _07713_, _07712_);
  and (_07715_, _07714_, _34796_);
  or (_07716_, _07715_, _07711_);
  or (_07717_, _07716_, _34772_);
  and (_07718_, _07717_, _34719_);
  and (_07719_, _07718_, _07707_);
  or (_07720_, _07719_, _07697_);
  and (_07721_, _07720_, _34700_);
  or (_07722_, _07721_, _07675_);
  and (_07723_, _07722_, _34840_);
  or (_07724_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_07725_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_07726_, _07725_, _07724_);
  and (_07727_, _07726_, _34581_);
  or (_07728_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_07729_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_07730_, _07729_, _07728_);
  and (_07731_, _07730_, _34796_);
  or (_07732_, _07731_, _07727_);
  and (_07733_, _07732_, _34790_);
  or (_07734_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_07735_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_07736_, _07735_, _07734_);
  and (_07737_, _07736_, _34581_);
  or (_07738_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_07739_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_07740_, _07739_, _07738_);
  and (_07741_, _07740_, _34796_);
  or (_07742_, _07741_, _07737_);
  and (_07743_, _07742_, _34772_);
  or (_07744_, _07743_, _07733_);
  and (_07745_, _07744_, _34719_);
  and (_07746_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_07747_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_07748_, _07747_, _07746_);
  and (_07749_, _07748_, _34581_);
  and (_07750_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_07751_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_07752_, _07751_, _07750_);
  and (_07753_, _07752_, _34796_);
  or (_07754_, _07753_, _07749_);
  and (_07755_, _07754_, _34790_);
  and (_07756_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_07757_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_07758_, _07757_, _07756_);
  and (_07759_, _07758_, _34581_);
  and (_07760_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_07761_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_07762_, _07761_, _07760_);
  and (_07763_, _07762_, _34796_);
  or (_07764_, _07763_, _07759_);
  and (_07765_, _07764_, _34772_);
  or (_07766_, _07765_, _07755_);
  and (_07767_, _07766_, _34803_);
  or (_07768_, _07767_, _07745_);
  and (_07769_, _07768_, _34700_);
  or (_07770_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_07771_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_07772_, _07771_, _34796_);
  and (_07773_, _07772_, _07770_);
  or (_07774_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_07775_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_07776_, _07775_, _34581_);
  and (_07777_, _07776_, _07774_);
  or (_07778_, _07777_, _07773_);
  and (_07779_, _07778_, _34790_);
  or (_07780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_07781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_07782_, _07781_, _34796_);
  and (_07783_, _07782_, _07780_);
  or (_07784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_07785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_07786_, _07785_, _34581_);
  and (_07787_, _07786_, _07784_);
  or (_07788_, _07787_, _07783_);
  and (_07789_, _07788_, _34772_);
  or (_07790_, _07789_, _07779_);
  and (_07791_, _07790_, _34719_);
  and (_07792_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_07793_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_07794_, _07793_, _07792_);
  and (_07795_, _07794_, _34581_);
  and (_07796_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_07797_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_07798_, _07797_, _07796_);
  and (_07799_, _07798_, _34796_);
  or (_07800_, _07799_, _07795_);
  and (_07801_, _07800_, _34790_);
  and (_07802_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_07803_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_07804_, _07803_, _07802_);
  and (_07805_, _07804_, _34581_);
  and (_07806_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_07807_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_07808_, _07807_, _07806_);
  and (_07809_, _07808_, _34796_);
  or (_07810_, _07809_, _07805_);
  and (_07811_, _07810_, _34772_);
  or (_07812_, _07811_, _07801_);
  and (_07813_, _07812_, _34803_);
  or (_07814_, _07813_, _07791_);
  and (_07815_, _07814_, _34789_);
  or (_07816_, _07815_, _07769_);
  and (_07817_, _07816_, _34638_);
  or (_07818_, _07817_, _07723_);
  or (_07819_, _07818_, _34985_);
  and (_07820_, _07819_, _07629_);
  or (_07821_, _07820_, _35178_);
  and (_07822_, _07821_, _07439_);
  or (_07823_, _07822_, _34788_);
  or (_07824_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_07825_, _07824_, _38997_);
  and (_38984_[2], _07825_, _07823_);
  and (_07826_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_07827_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_07828_, _07827_, _07826_);
  and (_07829_, _07828_, _34796_);
  and (_07830_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_07831_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_07832_, _07831_, _07830_);
  and (_07833_, _07832_, _34581_);
  or (_07834_, _07833_, _07829_);
  or (_07835_, _07834_, _34790_);
  and (_07836_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_07837_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_07838_, _07837_, _07836_);
  and (_07839_, _07838_, _34796_);
  and (_07840_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_07841_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_07842_, _07841_, _07840_);
  and (_07843_, _07842_, _34581_);
  or (_07844_, _07843_, _07839_);
  or (_07845_, _07844_, _34772_);
  and (_07846_, _07845_, _34803_);
  and (_07847_, _07846_, _07835_);
  or (_07848_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_07849_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_07850_, _07849_, _34581_);
  and (_07851_, _07850_, _07848_);
  or (_07852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_07853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_07854_, _07853_, _34796_);
  and (_07855_, _07854_, _07852_);
  or (_07856_, _07855_, _07851_);
  or (_07857_, _07856_, _34790_);
  or (_07858_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_07859_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_07860_, _07859_, _34581_);
  and (_07861_, _07860_, _07858_);
  or (_07862_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_07863_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_07864_, _07863_, _34796_);
  and (_07865_, _07864_, _07862_);
  or (_07866_, _07865_, _07861_);
  or (_07867_, _07866_, _34772_);
  and (_07868_, _07867_, _34719_);
  and (_07869_, _07868_, _07857_);
  or (_07870_, _07869_, _07847_);
  or (_07871_, _07870_, _34700_);
  and (_07872_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_07873_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_07874_, _07873_, _34581_);
  or (_07875_, _07874_, _07872_);
  and (_07876_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_07877_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_07878_, _07877_, _34796_);
  or (_07879_, _07878_, _07876_);
  and (_07880_, _07879_, _07875_);
  or (_07881_, _07880_, _34790_);
  and (_07882_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_07883_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_07884_, _07883_, _34581_);
  or (_07885_, _07884_, _07882_);
  and (_07886_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_07887_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_07888_, _07887_, _34796_);
  or (_07889_, _07888_, _07886_);
  and (_07890_, _07889_, _07885_);
  or (_07891_, _07890_, _34772_);
  and (_07892_, _07891_, _34803_);
  and (_07893_, _07892_, _07881_);
  or (_07894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_07895_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_07896_, _07895_, _07894_);
  or (_07897_, _07896_, _34796_);
  or (_07898_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_07899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_07900_, _07899_, _07898_);
  or (_07901_, _07900_, _34581_);
  and (_07902_, _07901_, _07897_);
  or (_07903_, _07902_, _34790_);
  or (_07904_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_07905_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_07906_, _07905_, _07904_);
  or (_07907_, _07906_, _34796_);
  or (_07908_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_07909_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_07910_, _07909_, _07908_);
  or (_07911_, _07910_, _34581_);
  and (_07912_, _07911_, _07907_);
  or (_07913_, _07912_, _34772_);
  and (_07914_, _07913_, _34719_);
  and (_07915_, _07914_, _07903_);
  or (_07916_, _07915_, _07893_);
  or (_07917_, _07916_, _34789_);
  and (_07918_, _07917_, _34840_);
  and (_07919_, _07918_, _07871_);
  and (_07920_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_07921_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_07922_, _07921_, _07920_);
  and (_07923_, _07922_, _34581_);
  and (_07924_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_07925_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_07926_, _07925_, _07924_);
  and (_07927_, _07926_, _34796_);
  or (_07928_, _07927_, _07923_);
  and (_07929_, _07928_, _34772_);
  and (_07930_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_07931_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_07932_, _07931_, _07930_);
  and (_07933_, _07932_, _34581_);
  and (_07934_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_07935_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_07936_, _07935_, _07934_);
  and (_07937_, _07936_, _34796_);
  or (_07938_, _07937_, _07933_);
  and (_07939_, _07938_, _34790_);
  or (_07940_, _07939_, _07929_);
  and (_07941_, _07940_, _34803_);
  or (_07942_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_07943_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_07944_, _07943_, _07942_);
  and (_07945_, _07944_, _34581_);
  or (_07946_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_07947_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_07948_, _07947_, _07946_);
  and (_07949_, _07948_, _34796_);
  or (_07950_, _07949_, _07945_);
  and (_07951_, _07950_, _34772_);
  or (_07952_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_07953_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_07954_, _07953_, _07952_);
  and (_07955_, _07954_, _34581_);
  or (_07956_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_07957_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_07958_, _07957_, _07956_);
  and (_07959_, _07958_, _34796_);
  or (_07960_, _07959_, _07955_);
  and (_07961_, _07960_, _34790_);
  or (_07962_, _07961_, _07951_);
  and (_07963_, _07962_, _34719_);
  or (_07964_, _07963_, _07941_);
  and (_07965_, _07964_, _34789_);
  and (_07966_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_07967_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_07968_, _07967_, _07966_);
  and (_07969_, _07968_, _34581_);
  and (_07970_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_07971_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_07972_, _07971_, _07970_);
  and (_07973_, _07972_, _34796_);
  or (_07974_, _07973_, _07969_);
  and (_07975_, _07974_, _34772_);
  and (_07976_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_07977_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_07978_, _07977_, _07976_);
  and (_07979_, _07978_, _34581_);
  and (_07980_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_07981_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_07982_, _07981_, _07980_);
  and (_07983_, _07982_, _34796_);
  or (_07984_, _07983_, _07979_);
  and (_07985_, _07984_, _34790_);
  or (_07986_, _07985_, _07975_);
  and (_07987_, _07986_, _34803_);
  or (_07988_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_07989_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_07990_, _07989_, _07988_);
  and (_07991_, _07990_, _34581_);
  or (_07992_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_07993_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_07994_, _07993_, _07992_);
  and (_07995_, _07994_, _34796_);
  or (_07996_, _07995_, _07991_);
  and (_07997_, _07996_, _34772_);
  or (_07998_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_07999_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_08000_, _07999_, _07998_);
  and (_08001_, _08000_, _34581_);
  or (_08002_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_08003_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_08004_, _08003_, _08002_);
  and (_08005_, _08004_, _34796_);
  or (_08006_, _08005_, _08001_);
  and (_08007_, _08006_, _34790_);
  or (_08008_, _08007_, _07997_);
  and (_08009_, _08008_, _34719_);
  or (_08010_, _08009_, _07987_);
  and (_08011_, _08010_, _34700_);
  or (_08012_, _08011_, _07965_);
  and (_08013_, _08012_, _34638_);
  or (_08014_, _08013_, _07919_);
  or (_08015_, _08014_, _34692_);
  and (_08016_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_08017_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_08018_, _08017_, _08016_);
  and (_08019_, _08018_, _34581_);
  and (_08020_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_08021_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_08022_, _08021_, _08020_);
  and (_08023_, _08022_, _34796_);
  or (_08024_, _08023_, _08019_);
  or (_08025_, _08024_, _34790_);
  and (_08026_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_08027_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_08028_, _08027_, _08026_);
  and (_08029_, _08028_, _34581_);
  and (_08030_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_08031_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_08032_, _08031_, _08030_);
  and (_08033_, _08032_, _34796_);
  or (_08034_, _08033_, _08029_);
  or (_08035_, _08034_, _34772_);
  and (_08036_, _08035_, _34803_);
  and (_08037_, _08036_, _08025_);
  or (_08038_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_08039_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_08040_, _08039_, _34796_);
  and (_08041_, _08040_, _08038_);
  or (_08042_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_08043_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_08044_, _08043_, _34581_);
  and (_08045_, _08044_, _08042_);
  or (_08046_, _08045_, _08041_);
  or (_08047_, _08046_, _34790_);
  or (_08048_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_08049_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_08050_, _08049_, _34796_);
  and (_08051_, _08050_, _08048_);
  or (_08052_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_08053_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_08054_, _08053_, _34581_);
  and (_08055_, _08054_, _08052_);
  or (_08056_, _08055_, _08051_);
  or (_08057_, _08056_, _34772_);
  and (_08058_, _08057_, _34719_);
  and (_08059_, _08058_, _08047_);
  or (_08060_, _08059_, _08037_);
  and (_08061_, _08060_, _34789_);
  and (_08062_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_08063_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_08064_, _08063_, _08062_);
  and (_08065_, _08064_, _34581_);
  and (_08066_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_08067_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_08068_, _08067_, _08066_);
  and (_08069_, _08068_, _34796_);
  or (_08070_, _08069_, _08065_);
  or (_08071_, _08070_, _34790_);
  and (_08072_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_08073_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_08074_, _08073_, _08072_);
  and (_08075_, _08074_, _34581_);
  and (_08076_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_08077_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_08078_, _08077_, _08076_);
  and (_08079_, _08078_, _34796_);
  or (_08080_, _08079_, _08075_);
  or (_08081_, _08080_, _34772_);
  and (_08082_, _08081_, _34803_);
  and (_08083_, _08082_, _08071_);
  or (_08084_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_08085_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_08086_, _08085_, _08084_);
  and (_08087_, _08086_, _34581_);
  or (_08088_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_08089_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_08090_, _08089_, _08088_);
  and (_08091_, _08090_, _34796_);
  or (_08092_, _08091_, _08087_);
  or (_08093_, _08092_, _34790_);
  or (_08094_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_08095_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_08096_, _08095_, _08094_);
  and (_08097_, _08096_, _34581_);
  or (_08098_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_08099_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_08100_, _08099_, _08098_);
  and (_08101_, _08100_, _34796_);
  or (_08102_, _08101_, _08097_);
  or (_08103_, _08102_, _34772_);
  and (_08104_, _08103_, _34719_);
  and (_08105_, _08104_, _08093_);
  or (_08106_, _08105_, _08083_);
  and (_08107_, _08106_, _34700_);
  or (_08108_, _08107_, _08061_);
  and (_08109_, _08108_, _34840_);
  or (_08110_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_08111_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_08112_, _08111_, _08110_);
  and (_08113_, _08112_, _34581_);
  or (_08114_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_08115_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_08116_, _08115_, _08114_);
  and (_08117_, _08116_, _34796_);
  or (_08118_, _08117_, _08113_);
  and (_08119_, _08118_, _34790_);
  or (_08120_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_08121_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_08122_, _08121_, _08120_);
  and (_08123_, _08122_, _34581_);
  or (_08124_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_08125_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_08126_, _08125_, _08124_);
  and (_08127_, _08126_, _34796_);
  or (_08128_, _08127_, _08123_);
  and (_08129_, _08128_, _34772_);
  or (_08130_, _08129_, _08119_);
  and (_08131_, _08130_, _34719_);
  and (_08132_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_08133_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_08134_, _08133_, _08132_);
  and (_08135_, _08134_, _34581_);
  and (_08136_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_08137_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_08138_, _08137_, _08136_);
  and (_08139_, _08138_, _34796_);
  or (_08140_, _08139_, _08135_);
  and (_08141_, _08140_, _34790_);
  and (_08142_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_08143_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_08144_, _08143_, _08142_);
  and (_08145_, _08144_, _34581_);
  and (_08146_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_08147_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_08148_, _08147_, _08146_);
  and (_08149_, _08148_, _34796_);
  or (_08150_, _08149_, _08145_);
  and (_08151_, _08150_, _34772_);
  or (_08152_, _08151_, _08141_);
  and (_08153_, _08152_, _34803_);
  or (_08154_, _08153_, _08131_);
  and (_08155_, _08154_, _34700_);
  or (_08156_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_08157_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  and (_08158_, _08157_, _34796_);
  and (_08159_, _08158_, _08156_);
  or (_08160_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_08161_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  and (_08162_, _08161_, _34581_);
  and (_08163_, _08162_, _08160_);
  or (_08164_, _08163_, _08159_);
  and (_08165_, _08164_, _34790_);
  or (_08166_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_08167_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_08168_, _08167_, _34796_);
  and (_08169_, _08168_, _08166_);
  or (_08170_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_08171_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  and (_08172_, _08171_, _34581_);
  and (_08173_, _08172_, _08170_);
  or (_08174_, _08173_, _08169_);
  and (_08175_, _08174_, _34772_);
  or (_08176_, _08175_, _08165_);
  and (_08177_, _08176_, _34719_);
  and (_08178_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  and (_08179_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_08180_, _08179_, _08178_);
  and (_08181_, _08180_, _34581_);
  and (_08182_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_08183_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _34796_);
  or (_08186_, _08185_, _08181_);
  and (_08187_, _08186_, _34790_);
  and (_08188_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  and (_08189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_08190_, _08189_, _08188_);
  and (_08191_, _08190_, _34581_);
  and (_08192_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_08193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_08194_, _08193_, _08192_);
  and (_08195_, _08194_, _34796_);
  or (_08196_, _08195_, _08191_);
  and (_08197_, _08196_, _34772_);
  or (_08198_, _08197_, _08187_);
  and (_08199_, _08198_, _34803_);
  or (_08200_, _08199_, _08177_);
  and (_08201_, _08200_, _34789_);
  or (_08202_, _08201_, _08155_);
  and (_08203_, _08202_, _34638_);
  or (_08204_, _08203_, _08109_);
  or (_08205_, _08204_, _34985_);
  and (_08206_, _08205_, _08015_);
  or (_08207_, _08206_, _34346_);
  and (_08208_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_08209_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_08210_, _08209_, _08208_);
  and (_08211_, _08210_, _34581_);
  and (_08212_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_08213_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_08214_, _08213_, _08212_);
  and (_08215_, _08214_, _34796_);
  or (_08216_, _08215_, _08211_);
  or (_08217_, _08216_, _34790_);
  and (_08218_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_08219_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_08220_, _08219_, _08218_);
  and (_08221_, _08220_, _34581_);
  and (_08222_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_08223_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_08224_, _08223_, _08222_);
  and (_08225_, _08224_, _34796_);
  or (_08226_, _08225_, _08221_);
  or (_08227_, _08226_, _34772_);
  and (_08228_, _08227_, _34803_);
  and (_08229_, _08228_, _08217_);
  or (_08230_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_08231_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_08232_, _08231_, _08230_);
  and (_08233_, _08232_, _34581_);
  or (_08234_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_08235_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_08236_, _08235_, _08234_);
  and (_08237_, _08236_, _34796_);
  or (_08238_, _08237_, _08233_);
  or (_08239_, _08238_, _34790_);
  or (_08240_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_08241_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_08242_, _08241_, _08240_);
  and (_08243_, _08242_, _34581_);
  or (_08244_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_08245_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_08246_, _08245_, _08244_);
  and (_08247_, _08246_, _34796_);
  or (_08248_, _08247_, _08243_);
  or (_08249_, _08248_, _34772_);
  and (_08250_, _08249_, _34719_);
  and (_08251_, _08250_, _08239_);
  or (_08252_, _08251_, _08229_);
  and (_08253_, _08252_, _34700_);
  and (_08254_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_08255_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_08256_, _08255_, _08254_);
  and (_08257_, _08256_, _34581_);
  and (_08258_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_08259_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_08260_, _08259_, _08258_);
  and (_08261_, _08260_, _34796_);
  or (_08262_, _08261_, _08257_);
  or (_08263_, _08262_, _34790_);
  and (_08264_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_08265_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_08266_, _08265_, _08264_);
  and (_08267_, _08266_, _34581_);
  and (_08268_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_08269_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_08270_, _08269_, _08268_);
  and (_08271_, _08270_, _34796_);
  or (_08272_, _08271_, _08267_);
  or (_08273_, _08272_, _34772_);
  and (_08274_, _08273_, _34803_);
  and (_08275_, _08274_, _08263_);
  or (_08276_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_08277_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_08278_, _08277_, _34796_);
  and (_08279_, _08278_, _08276_);
  or (_08280_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_08281_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_08282_, _08281_, _34581_);
  and (_08283_, _08282_, _08280_);
  or (_08284_, _08283_, _08279_);
  or (_08285_, _08284_, _34790_);
  or (_08286_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_08287_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_08288_, _08287_, _34796_);
  and (_08289_, _08288_, _08286_);
  or (_08290_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_08291_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_08292_, _08291_, _34581_);
  and (_08293_, _08292_, _08290_);
  or (_08294_, _08293_, _08289_);
  or (_08295_, _08294_, _34772_);
  and (_08296_, _08295_, _34719_);
  and (_08297_, _08296_, _08285_);
  or (_08298_, _08297_, _08275_);
  and (_08299_, _08298_, _34789_);
  or (_08300_, _08299_, _08253_);
  and (_08301_, _08300_, _34840_);
  and (_08302_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_08303_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_08304_, _08303_, _08302_);
  and (_08305_, _08304_, _34581_);
  and (_08306_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_08307_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_08308_, _08307_, _08306_);
  and (_08309_, _08308_, _34796_);
  or (_08310_, _08309_, _08305_);
  and (_08311_, _08310_, _34772_);
  and (_08312_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_08313_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_08314_, _08313_, _08312_);
  and (_08315_, _08314_, _34581_);
  and (_08316_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_08317_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_08318_, _08317_, _08316_);
  and (_08319_, _08318_, _34796_);
  or (_08320_, _08319_, _08315_);
  and (_08321_, _08320_, _34790_);
  or (_08322_, _08321_, _08311_);
  and (_08323_, _08322_, _34803_);
  or (_08324_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_08325_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_08326_, _08325_, _34796_);
  and (_08327_, _08326_, _08324_);
  or (_08328_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_08329_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_08330_, _08329_, _34581_);
  and (_08331_, _08330_, _08328_);
  or (_08332_, _08331_, _08327_);
  and (_08333_, _08332_, _34772_);
  or (_08334_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_08335_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_08336_, _08335_, _34796_);
  and (_08337_, _08336_, _08334_);
  or (_08338_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_08339_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_08340_, _08339_, _34581_);
  and (_08341_, _08340_, _08338_);
  or (_08342_, _08341_, _08337_);
  and (_08343_, _08342_, _34790_);
  or (_08344_, _08343_, _08333_);
  and (_08345_, _08344_, _34719_);
  or (_08346_, _08345_, _08323_);
  and (_08347_, _08346_, _34789_);
  and (_08348_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_08349_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_08350_, _08349_, _08348_);
  and (_08351_, _08350_, _34581_);
  and (_08352_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_08353_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_08354_, _08353_, _08352_);
  and (_08355_, _08354_, _34796_);
  or (_08356_, _08355_, _08351_);
  and (_08357_, _08356_, _34772_);
  and (_08358_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_08359_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_08360_, _08359_, _08358_);
  and (_08361_, _08360_, _34581_);
  and (_08362_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_08363_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_08364_, _08363_, _08362_);
  and (_08365_, _08364_, _34796_);
  or (_08366_, _08365_, _08361_);
  and (_08367_, _08366_, _34790_);
  or (_08368_, _08367_, _08357_);
  and (_08369_, _08368_, _34803_);
  or (_08370_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_08371_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_08372_, _08371_, _08370_);
  and (_08373_, _08372_, _34581_);
  or (_08374_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_08375_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_08376_, _08375_, _08374_);
  and (_08377_, _08376_, _34796_);
  or (_08378_, _08377_, _08373_);
  and (_08379_, _08378_, _34772_);
  or (_08380_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_08381_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_08382_, _08381_, _08380_);
  and (_08383_, _08382_, _34581_);
  or (_08384_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_08385_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_08386_, _08385_, _08384_);
  and (_08387_, _08386_, _34796_);
  or (_08388_, _08387_, _08383_);
  and (_08389_, _08388_, _34790_);
  or (_08390_, _08389_, _08379_);
  and (_08391_, _08390_, _34719_);
  or (_08392_, _08391_, _08369_);
  and (_08393_, _08392_, _34700_);
  or (_08394_, _08393_, _08347_);
  and (_08395_, _08394_, _34638_);
  or (_08396_, _08395_, _08301_);
  or (_08397_, _08396_, _34692_);
  and (_08398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_08399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_08400_, _08399_, _08398_);
  and (_08401_, _08400_, _34581_);
  and (_08402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_08403_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_08404_, _08403_, _08402_);
  and (_08405_, _08404_, _34796_);
  or (_08406_, _08405_, _08401_);
  or (_08407_, _08406_, _34790_);
  and (_08408_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_08409_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_08410_, _08409_, _08408_);
  and (_08411_, _08410_, _34581_);
  and (_08412_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_08413_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_08414_, _08413_, _08412_);
  and (_08415_, _08414_, _34796_);
  or (_08416_, _08415_, _08411_);
  or (_08417_, _08416_, _34772_);
  and (_08418_, _08417_, _34803_);
  and (_08419_, _08418_, _08407_);
  or (_08420_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_08421_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_08422_, _08421_, _34796_);
  and (_08423_, _08422_, _08420_);
  or (_08424_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_08425_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_08426_, _08425_, _34581_);
  and (_08427_, _08426_, _08424_);
  or (_08428_, _08427_, _08423_);
  or (_08429_, _08428_, _34790_);
  or (_08430_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_08431_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_08432_, _08431_, _34796_);
  and (_08433_, _08432_, _08430_);
  or (_08434_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_08435_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_08436_, _08435_, _34581_);
  and (_08437_, _08436_, _08434_);
  or (_08438_, _08437_, _08433_);
  or (_08439_, _08438_, _34772_);
  and (_08440_, _08439_, _34719_);
  and (_08441_, _08440_, _08429_);
  or (_08442_, _08441_, _08419_);
  and (_08443_, _08442_, _34789_);
  and (_08444_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_08445_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_08446_, _08445_, _08444_);
  and (_08447_, _08446_, _34581_);
  and (_08448_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_08449_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_08450_, _08449_, _08448_);
  and (_08451_, _08450_, _34796_);
  or (_08452_, _08451_, _08447_);
  or (_08453_, _08452_, _34790_);
  and (_08454_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_08455_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_08456_, _08455_, _08454_);
  and (_08457_, _08456_, _34581_);
  and (_08458_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_08459_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_08460_, _08459_, _08458_);
  and (_08461_, _08460_, _34796_);
  or (_08462_, _08461_, _08457_);
  or (_08463_, _08462_, _34772_);
  and (_08464_, _08463_, _34803_);
  and (_08465_, _08464_, _08453_);
  or (_08466_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_08467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_08468_, _08467_, _08466_);
  and (_08469_, _08468_, _34581_);
  or (_08470_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_08471_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_08472_, _08471_, _08470_);
  and (_08473_, _08472_, _34796_);
  or (_08474_, _08473_, _08469_);
  or (_08475_, _08474_, _34790_);
  or (_08476_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_08477_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_08478_, _08477_, _08476_);
  and (_08479_, _08478_, _34581_);
  or (_08480_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_08481_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_08482_, _08481_, _08480_);
  and (_08483_, _08482_, _34796_);
  or (_08484_, _08483_, _08479_);
  or (_08485_, _08484_, _34772_);
  and (_08486_, _08485_, _34719_);
  and (_08487_, _08486_, _08475_);
  or (_08488_, _08487_, _08465_);
  and (_08489_, _08488_, _34700_);
  or (_08490_, _08489_, _08443_);
  and (_08491_, _08490_, _34840_);
  or (_08492_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_08493_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_08494_, _08493_, _08492_);
  and (_08495_, _08494_, _34581_);
  or (_08496_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_08497_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_08498_, _08497_, _08496_);
  and (_08499_, _08498_, _34796_);
  or (_08500_, _08499_, _08495_);
  and (_08501_, _08500_, _34790_);
  or (_08502_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_08503_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_08504_, _08503_, _08502_);
  and (_08505_, _08504_, _34581_);
  or (_08506_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_08507_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_08508_, _08507_, _08506_);
  and (_08509_, _08508_, _34796_);
  or (_08510_, _08509_, _08505_);
  and (_08511_, _08510_, _34772_);
  or (_08512_, _08511_, _08501_);
  and (_08513_, _08512_, _34719_);
  and (_08514_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_08515_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_08516_, _08515_, _08514_);
  and (_08517_, _08516_, _34581_);
  and (_08518_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_08519_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_08520_, _08519_, _08518_);
  and (_08521_, _08520_, _34796_);
  or (_08522_, _08521_, _08517_);
  and (_08523_, _08522_, _34790_);
  and (_08524_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_08525_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_08526_, _08525_, _08524_);
  and (_08527_, _08526_, _34581_);
  and (_08528_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_08529_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_08530_, _08529_, _08528_);
  and (_08531_, _08530_, _34796_);
  or (_08532_, _08531_, _08527_);
  and (_08533_, _08532_, _34772_);
  or (_08534_, _08533_, _08523_);
  and (_08535_, _08534_, _34803_);
  or (_08536_, _08535_, _08513_);
  and (_08537_, _08536_, _34700_);
  or (_08538_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_08539_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_08540_, _08539_, _34796_);
  and (_08541_, _08540_, _08538_);
  or (_08542_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_08543_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_08544_, _08543_, _34581_);
  and (_08545_, _08544_, _08542_);
  or (_08546_, _08545_, _08541_);
  and (_08547_, _08546_, _34790_);
  or (_08548_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_08549_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_08550_, _08549_, _34796_);
  and (_08551_, _08550_, _08548_);
  or (_08552_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_08553_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_08554_, _08553_, _34581_);
  and (_08555_, _08554_, _08552_);
  or (_08556_, _08555_, _08551_);
  and (_08557_, _08556_, _34772_);
  or (_08558_, _08557_, _08547_);
  and (_08559_, _08558_, _34719_);
  and (_08560_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_08561_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_08562_, _08561_, _08560_);
  and (_08563_, _08562_, _34581_);
  and (_08564_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_08565_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_08566_, _08565_, _08564_);
  and (_08567_, _08566_, _34796_);
  or (_08568_, _08567_, _08563_);
  and (_08569_, _08568_, _34790_);
  and (_08570_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_08571_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_08572_, _08571_, _08570_);
  and (_08573_, _08572_, _34581_);
  and (_08574_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_08575_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_08576_, _08575_, _08574_);
  and (_08577_, _08576_, _34796_);
  or (_08578_, _08577_, _08573_);
  and (_08579_, _08578_, _34772_);
  or (_08580_, _08579_, _08569_);
  and (_08581_, _08580_, _34803_);
  or (_08582_, _08581_, _08559_);
  and (_08583_, _08582_, _34789_);
  or (_08584_, _08583_, _08537_);
  and (_08585_, _08584_, _34638_);
  or (_08586_, _08585_, _08491_);
  or (_08587_, _08586_, _34985_);
  and (_08588_, _08587_, _08397_);
  or (_08589_, _08588_, _35178_);
  and (_08590_, _08589_, _08207_);
  or (_08591_, _08590_, _34788_);
  or (_08592_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_08593_, _08592_, _38997_);
  and (_38984_[3], _08593_, _08591_);
  and (_08594_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_08595_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_08596_, _08595_, _08594_);
  and (_08597_, _08596_, _34581_);
  and (_08598_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_08599_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_08600_, _08599_, _08598_);
  and (_08601_, _08600_, _34796_);
  or (_08602_, _08601_, _08597_);
  or (_08603_, _08602_, _34790_);
  and (_08604_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_08605_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_08606_, _08605_, _08604_);
  and (_08607_, _08606_, _34581_);
  and (_08608_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_08609_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_08610_, _08609_, _08608_);
  and (_08611_, _08610_, _34796_);
  or (_08612_, _08611_, _08607_);
  or (_08613_, _08612_, _34772_);
  and (_08614_, _08613_, _34803_);
  and (_08615_, _08614_, _08603_);
  or (_08616_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_08617_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_08618_, _08617_, _08616_);
  and (_08619_, _08618_, _34581_);
  or (_08620_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_08621_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_08622_, _08621_, _08620_);
  and (_08623_, _08622_, _34796_);
  or (_08624_, _08623_, _08619_);
  or (_08625_, _08624_, _34790_);
  or (_08626_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_08627_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_08628_, _08627_, _08626_);
  and (_08629_, _08628_, _34581_);
  or (_08630_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_08631_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_08632_, _08631_, _08630_);
  and (_08633_, _08632_, _34796_);
  or (_08634_, _08633_, _08629_);
  or (_08635_, _08634_, _34772_);
  and (_08636_, _08635_, _34719_);
  and (_08637_, _08636_, _08625_);
  or (_08638_, _08637_, _08615_);
  or (_08639_, _08638_, _34789_);
  and (_08640_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_08641_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_08642_, _08641_, _08640_);
  and (_08643_, _08642_, _34581_);
  and (_08644_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_08645_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_08646_, _08645_, _08644_);
  and (_08647_, _08646_, _34796_);
  or (_08648_, _08647_, _08643_);
  or (_08649_, _08648_, _34790_);
  and (_08650_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_08651_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_08652_, _08651_, _08650_);
  and (_08653_, _08652_, _34581_);
  and (_08654_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_08655_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_08656_, _08655_, _08654_);
  and (_08657_, _08656_, _34796_);
  or (_08658_, _08657_, _08653_);
  or (_08659_, _08658_, _34772_);
  and (_08660_, _08659_, _34803_);
  and (_08661_, _08660_, _08649_);
  or (_08662_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_08663_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_08664_, _08663_, _34796_);
  and (_08665_, _08664_, _08662_);
  or (_08666_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_08667_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_08668_, _08667_, _34581_);
  and (_08669_, _08668_, _08666_);
  or (_08670_, _08669_, _08665_);
  or (_08671_, _08670_, _34790_);
  or (_08672_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_08673_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_08674_, _08673_, _34796_);
  and (_08675_, _08674_, _08672_);
  or (_08676_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_08677_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_08678_, _08677_, _34581_);
  and (_08679_, _08678_, _08676_);
  or (_08680_, _08679_, _08675_);
  or (_08681_, _08680_, _34772_);
  and (_08682_, _08681_, _34719_);
  and (_08683_, _08682_, _08671_);
  or (_08684_, _08683_, _08661_);
  or (_08685_, _08684_, _34700_);
  and (_08686_, _08685_, _34840_);
  and (_08687_, _08686_, _08639_);
  and (_08688_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_08689_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_08690_, _08689_, _08688_);
  and (_08691_, _08690_, _34581_);
  and (_08692_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_08693_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_08694_, _08693_, _08692_);
  and (_08695_, _08694_, _34796_);
  or (_08696_, _08695_, _08691_);
  and (_08697_, _08696_, _34772_);
  and (_08698_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_08699_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_08700_, _08699_, _08698_);
  and (_08701_, _08700_, _34581_);
  and (_08702_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_08703_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_08704_, _08703_, _08702_);
  and (_08705_, _08704_, _34796_);
  or (_08706_, _08705_, _08701_);
  and (_08707_, _08706_, _34790_);
  or (_08708_, _08707_, _34719_);
  or (_08709_, _08708_, _08697_);
  or (_08710_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_08711_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_08712_, _08711_, _34796_);
  and (_08713_, _08712_, _08710_);
  or (_08714_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_08715_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_08716_, _08715_, _34581_);
  and (_08717_, _08716_, _08714_);
  or (_08718_, _08717_, _08713_);
  and (_08719_, _08718_, _34772_);
  or (_08720_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_08721_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_08722_, _08721_, _34796_);
  and (_08723_, _08722_, _08720_);
  or (_08724_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_08725_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_08726_, _08725_, _34581_);
  and (_08727_, _08726_, _08724_);
  or (_08728_, _08727_, _08723_);
  and (_08729_, _08728_, _34790_);
  or (_08730_, _08729_, _34803_);
  or (_08731_, _08730_, _08719_);
  and (_08732_, _08731_, _08709_);
  or (_08733_, _08732_, _34700_);
  and (_08734_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_08735_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_08736_, _08735_, _08734_);
  and (_08737_, _08736_, _34581_);
  and (_08738_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_08739_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_08740_, _08739_, _08738_);
  and (_08741_, _08740_, _34796_);
  or (_08742_, _08741_, _08737_);
  and (_08743_, _08742_, _34772_);
  and (_08744_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_08745_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_08746_, _08745_, _08744_);
  and (_08747_, _08746_, _34581_);
  and (_08748_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_08749_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_08750_, _08749_, _08748_);
  and (_08751_, _08750_, _34796_);
  or (_08752_, _08751_, _08747_);
  and (_08753_, _08752_, _34790_);
  or (_08754_, _08753_, _34719_);
  or (_08755_, _08754_, _08743_);
  or (_08756_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_08757_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_08758_, _08757_, _08756_);
  and (_08759_, _08758_, _34581_);
  or (_08760_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_08761_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_08762_, _08761_, _08760_);
  and (_08763_, _08762_, _34796_);
  or (_08764_, _08763_, _08759_);
  and (_08765_, _08764_, _34772_);
  or (_08766_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_08767_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_08768_, _08767_, _08766_);
  and (_08769_, _08768_, _34581_);
  or (_08770_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_08771_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_08772_, _08771_, _08770_);
  and (_08773_, _08772_, _34796_);
  or (_08774_, _08773_, _08769_);
  and (_08775_, _08774_, _34790_);
  or (_08776_, _08775_, _34803_);
  or (_08777_, _08776_, _08765_);
  and (_08778_, _08777_, _08755_);
  or (_08779_, _08778_, _34789_);
  and (_08780_, _08779_, _34638_);
  and (_08781_, _08780_, _08733_);
  or (_08782_, _08781_, _08687_);
  or (_08783_, _08782_, _34692_);
  and (_08784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and (_08785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_08786_, _08785_, _08784_);
  and (_08787_, _08786_, _34581_);
  and (_08788_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and (_08789_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_08790_, _08789_, _08788_);
  and (_08791_, _08790_, _34796_);
  or (_08792_, _08791_, _08787_);
  and (_08793_, _08792_, _34772_);
  and (_08794_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and (_08795_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_08796_, _08795_, _08794_);
  and (_08797_, _08796_, _34581_);
  and (_08798_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and (_08799_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_08800_, _08799_, _08798_);
  and (_08801_, _08800_, _34796_);
  or (_08802_, _08801_, _08797_);
  and (_08803_, _08802_, _34790_);
  or (_08804_, _08803_, _34719_);
  or (_08805_, _08804_, _08793_);
  or (_08806_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_08807_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and (_08808_, _08807_, _08806_);
  and (_08809_, _08808_, _34581_);
  or (_08810_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_08811_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  and (_08812_, _08811_, _08810_);
  and (_08813_, _08812_, _34796_);
  or (_08814_, _08813_, _08809_);
  and (_08815_, _08814_, _34772_);
  or (_08816_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_08817_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and (_08818_, _08817_, _08816_);
  and (_08819_, _08818_, _34581_);
  or (_08820_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_08821_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  and (_08822_, _08821_, _08820_);
  and (_08823_, _08822_, _34796_);
  or (_08824_, _08823_, _08819_);
  and (_08825_, _08824_, _34790_);
  or (_08826_, _08825_, _34803_);
  or (_08827_, _08826_, _08815_);
  and (_08828_, _08827_, _08805_);
  or (_08829_, _08828_, _34700_);
  and (_08830_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_08831_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_08832_, _08831_, _08830_);
  and (_08833_, _08832_, _34581_);
  and (_08834_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_08835_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_08836_, _08835_, _08834_);
  and (_08837_, _08836_, _34796_);
  or (_08838_, _08837_, _08833_);
  and (_08839_, _08838_, _34772_);
  and (_08840_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_08841_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_08842_, _08841_, _08840_);
  and (_08843_, _08842_, _34581_);
  and (_08844_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_08845_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_08846_, _08845_, _08844_);
  and (_08847_, _08846_, _34796_);
  or (_08848_, _08847_, _08843_);
  and (_08849_, _08848_, _34790_);
  or (_08850_, _08849_, _34719_);
  or (_08851_, _08850_, _08839_);
  or (_08852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_08853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_08854_, _08853_, _08852_);
  and (_08855_, _08854_, _34581_);
  or (_08856_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_08857_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_08858_, _08857_, _08856_);
  and (_08859_, _08858_, _34796_);
  or (_08860_, _08859_, _08855_);
  and (_08861_, _08860_, _34772_);
  or (_08862_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_08863_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_08864_, _08863_, _08862_);
  and (_08865_, _08864_, _34581_);
  or (_08866_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_08867_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_08868_, _08867_, _08866_);
  and (_08869_, _08868_, _34796_);
  or (_08870_, _08869_, _08865_);
  and (_08871_, _08870_, _34790_);
  or (_08872_, _08871_, _34803_);
  or (_08873_, _08872_, _08861_);
  and (_08874_, _08873_, _08851_);
  or (_08875_, _08874_, _34789_);
  and (_08876_, _08875_, _34638_);
  and (_08877_, _08876_, _08829_);
  and (_08878_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_08879_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_08880_, _08879_, _08878_);
  and (_08881_, _08880_, _34796_);
  and (_08882_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_08883_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_08884_, _08883_, _08882_);
  and (_08885_, _08884_, _34581_);
  or (_08886_, _08885_, _08881_);
  or (_08887_, _08886_, _34790_);
  and (_08888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_08889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_08890_, _08889_, _08888_);
  and (_08891_, _08890_, _34796_);
  and (_08892_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_08893_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_08894_, _08893_, _08892_);
  and (_08895_, _08894_, _34581_);
  or (_08896_, _08895_, _08891_);
  or (_08897_, _08896_, _34772_);
  and (_08898_, _08897_, _34803_);
  and (_08899_, _08898_, _08887_);
  or (_08900_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_08901_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_08902_, _08901_, _34581_);
  and (_08903_, _08902_, _08900_);
  or (_08904_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_08905_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_08906_, _08905_, _34796_);
  and (_08907_, _08906_, _08904_);
  or (_08908_, _08907_, _08903_);
  or (_08909_, _08908_, _34790_);
  or (_08910_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_08911_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_08912_, _08911_, _34581_);
  and (_08913_, _08912_, _08910_);
  or (_08914_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_08915_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_08916_, _08915_, _34796_);
  and (_08917_, _08916_, _08914_);
  or (_08918_, _08917_, _08913_);
  or (_08919_, _08918_, _34772_);
  and (_08920_, _08919_, _34719_);
  and (_08921_, _08920_, _08909_);
  or (_08922_, _08921_, _08899_);
  and (_08923_, _08922_, _34789_);
  and (_08924_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_08925_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_08926_, _08925_, _34581_);
  or (_08927_, _08926_, _08924_);
  and (_08928_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_08929_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_08930_, _08929_, _34796_);
  or (_08931_, _08930_, _08928_);
  and (_08932_, _08931_, _08927_);
  or (_08933_, _08932_, _34790_);
  and (_08934_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_08935_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_08936_, _08935_, _34581_);
  or (_08937_, _08936_, _08934_);
  and (_08938_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_08939_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_08940_, _08939_, _34796_);
  or (_08941_, _08940_, _08938_);
  and (_08942_, _08941_, _08937_);
  or (_08943_, _08942_, _34772_);
  and (_08944_, _08943_, _34803_);
  and (_08945_, _08944_, _08933_);
  or (_08946_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_08947_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_08948_, _08947_, _08946_);
  or (_08949_, _08948_, _34796_);
  or (_08950_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_08951_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_08952_, _08951_, _08950_);
  or (_08953_, _08952_, _34581_);
  and (_08954_, _08953_, _08949_);
  or (_08955_, _08954_, _34790_);
  or (_08956_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_08957_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_08958_, _08957_, _08956_);
  or (_08959_, _08958_, _34796_);
  or (_08960_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_08961_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_08962_, _08961_, _08960_);
  or (_08963_, _08962_, _34581_);
  and (_08964_, _08963_, _08959_);
  or (_08965_, _08964_, _34772_);
  and (_08966_, _08965_, _34719_);
  and (_08967_, _08966_, _08955_);
  or (_08968_, _08967_, _08945_);
  and (_08969_, _08968_, _34700_);
  or (_08970_, _08969_, _08923_);
  and (_08971_, _08970_, _34840_);
  or (_08972_, _08971_, _08877_);
  or (_08973_, _08972_, _34985_);
  and (_08974_, _08973_, _08783_);
  or (_08975_, _08974_, _34346_);
  and (_08976_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_08977_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_08978_, _08977_, _08976_);
  and (_08979_, _08978_, _34581_);
  and (_08980_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_08981_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_08982_, _08981_, _08980_);
  and (_08983_, _08982_, _34796_);
  or (_08984_, _08983_, _08979_);
  or (_08985_, _08984_, _34790_);
  and (_08986_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_08987_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_08988_, _08987_, _08986_);
  and (_08989_, _08988_, _34581_);
  and (_08990_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_08991_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_08992_, _08991_, _08990_);
  and (_08993_, _08992_, _34796_);
  or (_08994_, _08993_, _08989_);
  or (_08995_, _08994_, _34772_);
  and (_08996_, _08995_, _34803_);
  and (_08997_, _08996_, _08985_);
  or (_08998_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_08999_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_09000_, _08999_, _08998_);
  and (_09001_, _09000_, _34581_);
  or (_09002_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_09003_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_09004_, _09003_, _09002_);
  and (_09005_, _09004_, _34796_);
  or (_09006_, _09005_, _09001_);
  or (_09007_, _09006_, _34790_);
  or (_09008_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_09009_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_09010_, _09009_, _09008_);
  and (_09011_, _09010_, _34581_);
  or (_09012_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_09013_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_09014_, _09013_, _09012_);
  and (_09015_, _09014_, _34796_);
  or (_09016_, _09015_, _09011_);
  or (_09017_, _09016_, _34772_);
  and (_09018_, _09017_, _34719_);
  and (_09019_, _09018_, _09007_);
  or (_09020_, _09019_, _08997_);
  and (_09021_, _09020_, _34700_);
  and (_09022_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_09023_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_09024_, _09023_, _09022_);
  and (_09025_, _09024_, _34581_);
  and (_09026_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_09027_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_09028_, _09027_, _09026_);
  and (_09029_, _09028_, _34796_);
  or (_09030_, _09029_, _09025_);
  or (_09031_, _09030_, _34790_);
  and (_09032_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_09033_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_09034_, _09033_, _09032_);
  and (_09035_, _09034_, _34581_);
  and (_09036_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_09037_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_09038_, _09037_, _09036_);
  and (_09039_, _09038_, _34796_);
  or (_09040_, _09039_, _09035_);
  or (_09041_, _09040_, _34772_);
  and (_09042_, _09041_, _34803_);
  and (_09043_, _09042_, _09031_);
  or (_09044_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_09045_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_09046_, _09045_, _34796_);
  and (_09047_, _09046_, _09044_);
  or (_09048_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_09049_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_09050_, _09049_, _34581_);
  and (_09051_, _09050_, _09048_);
  or (_09052_, _09051_, _09047_);
  or (_09053_, _09052_, _34790_);
  or (_09054_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_09055_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_09056_, _09055_, _34796_);
  and (_09057_, _09056_, _09054_);
  or (_09058_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_09059_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_09060_, _09059_, _34581_);
  and (_09061_, _09060_, _09058_);
  or (_09062_, _09061_, _09057_);
  or (_09063_, _09062_, _34772_);
  and (_09064_, _09063_, _34719_);
  and (_09065_, _09064_, _09053_);
  or (_09066_, _09065_, _09043_);
  and (_09067_, _09066_, _34789_);
  or (_09068_, _09067_, _09021_);
  and (_09069_, _09068_, _34840_);
  and (_09070_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_09071_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_09072_, _09071_, _09070_);
  and (_09073_, _09072_, _34581_);
  and (_09074_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_09075_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_09076_, _09075_, _09074_);
  and (_09077_, _09076_, _34796_);
  or (_09078_, _09077_, _09073_);
  and (_09079_, _09078_, _34772_);
  and (_09080_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_09081_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_09082_, _09081_, _09080_);
  and (_09083_, _09082_, _34581_);
  and (_09084_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_09085_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_09086_, _09085_, _09084_);
  and (_09087_, _09086_, _34796_);
  or (_09088_, _09087_, _09083_);
  and (_09089_, _09088_, _34790_);
  or (_09090_, _09089_, _09079_);
  and (_09091_, _09090_, _34803_);
  or (_09092_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_09093_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_09094_, _09093_, _34796_);
  and (_09095_, _09094_, _09092_);
  or (_09096_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_09097_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_09098_, _09097_, _34581_);
  and (_09099_, _09098_, _09096_);
  or (_09100_, _09099_, _09095_);
  and (_09101_, _09100_, _34772_);
  or (_09102_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_09103_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_09104_, _09103_, _34796_);
  and (_09105_, _09104_, _09102_);
  or (_09106_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_09107_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_09108_, _09107_, _34581_);
  and (_09109_, _09108_, _09106_);
  or (_09110_, _09109_, _09105_);
  and (_09111_, _09110_, _34790_);
  or (_09112_, _09111_, _09101_);
  and (_09113_, _09112_, _34719_);
  or (_09114_, _09113_, _09091_);
  and (_09115_, _09114_, _34789_);
  and (_09116_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_09117_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_09118_, _09117_, _09116_);
  and (_09119_, _09118_, _34581_);
  and (_09120_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_09121_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_09122_, _09121_, _09120_);
  and (_09123_, _09122_, _34796_);
  or (_09124_, _09123_, _09119_);
  and (_09125_, _09124_, _34772_);
  and (_09126_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_09127_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_09128_, _09127_, _09126_);
  and (_09129_, _09128_, _34581_);
  and (_09130_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_09131_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_09132_, _09131_, _09130_);
  and (_09133_, _09132_, _34796_);
  or (_09134_, _09133_, _09129_);
  and (_09135_, _09134_, _34790_);
  or (_09136_, _09135_, _09125_);
  and (_09137_, _09136_, _34803_);
  or (_09138_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_09139_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_09140_, _09139_, _09138_);
  and (_09141_, _09140_, _34581_);
  or (_09142_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_09143_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_09144_, _09143_, _09142_);
  and (_09145_, _09144_, _34796_);
  or (_09146_, _09145_, _09141_);
  and (_09147_, _09146_, _34772_);
  or (_09148_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_09149_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_09150_, _09149_, _09148_);
  and (_09151_, _09150_, _34581_);
  or (_09152_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_09153_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_09154_, _09153_, _09152_);
  and (_09155_, _09154_, _34796_);
  or (_09156_, _09155_, _09151_);
  and (_09157_, _09156_, _34790_);
  or (_09158_, _09157_, _09147_);
  and (_09159_, _09158_, _34719_);
  or (_09160_, _09159_, _09137_);
  and (_09161_, _09160_, _34700_);
  or (_09162_, _09161_, _09115_);
  and (_09163_, _09162_, _34638_);
  or (_09164_, _09163_, _09069_);
  or (_09165_, _09164_, _34692_);
  and (_09166_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_09167_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_09168_, _09167_, _09166_);
  and (_09169_, _09168_, _34581_);
  and (_09170_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_09171_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_09172_, _09171_, _09170_);
  and (_09173_, _09172_, _34796_);
  or (_09174_, _09173_, _09169_);
  or (_09175_, _09174_, _34790_);
  and (_09176_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_09177_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_09178_, _09177_, _09176_);
  and (_09179_, _09178_, _34581_);
  and (_09180_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_09181_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_09182_, _09181_, _09180_);
  and (_09183_, _09182_, _34796_);
  or (_09184_, _09183_, _09179_);
  or (_09185_, _09184_, _34772_);
  and (_09186_, _09185_, _34803_);
  and (_09187_, _09186_, _09175_);
  or (_09188_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_09189_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_09190_, _09189_, _34796_);
  and (_09191_, _09190_, _09188_);
  or (_09192_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_09193_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_09194_, _09193_, _34581_);
  and (_09195_, _09194_, _09192_);
  or (_09196_, _09195_, _09191_);
  or (_09197_, _09196_, _34790_);
  or (_09198_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_09199_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_09200_, _09199_, _34796_);
  and (_09201_, _09200_, _09198_);
  or (_09202_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_09203_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_09204_, _09203_, _34581_);
  and (_09205_, _09204_, _09202_);
  or (_09206_, _09205_, _09201_);
  or (_09207_, _09206_, _34772_);
  and (_09208_, _09207_, _34719_);
  and (_09209_, _09208_, _09197_);
  or (_09210_, _09209_, _09187_);
  and (_09211_, _09210_, _34789_);
  and (_09212_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_09213_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_09214_, _09213_, _09212_);
  and (_09215_, _09214_, _34581_);
  and (_09216_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_09217_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_09218_, _09217_, _09216_);
  and (_09219_, _09218_, _34796_);
  or (_09220_, _09219_, _09215_);
  or (_09221_, _09220_, _34790_);
  and (_09222_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_09223_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_09224_, _09223_, _09222_);
  and (_09225_, _09224_, _34581_);
  and (_09226_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_09227_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_09228_, _09227_, _09226_);
  and (_09229_, _09228_, _34796_);
  or (_09230_, _09229_, _09225_);
  or (_09231_, _09230_, _34772_);
  and (_09232_, _09231_, _34803_);
  and (_09233_, _09232_, _09221_);
  or (_09234_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_09235_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_09236_, _09235_, _09234_);
  and (_09237_, _09236_, _34581_);
  or (_09238_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_09239_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_09240_, _09239_, _09238_);
  and (_09241_, _09240_, _34796_);
  or (_09242_, _09241_, _09237_);
  or (_09243_, _09242_, _34790_);
  or (_09244_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_09245_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_09246_, _09245_, _09244_);
  and (_09247_, _09246_, _34581_);
  or (_09248_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_09249_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_09250_, _09249_, _09248_);
  and (_09251_, _09250_, _34796_);
  or (_09252_, _09251_, _09247_);
  or (_09253_, _09252_, _34772_);
  and (_09254_, _09253_, _34719_);
  and (_09255_, _09254_, _09243_);
  or (_09256_, _09255_, _09233_);
  and (_09257_, _09256_, _34700_);
  or (_09258_, _09257_, _09211_);
  and (_09259_, _09258_, _34840_);
  or (_09260_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_09261_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_09262_, _09261_, _09260_);
  and (_09263_, _09262_, _34581_);
  or (_09264_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_09265_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_09266_, _09265_, _09264_);
  and (_09267_, _09266_, _34796_);
  or (_09268_, _09267_, _09263_);
  and (_09269_, _09268_, _34790_);
  or (_09270_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_09271_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_09272_, _09271_, _09270_);
  and (_09273_, _09272_, _34581_);
  or (_09274_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_09275_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_09276_, _09275_, _09274_);
  and (_09277_, _09276_, _34796_);
  or (_09278_, _09277_, _09273_);
  and (_09279_, _09278_, _34772_);
  or (_09280_, _09279_, _09269_);
  and (_09281_, _09280_, _34719_);
  and (_09282_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_09283_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_09284_, _09283_, _09282_);
  and (_09285_, _09284_, _34581_);
  and (_09286_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_09287_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_09288_, _09287_, _09286_);
  and (_09289_, _09288_, _34796_);
  or (_09290_, _09289_, _09285_);
  and (_09291_, _09290_, _34790_);
  and (_09292_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_09293_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_09294_, _09293_, _09292_);
  and (_09295_, _09294_, _34581_);
  and (_09296_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_09297_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_09298_, _09297_, _09296_);
  and (_09299_, _09298_, _34796_);
  or (_09300_, _09299_, _09295_);
  and (_09301_, _09300_, _34772_);
  or (_09302_, _09301_, _09291_);
  and (_09303_, _09302_, _34803_);
  or (_09304_, _09303_, _09281_);
  and (_09305_, _09304_, _34700_);
  or (_09306_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_09307_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_09308_, _09307_, _34796_);
  and (_09309_, _09308_, _09306_);
  or (_09310_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_09311_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_09312_, _09311_, _34581_);
  and (_09313_, _09312_, _09310_);
  or (_09314_, _09313_, _09309_);
  and (_09315_, _09314_, _34790_);
  or (_09316_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_09317_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_09318_, _09317_, _34796_);
  and (_09319_, _09318_, _09316_);
  or (_09320_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_09321_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_09322_, _09321_, _34581_);
  and (_09323_, _09322_, _09320_);
  or (_09324_, _09323_, _09319_);
  and (_09325_, _09324_, _34772_);
  or (_09326_, _09325_, _09315_);
  and (_09327_, _09326_, _34719_);
  and (_09328_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_09329_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_09330_, _09329_, _09328_);
  and (_09331_, _09330_, _34581_);
  and (_09332_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_09333_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_09334_, _09333_, _09332_);
  and (_09335_, _09334_, _34796_);
  or (_09336_, _09335_, _09331_);
  and (_09337_, _09336_, _34790_);
  and (_09338_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_09339_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_09340_, _09339_, _09338_);
  and (_09341_, _09340_, _34581_);
  and (_09342_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_09343_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_09344_, _09343_, _09342_);
  and (_09345_, _09344_, _34796_);
  or (_09346_, _09345_, _09341_);
  and (_09347_, _09346_, _34772_);
  or (_09348_, _09347_, _09337_);
  and (_09349_, _09348_, _34803_);
  or (_09350_, _09349_, _09327_);
  and (_09351_, _09350_, _34789_);
  or (_09352_, _09351_, _09305_);
  and (_09353_, _09352_, _34638_);
  or (_09354_, _09353_, _09259_);
  or (_09355_, _09354_, _34985_);
  and (_09356_, _09355_, _09165_);
  or (_09357_, _09356_, _35178_);
  and (_09358_, _09357_, _08975_);
  or (_09359_, _09358_, _34788_);
  or (_09360_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_09361_, _09360_, _38997_);
  and (_38984_[4], _09361_, _09359_);
  and (_09362_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_09363_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_09364_, _09363_, _09362_);
  and (_09365_, _09364_, _34581_);
  and (_09366_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_09367_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_09368_, _09367_, _09366_);
  and (_09369_, _09368_, _34796_);
  or (_09370_, _09369_, _09365_);
  or (_09371_, _09370_, _34790_);
  and (_09372_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_09373_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_09374_, _09373_, _09372_);
  and (_09375_, _09374_, _34581_);
  and (_09376_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_09377_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_09378_, _09377_, _09376_);
  and (_09379_, _09378_, _34796_);
  or (_09380_, _09379_, _09375_);
  or (_09381_, _09380_, _34772_);
  and (_09382_, _09381_, _34803_);
  and (_09383_, _09382_, _09371_);
  or (_09384_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_09385_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_09386_, _09385_, _09384_);
  and (_09387_, _09386_, _34581_);
  or (_09388_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_09389_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_09390_, _09389_, _09388_);
  and (_09391_, _09390_, _34796_);
  or (_09392_, _09391_, _09387_);
  or (_09393_, _09392_, _34790_);
  or (_09394_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_09395_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_09396_, _09395_, _09394_);
  and (_09397_, _09396_, _34581_);
  or (_09398_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_09399_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_09400_, _09399_, _09398_);
  and (_09401_, _09400_, _34796_);
  or (_09402_, _09401_, _09397_);
  or (_09403_, _09402_, _34772_);
  and (_09404_, _09403_, _34719_);
  and (_09405_, _09404_, _09393_);
  or (_09406_, _09405_, _09383_);
  and (_09407_, _09406_, _34700_);
  and (_09408_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_09409_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_09410_, _09409_, _09408_);
  and (_09411_, _09410_, _34581_);
  and (_09412_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_09413_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_09414_, _09413_, _09412_);
  and (_09415_, _09414_, _34796_);
  or (_09416_, _09415_, _09411_);
  or (_09417_, _09416_, _34790_);
  and (_09418_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_09419_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_09420_, _09419_, _09418_);
  and (_09421_, _09420_, _34581_);
  and (_09422_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_09423_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_09424_, _09423_, _09422_);
  and (_09425_, _09424_, _34796_);
  or (_09426_, _09425_, _09421_);
  or (_09427_, _09426_, _34772_);
  and (_09428_, _09427_, _34803_);
  and (_09429_, _09428_, _09417_);
  or (_09430_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_09431_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_09432_, _09431_, _34796_);
  and (_09433_, _09432_, _09430_);
  or (_09434_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_09435_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_09436_, _09435_, _34581_);
  and (_09437_, _09436_, _09434_);
  or (_09438_, _09437_, _09433_);
  or (_09439_, _09438_, _34790_);
  or (_09440_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_09441_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_09442_, _09441_, _34796_);
  and (_09443_, _09442_, _09440_);
  or (_09444_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_09445_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_09446_, _09445_, _34581_);
  and (_09447_, _09446_, _09444_);
  or (_09448_, _09447_, _09443_);
  or (_09449_, _09448_, _34772_);
  and (_09450_, _09449_, _34719_);
  and (_09451_, _09450_, _09439_);
  or (_09452_, _09451_, _09429_);
  and (_09453_, _09452_, _34789_);
  or (_09454_, _09453_, _09407_);
  and (_09455_, _09454_, _34840_);
  and (_09456_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_09457_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_09458_, _09457_, _09456_);
  and (_09459_, _09458_, _34581_);
  and (_09460_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_09461_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_09462_, _09461_, _09460_);
  and (_09463_, _09462_, _34796_);
  or (_09464_, _09463_, _09459_);
  and (_09465_, _09464_, _34772_);
  and (_09466_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_09467_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_09468_, _09467_, _09466_);
  and (_09469_, _09468_, _34581_);
  and (_09470_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_09471_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_09472_, _09471_, _09470_);
  and (_09473_, _09472_, _34796_);
  or (_09474_, _09473_, _09469_);
  and (_09475_, _09474_, _34790_);
  or (_09476_, _09475_, _09465_);
  and (_09477_, _09476_, _34803_);
  or (_09478_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_09479_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_09480_, _09479_, _34796_);
  and (_09481_, _09480_, _09478_);
  or (_09482_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_09483_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_09484_, _09483_, _34581_);
  and (_09485_, _09484_, _09482_);
  or (_09486_, _09485_, _09481_);
  and (_09487_, _09486_, _34772_);
  or (_09488_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_09489_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_09490_, _09489_, _34796_);
  and (_09491_, _09490_, _09488_);
  or (_09492_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_09493_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_09494_, _09493_, _34581_);
  and (_09495_, _09494_, _09492_);
  or (_09496_, _09495_, _09491_);
  and (_09497_, _09496_, _34790_);
  or (_09498_, _09497_, _09487_);
  and (_09499_, _09498_, _34719_);
  or (_09500_, _09499_, _09477_);
  and (_09501_, _09500_, _34789_);
  and (_09502_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_09503_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_09504_, _09503_, _09502_);
  and (_09505_, _09504_, _34581_);
  and (_09506_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_09507_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_09508_, _09507_, _09506_);
  and (_09509_, _09508_, _34796_);
  or (_09510_, _09509_, _09505_);
  and (_09511_, _09510_, _34772_);
  and (_09512_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_09513_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_09514_, _09513_, _09512_);
  and (_09515_, _09514_, _34581_);
  and (_09516_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_09517_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_09518_, _09517_, _09516_);
  and (_09519_, _09518_, _34796_);
  or (_09520_, _09519_, _09515_);
  and (_09521_, _09520_, _34790_);
  or (_09522_, _09521_, _09511_);
  and (_09523_, _09522_, _34803_);
  or (_09524_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_09525_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_09526_, _09525_, _09524_);
  and (_09527_, _09526_, _34581_);
  or (_09528_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_09529_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_09530_, _09529_, _09528_);
  and (_09531_, _09530_, _34796_);
  or (_09532_, _09531_, _09527_);
  and (_09533_, _09532_, _34772_);
  or (_09534_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_09535_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_09536_, _09535_, _09534_);
  and (_09537_, _09536_, _34581_);
  or (_09538_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_09539_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_09540_, _09539_, _09538_);
  and (_09541_, _09540_, _34796_);
  or (_09542_, _09541_, _09537_);
  and (_09543_, _09542_, _34790_);
  or (_09544_, _09543_, _09533_);
  and (_09545_, _09544_, _34719_);
  or (_09546_, _09545_, _09523_);
  and (_09547_, _09546_, _34700_);
  or (_09548_, _09547_, _09501_);
  and (_09549_, _09548_, _34638_);
  or (_09550_, _09549_, _09455_);
  or (_09551_, _09550_, _34692_);
  and (_09552_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_09553_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_09554_, _09553_, _09552_);
  and (_09555_, _09554_, _34581_);
  and (_09556_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_09557_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_09558_, _09557_, _09556_);
  and (_09559_, _09558_, _34796_);
  or (_09560_, _09559_, _09555_);
  or (_09561_, _09560_, _34790_);
  and (_09562_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_09563_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_09564_, _09563_, _09562_);
  and (_09565_, _09564_, _34581_);
  and (_09566_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_09567_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_09568_, _09567_, _09566_);
  and (_09569_, _09568_, _34796_);
  or (_09570_, _09569_, _09565_);
  or (_09571_, _09570_, _34772_);
  and (_09572_, _09571_, _34803_);
  and (_09573_, _09572_, _09561_);
  or (_09574_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_09575_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_09576_, _09575_, _34796_);
  and (_09577_, _09576_, _09574_);
  or (_09578_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_09579_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_09580_, _09579_, _34581_);
  and (_09581_, _09580_, _09578_);
  or (_09582_, _09581_, _09577_);
  or (_09583_, _09582_, _34790_);
  or (_09584_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_09585_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_09586_, _09585_, _34796_);
  and (_09587_, _09586_, _09584_);
  or (_09588_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_09589_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_09590_, _09589_, _34581_);
  and (_09591_, _09590_, _09588_);
  or (_09592_, _09591_, _09587_);
  or (_09593_, _09592_, _34772_);
  and (_09594_, _09593_, _34719_);
  and (_09595_, _09594_, _09583_);
  or (_09596_, _09595_, _09573_);
  and (_09597_, _09596_, _34789_);
  and (_09598_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_09599_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_09600_, _09599_, _09598_);
  and (_09601_, _09600_, _34581_);
  and (_09602_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_09603_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_09604_, _09603_, _09602_);
  and (_09605_, _09604_, _34796_);
  or (_09606_, _09605_, _09601_);
  or (_09607_, _09606_, _34790_);
  and (_09608_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_09609_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_09610_, _09609_, _09608_);
  and (_09611_, _09610_, _34581_);
  and (_09612_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_09613_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_09614_, _09613_, _09612_);
  and (_09615_, _09614_, _34796_);
  or (_09616_, _09615_, _09611_);
  or (_09617_, _09616_, _34772_);
  and (_09618_, _09617_, _34803_);
  and (_09619_, _09618_, _09607_);
  or (_09620_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_09621_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_09622_, _09621_, _09620_);
  and (_09623_, _09622_, _34581_);
  or (_09624_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_09625_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_09626_, _09625_, _09624_);
  and (_09627_, _09626_, _34796_);
  or (_09628_, _09627_, _09623_);
  or (_09629_, _09628_, _34790_);
  or (_09630_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_09631_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_09632_, _09631_, _09630_);
  and (_09633_, _09632_, _34581_);
  or (_09634_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_09635_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_09636_, _09635_, _09634_);
  and (_09637_, _09636_, _34796_);
  or (_09638_, _09637_, _09633_);
  or (_09639_, _09638_, _34772_);
  and (_09640_, _09639_, _34719_);
  and (_09641_, _09640_, _09629_);
  or (_09642_, _09641_, _09619_);
  and (_09643_, _09642_, _34700_);
  or (_09644_, _09643_, _09597_);
  and (_09645_, _09644_, _34840_);
  or (_09646_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_09647_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_09648_, _09647_, _09646_);
  and (_09649_, _09648_, _34581_);
  or (_09650_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_09651_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_09652_, _09651_, _09650_);
  and (_09653_, _09652_, _34796_);
  or (_09654_, _09653_, _09649_);
  and (_09655_, _09654_, _34790_);
  or (_09656_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_09657_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_09658_, _09657_, _09656_);
  and (_09659_, _09658_, _34581_);
  or (_09660_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_09661_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_09662_, _09661_, _09660_);
  and (_09663_, _09662_, _34796_);
  or (_09664_, _09663_, _09659_);
  and (_09665_, _09664_, _34772_);
  or (_09666_, _09665_, _09655_);
  and (_09667_, _09666_, _34719_);
  and (_09668_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_09669_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_09670_, _09669_, _09668_);
  and (_09671_, _09670_, _34581_);
  and (_09672_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_09673_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_09674_, _09673_, _09672_);
  and (_09675_, _09674_, _34796_);
  or (_09676_, _09675_, _09671_);
  and (_09677_, _09676_, _34790_);
  and (_09678_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_09679_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_09680_, _09679_, _09678_);
  and (_09681_, _09680_, _34581_);
  and (_09682_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_09683_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_09684_, _09683_, _09682_);
  and (_09685_, _09684_, _34796_);
  or (_09686_, _09685_, _09681_);
  and (_09687_, _09686_, _34772_);
  or (_09688_, _09687_, _09677_);
  and (_09689_, _09688_, _34803_);
  or (_09690_, _09689_, _09667_);
  and (_09691_, _09690_, _34700_);
  or (_09692_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_09693_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_09694_, _09693_, _34796_);
  and (_09695_, _09694_, _09692_);
  or (_09696_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_09697_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_09698_, _09697_, _34581_);
  and (_09699_, _09698_, _09696_);
  or (_09700_, _09699_, _09695_);
  and (_09701_, _09700_, _34790_);
  or (_09702_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_09703_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_09704_, _09703_, _34796_);
  and (_09705_, _09704_, _09702_);
  or (_09706_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_09707_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_09708_, _09707_, _34581_);
  and (_09709_, _09708_, _09706_);
  or (_09710_, _09709_, _09705_);
  and (_09711_, _09710_, _34772_);
  or (_09712_, _09711_, _09701_);
  and (_09713_, _09712_, _34719_);
  and (_09714_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_09715_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_09716_, _09715_, _09714_);
  and (_09717_, _09716_, _34581_);
  and (_09718_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_09719_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_09720_, _09719_, _09718_);
  and (_09721_, _09720_, _34796_);
  or (_09722_, _09721_, _09717_);
  and (_09723_, _09722_, _34790_);
  and (_09724_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_09725_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_09726_, _09725_, _09724_);
  and (_09727_, _09726_, _34581_);
  and (_09728_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_09729_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_09730_, _09729_, _09728_);
  and (_09731_, _09730_, _34796_);
  or (_09732_, _09731_, _09727_);
  and (_09733_, _09732_, _34772_);
  or (_09734_, _09733_, _09723_);
  and (_09735_, _09734_, _34803_);
  or (_09736_, _09735_, _09713_);
  and (_09737_, _09736_, _34789_);
  or (_09738_, _09737_, _09691_);
  and (_09739_, _09738_, _34638_);
  or (_09740_, _09739_, _09645_);
  or (_09741_, _09740_, _34985_);
  and (_09742_, _09741_, _09551_);
  or (_09743_, _09742_, _34346_);
  and (_09744_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_09745_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_09746_, _09745_, _09744_);
  and (_09747_, _09746_, _34581_);
  and (_09748_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_09749_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_09750_, _09749_, _09748_);
  and (_09751_, _09750_, _34796_);
  or (_09752_, _09751_, _09747_);
  and (_09753_, _09752_, _34772_);
  and (_09754_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_09755_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_09756_, _09755_, _09754_);
  and (_09757_, _09756_, _34581_);
  and (_09758_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_09759_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_09760_, _09759_, _09758_);
  and (_09761_, _09760_, _34796_);
  or (_09762_, _09761_, _09757_);
  and (_09763_, _09762_, _34790_);
  or (_09764_, _09763_, _09753_);
  and (_09765_, _09764_, _34803_);
  or (_09766_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_09767_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_09768_, _09767_, _34796_);
  and (_09769_, _09768_, _09766_);
  or (_09770_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_09771_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_09772_, _09771_, _34581_);
  and (_09773_, _09772_, _09770_);
  or (_09774_, _09773_, _09769_);
  and (_09775_, _09774_, _34772_);
  or (_09776_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_09777_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_09778_, _09777_, _34796_);
  and (_09779_, _09778_, _09776_);
  or (_09780_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_09781_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_09782_, _09781_, _34581_);
  and (_09783_, _09782_, _09780_);
  or (_09784_, _09783_, _09779_);
  and (_09785_, _09784_, _34790_);
  or (_09786_, _09785_, _09775_);
  and (_09787_, _09786_, _34719_);
  or (_09788_, _09787_, _09765_);
  and (_09789_, _09788_, _34789_);
  and (_09790_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_09791_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_09792_, _09791_, _09790_);
  and (_09793_, _09792_, _34581_);
  and (_09794_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_09795_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_09796_, _09795_, _09794_);
  and (_09797_, _09796_, _34796_);
  or (_09798_, _09797_, _09793_);
  and (_09799_, _09798_, _34772_);
  and (_09800_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_09801_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_09802_, _09801_, _09800_);
  and (_09803_, _09802_, _34581_);
  and (_09804_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_09805_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_09806_, _09805_, _09804_);
  and (_09807_, _09806_, _34796_);
  or (_09808_, _09807_, _09803_);
  and (_09809_, _09808_, _34790_);
  or (_09810_, _09809_, _09799_);
  and (_09811_, _09810_, _34803_);
  or (_09812_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_09813_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_09814_, _09813_, _09812_);
  and (_09815_, _09814_, _34581_);
  or (_09816_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_09817_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_09818_, _09817_, _09816_);
  and (_09819_, _09818_, _34796_);
  or (_09820_, _09819_, _09815_);
  and (_09821_, _09820_, _34772_);
  or (_09822_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_09823_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_09824_, _09823_, _09822_);
  and (_09825_, _09824_, _34581_);
  or (_09826_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_09827_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_09828_, _09827_, _09826_);
  and (_09829_, _09828_, _34796_);
  or (_09830_, _09829_, _09825_);
  and (_09831_, _09830_, _34790_);
  or (_09832_, _09831_, _09821_);
  and (_09833_, _09832_, _34719_);
  or (_09834_, _09833_, _09811_);
  and (_09835_, _09834_, _34700_);
  or (_09836_, _09835_, _09789_);
  and (_09837_, _09836_, _34638_);
  and (_09838_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_09839_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_09840_, _09839_, _09838_);
  and (_09841_, _09840_, _34581_);
  and (_09842_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_09843_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_09844_, _09843_, _09842_);
  and (_09845_, _09844_, _34796_);
  or (_09846_, _09845_, _09841_);
  or (_09847_, _09846_, _34790_);
  and (_09848_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_09849_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_09850_, _09849_, _09848_);
  and (_09851_, _09850_, _34581_);
  and (_09852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_09853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_09854_, _09853_, _09852_);
  and (_09855_, _09854_, _34796_);
  or (_09856_, _09855_, _09851_);
  or (_09857_, _09856_, _34772_);
  and (_09858_, _09857_, _34803_);
  and (_09859_, _09858_, _09847_);
  or (_09860_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_09861_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_09862_, _09861_, _09860_);
  and (_09863_, _09862_, _34581_);
  or (_09864_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_09865_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_09866_, _09865_, _09864_);
  and (_09867_, _09866_, _34796_);
  or (_09868_, _09867_, _09863_);
  or (_09869_, _09868_, _34790_);
  or (_09870_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_09871_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_09872_, _09871_, _09870_);
  and (_09873_, _09872_, _34581_);
  or (_09874_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_09875_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_09876_, _09875_, _09874_);
  and (_09877_, _09876_, _34796_);
  or (_09878_, _09877_, _09873_);
  or (_09879_, _09878_, _34772_);
  and (_09880_, _09879_, _34719_);
  and (_09881_, _09880_, _09869_);
  or (_09882_, _09881_, _09859_);
  and (_09883_, _09882_, _34700_);
  and (_09884_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_09885_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_09886_, _09885_, _09884_);
  and (_09887_, _09886_, _34581_);
  and (_09888_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_09889_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_09890_, _09889_, _09888_);
  and (_09891_, _09890_, _34796_);
  or (_09892_, _09891_, _09887_);
  or (_09893_, _09892_, _34790_);
  and (_09894_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_09895_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_09896_, _09895_, _09894_);
  and (_09897_, _09896_, _34581_);
  and (_09898_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_09899_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_09900_, _09899_, _09898_);
  and (_09901_, _09900_, _34796_);
  or (_09902_, _09901_, _09897_);
  or (_09903_, _09902_, _34772_);
  and (_09904_, _09903_, _34803_);
  and (_09905_, _09904_, _09893_);
  or (_09906_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_09907_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_09908_, _09907_, _34796_);
  and (_09909_, _09908_, _09906_);
  or (_09910_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_09911_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_09912_, _09911_, _34581_);
  and (_09913_, _09912_, _09910_);
  or (_09914_, _09913_, _09909_);
  or (_09915_, _09914_, _34790_);
  or (_09916_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_09917_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_09918_, _09917_, _34796_);
  and (_09919_, _09918_, _09916_);
  or (_09920_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_09921_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_09922_, _09921_, _34581_);
  and (_09923_, _09922_, _09920_);
  or (_09924_, _09923_, _09919_);
  or (_09925_, _09924_, _34772_);
  and (_09926_, _09925_, _34719_);
  and (_09927_, _09926_, _09915_);
  or (_09928_, _09927_, _09905_);
  and (_09929_, _09928_, _34789_);
  or (_09930_, _09929_, _09883_);
  and (_09931_, _09930_, _34840_);
  or (_09932_, _09931_, _09837_);
  or (_09933_, _09932_, _34692_);
  and (_09934_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_09935_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_09936_, _09935_, _09934_);
  and (_09937_, _09936_, _34796_);
  and (_09938_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_09939_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_09940_, _09939_, _09938_);
  and (_09941_, _09940_, _34581_);
  or (_09942_, _09941_, _09937_);
  or (_09943_, _09942_, _34790_);
  and (_09944_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_09945_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_09946_, _09945_, _09944_);
  and (_09947_, _09946_, _34796_);
  and (_09948_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_09949_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_09950_, _09949_, _09948_);
  and (_09951_, _09950_, _34581_);
  or (_09952_, _09951_, _09947_);
  or (_09953_, _09952_, _34772_);
  and (_09954_, _09953_, _34803_);
  and (_09955_, _09954_, _09943_);
  or (_09956_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_09957_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_09958_, _09957_, _34581_);
  and (_09959_, _09958_, _09956_);
  or (_09960_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_09961_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_09962_, _09961_, _34796_);
  and (_09963_, _09962_, _09960_);
  or (_09964_, _09963_, _09959_);
  or (_09965_, _09964_, _34790_);
  or (_09966_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_09967_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_09968_, _09967_, _34581_);
  and (_09969_, _09968_, _09966_);
  or (_09970_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_09971_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_09972_, _09971_, _34796_);
  and (_09973_, _09972_, _09970_);
  or (_09974_, _09973_, _09969_);
  or (_09975_, _09974_, _34772_);
  and (_09976_, _09975_, _34719_);
  and (_09977_, _09976_, _09965_);
  or (_09978_, _09977_, _09955_);
  and (_09979_, _09978_, _34789_);
  and (_09980_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_09981_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_09982_, _09981_, _34581_);
  or (_09983_, _09982_, _09980_);
  and (_09984_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_09985_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_09986_, _09985_, _34796_);
  or (_09987_, _09986_, _09984_);
  and (_09988_, _09987_, _09983_);
  or (_09989_, _09988_, _34790_);
  and (_09990_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_09991_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_09992_, _09991_, _34581_);
  or (_09993_, _09992_, _09990_);
  and (_09994_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_09995_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_09996_, _09995_, _34796_);
  or (_09997_, _09996_, _09994_);
  and (_09998_, _09997_, _09993_);
  or (_09999_, _09998_, _34772_);
  and (_10000_, _09999_, _34803_);
  and (_10001_, _10000_, _09989_);
  or (_10002_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_10003_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_10004_, _10003_, _10002_);
  or (_10005_, _10004_, _34796_);
  or (_10006_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_10007_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_10008_, _10007_, _10006_);
  or (_10009_, _10008_, _34581_);
  and (_10010_, _10009_, _10005_);
  or (_10011_, _10010_, _34790_);
  or (_10012_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_10013_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_10014_, _10013_, _10012_);
  or (_10015_, _10014_, _34796_);
  or (_10016_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_10017_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_10018_, _10017_, _10016_);
  or (_10019_, _10018_, _34581_);
  and (_10020_, _10019_, _10015_);
  or (_10021_, _10020_, _34772_);
  and (_10022_, _10021_, _34719_);
  and (_10023_, _10022_, _10011_);
  or (_10024_, _10023_, _10001_);
  and (_10025_, _10024_, _34700_);
  or (_10026_, _10025_, _09979_);
  and (_10027_, _10026_, _34840_);
  and (_10028_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_10029_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_10030_, _10029_, _10028_);
  and (_10031_, _10030_, _34581_);
  and (_10032_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_10033_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_10034_, _10033_, _10032_);
  and (_10035_, _10034_, _34796_);
  or (_10036_, _10035_, _10031_);
  and (_10037_, _10036_, _34772_);
  and (_10038_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_10039_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_10040_, _10039_, _10038_);
  and (_10041_, _10040_, _34581_);
  and (_10042_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_10043_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_10044_, _10043_, _10042_);
  and (_10045_, _10044_, _34796_);
  or (_10046_, _10045_, _10041_);
  and (_10047_, _10046_, _34790_);
  or (_10048_, _10047_, _10037_);
  and (_10049_, _10048_, _34803_);
  or (_10050_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_10051_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_10052_, _10051_, _10050_);
  and (_10053_, _10052_, _34581_);
  or (_10054_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_10055_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_10056_, _10055_, _10054_);
  and (_10057_, _10056_, _34796_);
  or (_10058_, _10057_, _10053_);
  and (_10059_, _10058_, _34772_);
  or (_10060_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_10061_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_10062_, _10061_, _10060_);
  and (_10063_, _10062_, _34581_);
  or (_10064_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_10065_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_10066_, _10065_, _10064_);
  and (_10067_, _10066_, _34796_);
  or (_10068_, _10067_, _10063_);
  and (_10069_, _10068_, _34790_);
  or (_10070_, _10069_, _10059_);
  and (_10071_, _10070_, _34719_);
  or (_10072_, _10071_, _10049_);
  and (_10073_, _10072_, _34700_);
  and (_10074_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  and (_10075_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_10076_, _10075_, _10074_);
  and (_10077_, _10076_, _34581_);
  and (_10078_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and (_10079_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_10080_, _10079_, _10078_);
  and (_10081_, _10080_, _34796_);
  or (_10082_, _10081_, _10077_);
  and (_10083_, _10082_, _34772_);
  and (_10084_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  and (_10085_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_10086_, _10085_, _10084_);
  and (_10087_, _10086_, _34581_);
  and (_10088_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and (_10089_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_10090_, _10089_, _10088_);
  and (_10091_, _10090_, _34796_);
  or (_10092_, _10091_, _10087_);
  and (_10093_, _10092_, _34790_);
  or (_10094_, _10093_, _10083_);
  and (_10095_, _10094_, _34803_);
  or (_10096_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_10097_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and (_10098_, _10097_, _10096_);
  and (_10099_, _10098_, _34581_);
  or (_10100_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_10101_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and (_10102_, _10101_, _10100_);
  and (_10103_, _10102_, _34796_);
  or (_10104_, _10103_, _10099_);
  and (_10105_, _10104_, _34772_);
  or (_10106_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_10107_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and (_10108_, _10107_, _10106_);
  and (_10109_, _10108_, _34581_);
  or (_10110_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_10111_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and (_10112_, _10111_, _10110_);
  and (_10113_, _10112_, _34796_);
  or (_10114_, _10113_, _10109_);
  and (_10115_, _10114_, _34790_);
  or (_10116_, _10115_, _10105_);
  and (_10117_, _10116_, _34719_);
  or (_10118_, _10117_, _10095_);
  and (_10119_, _10118_, _34789_);
  or (_10120_, _10119_, _10073_);
  and (_10121_, _10120_, _34638_);
  or (_10122_, _10121_, _10027_);
  or (_10123_, _10122_, _34985_);
  and (_10124_, _10123_, _09933_);
  or (_10125_, _10124_, _35178_);
  and (_10126_, _10125_, _09743_);
  or (_10127_, _10126_, _34788_);
  or (_10128_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_10129_, _10128_, _38997_);
  and (_38984_[5], _10129_, _10127_);
  and (_10130_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_10131_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_10132_, _10131_, _10130_);
  and (_10133_, _10132_, _34581_);
  and (_10134_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_10135_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_10136_, _10135_, _10134_);
  and (_10137_, _10136_, _34796_);
  or (_10138_, _10137_, _10133_);
  or (_10139_, _10138_, _34790_);
  and (_10140_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_10141_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_10142_, _10141_, _10140_);
  and (_10143_, _10142_, _34581_);
  and (_10144_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_10145_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_10146_, _10145_, _10144_);
  and (_10147_, _10146_, _34796_);
  or (_10148_, _10147_, _10143_);
  or (_10149_, _10148_, _34772_);
  and (_10150_, _10149_, _34803_);
  and (_10151_, _10150_, _10139_);
  or (_10152_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_10153_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_10154_, _10153_, _10152_);
  and (_10155_, _10154_, _34581_);
  or (_10156_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_10157_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_10158_, _10157_, _10156_);
  and (_10159_, _10158_, _34796_);
  or (_10160_, _10159_, _10155_);
  or (_10161_, _10160_, _34790_);
  or (_10162_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_10163_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_10164_, _10163_, _10162_);
  and (_10165_, _10164_, _34581_);
  or (_10166_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_10167_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_10168_, _10167_, _10166_);
  and (_10169_, _10168_, _34796_);
  or (_10170_, _10169_, _10165_);
  or (_10171_, _10170_, _34772_);
  and (_10172_, _10171_, _34719_);
  and (_10173_, _10172_, _10161_);
  or (_10174_, _10173_, _10151_);
  and (_10175_, _10174_, _34700_);
  and (_10176_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_10177_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_10178_, _10177_, _10176_);
  and (_10179_, _10178_, _34581_);
  and (_10180_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_10181_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_10182_, _10181_, _10180_);
  and (_10183_, _10182_, _34796_);
  or (_10184_, _10183_, _10179_);
  or (_10185_, _10184_, _34790_);
  and (_10186_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_10187_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_10188_, _10187_, _10186_);
  and (_10189_, _10188_, _34581_);
  and (_10190_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_10191_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_10192_, _10191_, _10190_);
  and (_10193_, _10192_, _34796_);
  or (_10194_, _10193_, _10189_);
  or (_10195_, _10194_, _34772_);
  and (_10196_, _10195_, _34803_);
  and (_10197_, _10196_, _10185_);
  or (_10198_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_10199_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_10200_, _10199_, _34796_);
  and (_10201_, _10200_, _10198_);
  or (_10202_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_10203_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_10204_, _10203_, _34581_);
  and (_10205_, _10204_, _10202_);
  or (_10206_, _10205_, _10201_);
  or (_10207_, _10206_, _34790_);
  or (_10208_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_10209_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_10210_, _10209_, _34796_);
  and (_10211_, _10210_, _10208_);
  or (_10212_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_10213_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_10214_, _10213_, _34581_);
  and (_10215_, _10214_, _10212_);
  or (_10216_, _10215_, _10211_);
  or (_10217_, _10216_, _34772_);
  and (_10218_, _10217_, _34719_);
  and (_10219_, _10218_, _10207_);
  or (_10220_, _10219_, _10197_);
  and (_10221_, _10220_, _34789_);
  or (_10222_, _10221_, _10175_);
  and (_10223_, _10222_, _34840_);
  and (_10224_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_10225_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _34581_);
  and (_10228_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_10229_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_10230_, _10229_, _10228_);
  and (_10231_, _10230_, _34796_);
  or (_10232_, _10231_, _10227_);
  and (_10233_, _10232_, _34772_);
  and (_10234_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_10235_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_10236_, _10235_, _10234_);
  and (_10237_, _10236_, _34581_);
  and (_10238_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_10239_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_10240_, _10239_, _10238_);
  and (_10241_, _10240_, _34796_);
  or (_10242_, _10241_, _10237_);
  and (_10243_, _10242_, _34790_);
  or (_10244_, _10243_, _10233_);
  and (_10245_, _10244_, _34803_);
  or (_10246_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_10247_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_10248_, _10247_, _34796_);
  and (_10249_, _10248_, _10246_);
  or (_10250_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_10251_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_10252_, _10251_, _34581_);
  and (_10253_, _10252_, _10250_);
  or (_10254_, _10253_, _10249_);
  and (_10255_, _10254_, _34772_);
  or (_10256_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_10257_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_10258_, _10257_, _34796_);
  and (_10259_, _10258_, _10256_);
  or (_10260_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_10261_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_10262_, _10261_, _34581_);
  and (_10263_, _10262_, _10260_);
  or (_10264_, _10263_, _10259_);
  and (_10265_, _10264_, _34790_);
  or (_10266_, _10265_, _10255_);
  and (_10267_, _10266_, _34719_);
  or (_10268_, _10267_, _10245_);
  and (_10269_, _10268_, _34789_);
  and (_10270_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_10271_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_10272_, _10271_, _10270_);
  and (_10273_, _10272_, _34581_);
  and (_10274_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_10275_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_10276_, _10275_, _10274_);
  and (_10277_, _10276_, _34796_);
  or (_10278_, _10277_, _10273_);
  and (_10279_, _10278_, _34772_);
  and (_10280_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_10281_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_10282_, _10281_, _10280_);
  and (_10283_, _10282_, _34581_);
  and (_10284_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_10285_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_10286_, _10285_, _10284_);
  and (_10287_, _10286_, _34796_);
  or (_10288_, _10287_, _10283_);
  and (_10289_, _10288_, _34790_);
  or (_10290_, _10289_, _10279_);
  and (_10291_, _10290_, _34803_);
  or (_10292_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_10293_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_10294_, _10293_, _10292_);
  and (_10295_, _10294_, _34581_);
  or (_10296_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_10297_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_10298_, _10297_, _10296_);
  and (_10299_, _10298_, _34796_);
  or (_10300_, _10299_, _10295_);
  and (_10301_, _10300_, _34772_);
  or (_10302_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_10303_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_10304_, _10303_, _10302_);
  and (_10305_, _10304_, _34581_);
  or (_10306_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_10307_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_10308_, _10307_, _10306_);
  and (_10309_, _10308_, _34796_);
  or (_10310_, _10309_, _10305_);
  and (_10311_, _10310_, _34790_);
  or (_10312_, _10311_, _10301_);
  and (_10313_, _10312_, _34719_);
  or (_10314_, _10313_, _10291_);
  and (_10315_, _10314_, _34700_);
  or (_10316_, _10315_, _10269_);
  and (_10317_, _10316_, _34638_);
  or (_10318_, _10317_, _10223_);
  or (_10319_, _10318_, _34692_);
  and (_10320_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_10321_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_10322_, _10321_, _10320_);
  and (_10323_, _10322_, _34581_);
  and (_10324_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_10325_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_10326_, _10325_, _10324_);
  and (_10327_, _10326_, _34796_);
  or (_10328_, _10327_, _10323_);
  or (_10329_, _10328_, _34790_);
  and (_10330_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_10331_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_10332_, _10331_, _10330_);
  and (_10333_, _10332_, _34581_);
  and (_10334_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_10335_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_10336_, _10335_, _10334_);
  and (_10337_, _10336_, _34796_);
  or (_10338_, _10337_, _10333_);
  or (_10339_, _10338_, _34772_);
  and (_10340_, _10339_, _34803_);
  and (_10341_, _10340_, _10329_);
  or (_10342_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_10343_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_10344_, _10343_, _34796_);
  and (_10345_, _10344_, _10342_);
  or (_10346_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_10347_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_10348_, _10347_, _34581_);
  and (_10349_, _10348_, _10346_);
  or (_10350_, _10349_, _10345_);
  or (_10351_, _10350_, _34790_);
  or (_10352_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_10353_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_10354_, _10353_, _34796_);
  and (_10355_, _10354_, _10352_);
  or (_10356_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_10357_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_10358_, _10357_, _34581_);
  and (_10359_, _10358_, _10356_);
  or (_10360_, _10359_, _10355_);
  or (_10361_, _10360_, _34772_);
  and (_10362_, _10361_, _34719_);
  and (_10363_, _10362_, _10351_);
  or (_10364_, _10363_, _10341_);
  and (_10365_, _10364_, _34789_);
  and (_10366_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_10367_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_10368_, _10367_, _10366_);
  and (_10369_, _10368_, _34581_);
  and (_10370_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_10371_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_10372_, _10371_, _10370_);
  and (_10373_, _10372_, _34796_);
  or (_10374_, _10373_, _10369_);
  or (_10375_, _10374_, _34790_);
  and (_10376_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_10377_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_10378_, _10377_, _10376_);
  and (_10379_, _10378_, _34581_);
  and (_10380_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_10381_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_10382_, _10381_, _10380_);
  and (_10383_, _10382_, _34796_);
  or (_10384_, _10383_, _10379_);
  or (_10385_, _10384_, _34772_);
  and (_10386_, _10385_, _34803_);
  and (_10387_, _10386_, _10375_);
  or (_10388_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_10389_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_10390_, _10389_, _10388_);
  and (_10391_, _10390_, _34581_);
  or (_10392_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_10393_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_10394_, _10393_, _10392_);
  and (_10395_, _10394_, _34796_);
  or (_10396_, _10395_, _10391_);
  or (_10397_, _10396_, _34790_);
  or (_10398_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_10399_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_10400_, _10399_, _10398_);
  and (_10401_, _10400_, _34581_);
  or (_10402_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_10403_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_10404_, _10403_, _10402_);
  and (_10405_, _10404_, _34796_);
  or (_10406_, _10405_, _10401_);
  or (_10407_, _10406_, _34772_);
  and (_10408_, _10407_, _34719_);
  and (_10409_, _10408_, _10397_);
  or (_10410_, _10409_, _10387_);
  and (_10411_, _10410_, _34700_);
  or (_10412_, _10411_, _10365_);
  and (_10413_, _10412_, _34840_);
  or (_10414_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_10415_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_10416_, _10415_, _10414_);
  and (_10417_, _10416_, _34581_);
  or (_10418_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_10419_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_10420_, _10419_, _10418_);
  and (_10421_, _10420_, _34796_);
  or (_10422_, _10421_, _10417_);
  and (_10423_, _10422_, _34790_);
  or (_10424_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_10425_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_10426_, _10425_, _10424_);
  and (_10427_, _10426_, _34581_);
  or (_10428_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_10429_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_10430_, _10429_, _10428_);
  and (_10431_, _10430_, _34796_);
  or (_10432_, _10431_, _10427_);
  and (_10433_, _10432_, _34772_);
  or (_10434_, _10433_, _10423_);
  and (_10435_, _10434_, _34719_);
  and (_10436_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_10437_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_10438_, _10437_, _10436_);
  and (_10439_, _10438_, _34581_);
  and (_10440_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_10441_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_10442_, _10441_, _10440_);
  and (_10443_, _10442_, _34796_);
  or (_10444_, _10443_, _10439_);
  and (_10445_, _10444_, _34790_);
  and (_10446_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_10447_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_10448_, _10447_, _10446_);
  and (_10449_, _10448_, _34581_);
  and (_10450_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_10451_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_10452_, _10451_, _10450_);
  and (_10453_, _10452_, _34796_);
  or (_10454_, _10453_, _10449_);
  and (_10455_, _10454_, _34772_);
  or (_10456_, _10455_, _10445_);
  and (_10457_, _10456_, _34803_);
  or (_10458_, _10457_, _10435_);
  and (_10459_, _10458_, _34700_);
  or (_10460_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_10461_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_10462_, _10461_, _34796_);
  and (_10463_, _10462_, _10460_);
  or (_10464_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_10465_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_10466_, _10465_, _34581_);
  and (_10467_, _10466_, _10464_);
  or (_10468_, _10467_, _10463_);
  and (_10469_, _10468_, _34790_);
  or (_10470_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_10471_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_10472_, _10471_, _34796_);
  and (_10473_, _10472_, _10470_);
  or (_10474_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_10475_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_10476_, _10475_, _34581_);
  and (_10477_, _10476_, _10474_);
  or (_10478_, _10477_, _10473_);
  and (_10479_, _10478_, _34772_);
  or (_10480_, _10479_, _10469_);
  and (_10481_, _10480_, _34719_);
  and (_10482_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_10483_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_10484_, _10483_, _10482_);
  and (_10485_, _10484_, _34581_);
  and (_10486_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_10487_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_10488_, _10487_, _10486_);
  and (_10489_, _10488_, _34796_);
  or (_10490_, _10489_, _10485_);
  and (_10491_, _10490_, _34790_);
  and (_10492_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_10493_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_10494_, _10493_, _10492_);
  and (_10495_, _10494_, _34581_);
  and (_10496_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_10497_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_10498_, _10497_, _10496_);
  and (_10499_, _10498_, _34796_);
  or (_10500_, _10499_, _10495_);
  and (_10501_, _10500_, _34772_);
  or (_10502_, _10501_, _10491_);
  and (_10503_, _10502_, _34803_);
  or (_10504_, _10503_, _10481_);
  and (_10505_, _10504_, _34789_);
  or (_10506_, _10505_, _10459_);
  and (_10507_, _10506_, _34638_);
  or (_10508_, _10507_, _10413_);
  or (_10509_, _10508_, _34985_);
  and (_10510_, _10509_, _10319_);
  or (_10511_, _10510_, _34346_);
  and (_10512_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_10513_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_10514_, _10513_, _10512_);
  and (_10515_, _10514_, _34581_);
  and (_10516_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_10517_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_10518_, _10517_, _10516_);
  and (_10519_, _10518_, _34796_);
  or (_10520_, _10519_, _10515_);
  or (_10521_, _10520_, _34790_);
  and (_10522_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_10523_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_10524_, _10523_, _10522_);
  and (_10525_, _10524_, _34581_);
  and (_10526_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_10527_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_10528_, _10527_, _10526_);
  and (_10529_, _10528_, _34796_);
  or (_10530_, _10529_, _10525_);
  or (_10531_, _10530_, _34772_);
  and (_10532_, _10531_, _34803_);
  and (_10533_, _10532_, _10521_);
  or (_10534_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_10535_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_10536_, _10535_, _10534_);
  and (_10537_, _10536_, _34581_);
  or (_10538_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_10539_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_10540_, _10539_, _10538_);
  and (_10541_, _10540_, _34796_);
  or (_10542_, _10541_, _10537_);
  or (_10543_, _10542_, _34790_);
  or (_10544_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_10545_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_10546_, _10545_, _10544_);
  and (_10547_, _10546_, _34581_);
  or (_10548_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_10549_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_10550_, _10549_, _10548_);
  and (_10551_, _10550_, _34796_);
  or (_10552_, _10551_, _10547_);
  or (_10553_, _10552_, _34772_);
  and (_10554_, _10553_, _34719_);
  and (_10555_, _10554_, _10543_);
  or (_10556_, _10555_, _10533_);
  and (_10557_, _10556_, _34700_);
  and (_10558_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_10559_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_10560_, _10559_, _10558_);
  and (_10561_, _10560_, _34581_);
  and (_10562_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_10563_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_10564_, _10563_, _10562_);
  and (_10565_, _10564_, _34796_);
  or (_10566_, _10565_, _10561_);
  or (_10567_, _10566_, _34790_);
  and (_10568_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_10569_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_10570_, _10569_, _10568_);
  and (_10571_, _10570_, _34581_);
  and (_10572_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_10573_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_10574_, _10573_, _10572_);
  and (_10575_, _10574_, _34796_);
  or (_10576_, _10575_, _10571_);
  or (_10577_, _10576_, _34772_);
  and (_10578_, _10577_, _34803_);
  and (_10579_, _10578_, _10567_);
  or (_10580_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_10581_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_10582_, _10581_, _34796_);
  and (_10583_, _10582_, _10580_);
  or (_10584_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_10585_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_10586_, _10585_, _34581_);
  and (_10587_, _10586_, _10584_);
  or (_10588_, _10587_, _10583_);
  or (_10589_, _10588_, _34790_);
  or (_10590_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_10591_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_10592_, _10591_, _34796_);
  and (_10593_, _10592_, _10590_);
  or (_10594_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_10595_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_10596_, _10595_, _34581_);
  and (_10597_, _10596_, _10594_);
  or (_10598_, _10597_, _10593_);
  or (_10599_, _10598_, _34772_);
  and (_10600_, _10599_, _34719_);
  and (_10601_, _10600_, _10589_);
  or (_10602_, _10601_, _10579_);
  and (_10603_, _10602_, _34789_);
  or (_10604_, _10603_, _10557_);
  and (_10605_, _10604_, _34840_);
  and (_10606_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_10607_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_10608_, _10607_, _10606_);
  and (_10609_, _10608_, _34581_);
  and (_10610_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_10611_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_10612_, _10611_, _10610_);
  and (_10613_, _10612_, _34796_);
  or (_10614_, _10613_, _10609_);
  and (_10615_, _10614_, _34772_);
  and (_10616_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_10617_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_10618_, _10617_, _10616_);
  and (_10619_, _10618_, _34581_);
  and (_10620_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_10621_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_10622_, _10621_, _10620_);
  and (_10623_, _10622_, _34796_);
  or (_10624_, _10623_, _10619_);
  and (_10625_, _10624_, _34790_);
  or (_10626_, _10625_, _10615_);
  and (_10627_, _10626_, _34803_);
  or (_10628_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_10629_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_10630_, _10629_, _34796_);
  and (_10631_, _10630_, _10628_);
  or (_10632_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_10633_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  and (_10634_, _10633_, _34581_);
  and (_10635_, _10634_, _10632_);
  or (_10636_, _10635_, _10631_);
  and (_10637_, _10636_, _34772_);
  or (_10638_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_10639_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  and (_10640_, _10639_, _34796_);
  and (_10641_, _10640_, _10638_);
  or (_10642_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_10643_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_10644_, _10643_, _34581_);
  and (_10645_, _10644_, _10642_);
  or (_10646_, _10645_, _10641_);
  and (_10647_, _10646_, _34790_);
  or (_10648_, _10647_, _10637_);
  and (_10649_, _10648_, _34719_);
  or (_10650_, _10649_, _10627_);
  and (_10651_, _10650_, _34789_);
  and (_10652_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_10653_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_10654_, _10653_, _10652_);
  and (_10655_, _10654_, _34581_);
  and (_10656_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_10657_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_10658_, _10657_, _10656_);
  and (_10659_, _10658_, _34796_);
  or (_10660_, _10659_, _10655_);
  and (_10661_, _10660_, _34772_);
  and (_10662_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_10663_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_10664_, _10663_, _10662_);
  and (_10665_, _10664_, _34581_);
  and (_10666_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_10667_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_10668_, _10667_, _10666_);
  and (_10669_, _10668_, _34796_);
  or (_10670_, _10669_, _10665_);
  and (_10671_, _10670_, _34790_);
  or (_10672_, _10671_, _10661_);
  and (_10673_, _10672_, _34803_);
  or (_10674_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_10675_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_10676_, _10675_, _10674_);
  and (_10677_, _10676_, _34581_);
  or (_10678_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_10679_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_10680_, _10679_, _10678_);
  and (_10681_, _10680_, _34796_);
  or (_10682_, _10681_, _10677_);
  and (_10683_, _10682_, _34772_);
  or (_10684_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_10685_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_10686_, _10685_, _10684_);
  and (_10687_, _10686_, _34581_);
  or (_10688_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_10689_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_10690_, _10689_, _10688_);
  and (_10691_, _10690_, _34796_);
  or (_10692_, _10691_, _10687_);
  and (_10693_, _10692_, _34790_);
  or (_10694_, _10693_, _10683_);
  and (_10695_, _10694_, _34719_);
  or (_10696_, _10695_, _10673_);
  and (_10697_, _10696_, _34700_);
  or (_10698_, _10697_, _10651_);
  and (_10699_, _10698_, _34638_);
  or (_10700_, _10699_, _10605_);
  or (_10701_, _10700_, _34692_);
  and (_10702_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_10703_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_10704_, _10703_, _10702_);
  and (_10705_, _10704_, _34581_);
  and (_10706_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_10707_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _34796_);
  or (_10710_, _10709_, _10705_);
  or (_10711_, _10710_, _34790_);
  and (_10712_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_10713_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_10714_, _10713_, _10712_);
  and (_10715_, _10714_, _34581_);
  and (_10716_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_10717_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_10718_, _10717_, _10716_);
  and (_10719_, _10718_, _34796_);
  or (_10720_, _10719_, _10715_);
  or (_10721_, _10720_, _34772_);
  and (_10722_, _10721_, _34803_);
  and (_10723_, _10722_, _10711_);
  or (_10724_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_10725_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_10726_, _10725_, _34796_);
  and (_10727_, _10726_, _10724_);
  or (_10728_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_10729_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_10730_, _10729_, _34581_);
  and (_10731_, _10730_, _10728_);
  or (_10732_, _10731_, _10727_);
  or (_10733_, _10732_, _34790_);
  or (_10734_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_10735_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_10736_, _10735_, _34796_);
  and (_10737_, _10736_, _10734_);
  or (_10738_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_10739_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_10740_, _10739_, _34581_);
  and (_10741_, _10740_, _10738_);
  or (_10742_, _10741_, _10737_);
  or (_10743_, _10742_, _34772_);
  and (_10744_, _10743_, _34719_);
  and (_10745_, _10744_, _10733_);
  or (_10746_, _10745_, _10723_);
  and (_10747_, _10746_, _34789_);
  and (_10748_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_10749_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_10750_, _10749_, _10748_);
  and (_10751_, _10750_, _34581_);
  and (_10752_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_10753_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_10754_, _10753_, _10752_);
  and (_10755_, _10754_, _34796_);
  or (_10756_, _10755_, _10751_);
  or (_10757_, _10756_, _34790_);
  and (_10758_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_10759_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_10760_, _10759_, _10758_);
  and (_10761_, _10760_, _34581_);
  and (_10762_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_10763_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_10764_, _10763_, _10762_);
  and (_10765_, _10764_, _34796_);
  or (_10766_, _10765_, _10761_);
  or (_10767_, _10766_, _34772_);
  and (_10768_, _10767_, _34803_);
  and (_10769_, _10768_, _10757_);
  or (_10770_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_10771_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_10772_, _10771_, _10770_);
  and (_10773_, _10772_, _34581_);
  or (_10774_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_10775_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_10776_, _10775_, _10774_);
  and (_10777_, _10776_, _34796_);
  or (_10778_, _10777_, _10773_);
  or (_10779_, _10778_, _34790_);
  or (_10780_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_10781_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_10782_, _10781_, _10780_);
  and (_10783_, _10782_, _34581_);
  or (_10784_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_10785_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_10786_, _10785_, _10784_);
  and (_10787_, _10786_, _34796_);
  or (_10788_, _10787_, _10783_);
  or (_10789_, _10788_, _34772_);
  and (_10790_, _10789_, _34719_);
  and (_10791_, _10790_, _10779_);
  or (_10792_, _10791_, _10769_);
  and (_10793_, _10792_, _34700_);
  or (_10794_, _10793_, _10747_);
  and (_10795_, _10794_, _34840_);
  or (_10796_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_10797_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_10798_, _10797_, _10796_);
  and (_10799_, _10798_, _34581_);
  or (_10800_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_10801_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_10802_, _10801_, _10800_);
  and (_10803_, _10802_, _34796_);
  or (_10804_, _10803_, _10799_);
  and (_10805_, _10804_, _34790_);
  or (_10806_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_10807_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_10808_, _10807_, _10806_);
  and (_10809_, _10808_, _34581_);
  or (_10810_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_10811_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_10812_, _10811_, _10810_);
  and (_10813_, _10812_, _34796_);
  or (_10814_, _10813_, _10809_);
  and (_10815_, _10814_, _34772_);
  or (_10816_, _10815_, _10805_);
  and (_10817_, _10816_, _34719_);
  and (_10818_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_10819_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_10820_, _10819_, _10818_);
  and (_10821_, _10820_, _34581_);
  and (_10822_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_10823_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_10824_, _10823_, _10822_);
  and (_10825_, _10824_, _34796_);
  or (_10826_, _10825_, _10821_);
  and (_10827_, _10826_, _34790_);
  and (_10828_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_10829_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_10830_, _10829_, _10828_);
  and (_10831_, _10830_, _34581_);
  and (_10832_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_10833_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_10834_, _10833_, _10832_);
  and (_10835_, _10834_, _34796_);
  or (_10836_, _10835_, _10831_);
  and (_10837_, _10836_, _34772_);
  or (_10838_, _10837_, _10827_);
  and (_10839_, _10838_, _34803_);
  or (_10840_, _10839_, _10817_);
  and (_10841_, _10840_, _34700_);
  or (_10842_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_10843_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_10844_, _10843_, _34796_);
  and (_10845_, _10844_, _10842_);
  or (_10846_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_10847_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_10848_, _10847_, _34581_);
  and (_10849_, _10848_, _10846_);
  or (_10850_, _10849_, _10845_);
  and (_10851_, _10850_, _34790_);
  or (_10852_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_10853_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_10854_, _10853_, _34796_);
  and (_10855_, _10854_, _10852_);
  or (_10856_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_10857_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_10858_, _10857_, _34581_);
  and (_10859_, _10858_, _10856_);
  or (_10860_, _10859_, _10855_);
  and (_10861_, _10860_, _34772_);
  or (_10862_, _10861_, _10851_);
  and (_10863_, _10862_, _34719_);
  and (_10864_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_10865_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_10866_, _10865_, _10864_);
  and (_10867_, _10866_, _34581_);
  and (_10868_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_10869_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_10870_, _10869_, _10868_);
  and (_10871_, _10870_, _34796_);
  or (_10872_, _10871_, _10867_);
  and (_10873_, _10872_, _34790_);
  and (_10874_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_10875_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_10876_, _10875_, _10874_);
  and (_10877_, _10876_, _34581_);
  and (_10878_, _34791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_10879_, _34473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_10880_, _10879_, _10878_);
  and (_10881_, _10880_, _34796_);
  or (_10882_, _10881_, _10877_);
  and (_10883_, _10882_, _34772_);
  or (_10884_, _10883_, _10873_);
  and (_10885_, _10884_, _34803_);
  or (_10886_, _10885_, _10863_);
  and (_10887_, _10886_, _34789_);
  or (_10888_, _10887_, _10841_);
  and (_10889_, _10888_, _34638_);
  or (_10890_, _10889_, _10795_);
  or (_10891_, _10890_, _34985_);
  and (_10892_, _10891_, _10701_);
  or (_10893_, _10892_, _35178_);
  and (_10894_, _10893_, _10511_);
  or (_10895_, _10894_, _34788_);
  or (_10896_, _35563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_10897_, _10896_, _38997_);
  and (_38984_[6], _10897_, _10895_);
  nor (_10898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_39040_, _10898_, rst);
  and (_10899_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_10900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_10901_, _10898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_10902_, _10901_, _10900_);
  not (_10903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_10904_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _10903_);
  or (_10905_, _10904_, _10902_);
  nor (_10906_, _10905_, _10899_);
  or (_10907_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_10908_, _10907_, _38997_);
  nor (_39041_, _10908_, _10906_);
  nor (_10909_, _10906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_10910_, _10909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_10911_, _10909_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_10912_, _10911_, _38997_);
  and (_39042_, _10912_, _10910_);
  not (_10913_, rxd_i);
  and (_10914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _10913_);
  nor (_10915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_10916_, _10915_);
  and (_10917_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and (_10918_, _10917_, _10916_);
  and (_10919_, _10918_, _10914_);
  not (_10920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_10921_, _10920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_10922_, _10921_, _10915_);
  or (_10923_, _10922_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or (_10924_, _10923_, _10919_);
  and (_10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _38997_);
  and (_39043_, _10925_, _10924_);
  and (_10926_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_10927_, _10926_, _10916_);
  nor (_10928_, _10915_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_10929_, _10928_, _10920_);
  nor (_10930_, _10929_, _10927_);
  not (_10931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_10932_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _10931_);
  not (_10933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_10934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _10933_);
  and (_10935_, _10934_, _10932_);
  not (_10936_, _10935_);
  or (_10937_, _10936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and (_10938_, _10935_, _10927_);
  and (_10939_, _10927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_10940_, _10939_, _10938_);
  and (_10941_, _10940_, _10937_);
  or (_10942_, _10941_, _10930_);
  and (_10943_, _10915_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_10944_, _10943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not (_10945_, _10944_);
  or (_10946_, _10945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_10947_, _10946_, _10942_);
  nand (_39044_, _10947_, _10925_);
  not (_10948_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not (_10949_, _10927_);
  nor (_10950_, _10920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_10951_, _10950_);
  not (_10952_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_10953_, _10915_, _10952_);
  and (_10954_, _10953_, _10951_);
  and (_10955_, _10954_, _10949_);
  nor (_10956_, _10955_, _10948_);
  and (_10957_, _10955_, rxd_i);
  or (_10958_, _10957_, rst);
  or (_39045_, _10958_, _10956_);
  nor (_10959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_10960_, _10959_, _10932_);
  and (_10961_, _10960_, _10939_);
  nand (_10962_, _10961_, _10913_);
  or (_10963_, _10961_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_10964_, _10963_, _38997_);
  and (_39046_[1], _10964_, _10962_);
  and (_10965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_10966_, _10965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_10967_, _10966_, _10931_);
  and (_10968_, _10967_, _10939_);
  and (_10969_, _10918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_10970_, _10969_, _10939_);
  nor (_10971_, _10966_, _10949_);
  or (_10972_, _10971_, _10970_);
  and (_10973_, _10972_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_10974_, _10973_, _10968_);
  and (_39047_[3], _10974_, _38997_);
  and (_10975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _38997_);
  nand (_10976_, _10975_, _10952_);
  nand (_10977_, _10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand (_39048_[7], _10977_, _10976_);
  and (_10978_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _10952_);
  not (_10979_, _10918_);
  not (_10980_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand (_10981_, _10922_, _10980_);
  and (_10982_, _10981_, _10979_);
  nand (_10983_, _10982_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand (_10984_, _10983_, _10949_);
  or (_10985_, _10935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_10986_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_10987_, _10986_, _10938_);
  and (_10988_, _10987_, _10985_);
  and (_10989_, _10988_, _10984_);
  or (_10990_, _10989_, _10944_);
  nand (_10991_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand (_10992_, _10991_, _10927_);
  or (_10993_, _10992_, _10936_);
  and (_10994_, _10993_, _10945_);
  or (_10995_, _10994_, rxd_i);
  and (_10996_, _10995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_10997_, _10996_, _10990_);
  or (_10998_, _10997_, _10978_);
  and (_39049_[11], _10998_, _38997_);
  and (_10999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_11000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_11001_, _10901_, _11000_);
  or (_11002_, _11001_, _10904_);
  nor (_11003_, _11002_, _10999_);
  or (_11004_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_11005_, _11004_, _38997_);
  nor (_39050_, _11005_, _11003_);
  nor (_11006_, _11003_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_11007_, _11006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_11008_, _11006_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_11009_, _11008_, _38997_);
  and (_39051_, _11009_, _11007_);
  not (_11010_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_11011_, _34233_, _33632_);
  and (_11012_, _34254_, _33662_);
  and (_11013_, _11012_, _11011_);
  and (_11014_, _11013_, _38997_);
  nand (_11015_, _11014_, _11010_);
  and (_11016_, _10943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  not (_11017_, _11016_);
  nor (_11018_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_11019_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_11020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_11021_, _11020_, _11019_);
  and (_11022_, _11021_, _11018_);
  not (_11023_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_11024_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_11025_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_11026_, _11025_, _11024_);
  and (_11027_, _11026_, _11023_);
  and (_11028_, _11027_, _11022_);
  or (_11029_, _11028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  not (_11030_, _11028_);
  or (_11031_, _11030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and (_11032_, _11031_, _11029_);
  or (_11033_, _11032_, _11017_);
  nor (_11034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_11035_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_11036_, _11035_, _11034_);
  and (_11037_, _10916_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_11038_, _11037_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_11039_, _11038_, _11036_);
  not (_11040_, _11039_);
  or (_11041_, _11040_, _11029_);
  and (_11042_, _11036_, _11037_);
  not (_11043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  or (_11044_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _11043_);
  or (_11045_, _11044_, _11042_);
  or (_11046_, _11045_, _11016_);
  and (_11047_, _11046_, _11041_);
  nand (_11048_, _11047_, _11033_);
  nor (_11049_, _11013_, rst);
  nand (_11050_, _11049_, _11048_);
  and (_39052_, _11050_, _11015_);
  nor (_11051_, _11030_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_11052_, _11042_, _11051_);
  and (_11053_, _11028_, _11016_);
  or (_11054_, _11043_, rst);
  nor (_11055_, _11054_, _11053_);
  and (_11056_, _11055_, _11052_);
  or (_39053_, _11056_, _11014_);
  or (_11057_, _11040_, _11051_);
  or (_11058_, _11042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_11059_, _10943_, _11043_);
  and (_11060_, _11059_, _11058_);
  and (_11061_, _11060_, _11057_);
  or (_11062_, _11061_, _11053_);
  and (_39054_, _11062_, _11049_);
  and (_11063_, _11038_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_11064_, _11063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_11065_, _11064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_11066_, _11065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_11067_, _11065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_11068_, _11067_, _11066_);
  and (_39055_[3], _11068_, _11049_);
  nor (_11069_, _11039_, _11016_);
  and (_11070_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_11071_, _11070_, _11049_);
  and (_11072_, _11014_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_39056_[10], _11072_, _11071_);
  not (_11073_, _33644_);
  nor (_11074_, _33571_, _33558_);
  and (_11075_, _11074_, _11073_);
  and (_11076_, _11075_, _33663_);
  and (_11077_, _11076_, _33633_);
  nand (_11078_, _11077_, _34221_);
  or (_11079_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_11080_, _11079_, _38997_);
  and (_39057_[7], _11080_, _11078_);
  and (_11081_, _33630_, _33591_);
  nor (_11082_, _33657_, _33604_);
  and (_11083_, _33661_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_11084_, _11083_, _34706_);
  and (_11085_, _11084_, _11082_);
  and (_11086_, _11085_, _11081_);
  and (_11087_, _11086_, _11075_);
  or (_11088_, _11087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  not (_11089_, _33662_);
  nor (_11090_, _11089_, _33657_);
  and (_11091_, _11090_, _34229_);
  and (_11092_, _11091_, _11011_);
  not (_11093_, _11092_);
  and (_11094_, _11093_, _11088_);
  nand (_11095_, _11087_, _35722_);
  and (_11096_, _11095_, _11094_);
  nor (_11097_, _11093_, _34221_);
  or (_11098_, _11097_, _11096_);
  and (_39058_[7], _11098_, _38997_);
  nor (_11099_, _10944_, _10938_);
  not (_11100_, _11099_);
  nor (_11101_, _10982_, _10927_);
  nor (_11102_, _11101_, _11100_);
  nor (_11103_, _11102_, _10952_);
  or (_11104_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_11105_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _10952_);
  or (_11106_, _11105_, _11099_);
  and (_11107_, _11106_, _38997_);
  and (_39049_[0], _11107_, _11104_);
  or (_11108_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_11109_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _10952_);
  or (_11110_, _11109_, _11099_);
  and (_11111_, _11110_, _38997_);
  and (_39049_[1], _11111_, _11108_);
  or (_11112_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_11113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _10952_);
  or (_11114_, _11113_, _11099_);
  and (_11115_, _11114_, _38997_);
  and (_39049_[2], _11115_, _11112_);
  or (_11116_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_11117_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _10952_);
  or (_11118_, _11117_, _11099_);
  and (_11119_, _11118_, _38997_);
  and (_39049_[3], _11119_, _11116_);
  or (_11120_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_11121_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _10952_);
  or (_11122_, _11121_, _11099_);
  and (_11123_, _11122_, _38997_);
  and (_39049_[4], _11123_, _11120_);
  or (_11124_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_11125_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _10952_);
  or (_11126_, _11125_, _11099_);
  and (_11127_, _11126_, _38997_);
  and (_39049_[5], _11127_, _11124_);
  or (_11128_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_11129_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _10952_);
  or (_11130_, _11129_, _11099_);
  and (_11131_, _11130_, _38997_);
  and (_39049_[6], _11131_, _11128_);
  or (_11132_, _11103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_11133_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _10952_);
  or (_11134_, _11133_, _11099_);
  and (_11135_, _11134_, _38997_);
  and (_39049_[7], _11135_, _11132_);
  nor (_11136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_11137_, _11136_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_11138_, _10936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_11139_, _10935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_11140_, _11139_, _10927_);
  and (_11141_, _11140_, _11138_);
  or (_11142_, _10918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_11143_, _11142_, _10981_);
  and (_11144_, _11143_, _10949_);
  or (_11145_, _11144_, _11141_);
  or (_11146_, _11145_, _10944_);
  or (_11147_, _10945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_11148_, _11147_, _10925_);
  and (_11149_, _11148_, _11146_);
  or (_39049_[8], _11149_, _11137_);
  and (_11150_, _10935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_11151_, _11150_, _10982_);
  or (_11152_, _11151_, _11102_);
  and (_11153_, _11152_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_11154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _10952_);
  nand (_11155_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_11156_, _11155_, _11099_);
  or (_11157_, _11156_, _11154_);
  or (_11158_, _11157_, _11153_);
  and (_39049_[9], _11158_, _38997_);
  not (_11159_, _11103_);
  and (_11160_, _11159_, _10975_);
  or (_11161_, _11151_, _11100_);
  and (_11162_, _10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_11163_, _11162_, _11161_);
  or (_39049_[10], _11163_, _11160_);
  or (_11164_, _10968_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_11165_, _10968_, _10913_);
  and (_11166_, _11165_, _38997_);
  and (_39046_[0], _11166_, _11164_);
  or (_11167_, _10970_, _10933_);
  or (_11168_, _10939_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_11169_, _11168_, _38997_);
  and (_39047_[0], _11169_, _11167_);
  and (_11170_, _10970_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_11171_, _10959_, _10965_);
  and (_11172_, _11171_, _10939_);
  or (_11173_, _11172_, _11170_);
  and (_39047_[1], _11173_, _38997_);
  and (_11174_, _10972_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_11175_, _10965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_11176_, _11175_, _10971_);
  or (_11177_, _11176_, _11174_);
  and (_39047_[2], _11177_, _38997_);
  and (_11178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _10952_);
  and (_11179_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_11180_, _11179_, _11178_);
  and (_39048_[0], _11180_, _38997_);
  and (_11181_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _10952_);
  and (_11182_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_11183_, _11182_, _11181_);
  and (_39048_[1], _11183_, _38997_);
  and (_11184_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _10952_);
  and (_11185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_11186_, _11185_, _11184_);
  and (_39048_[2], _11186_, _38997_);
  and (_11187_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _10952_);
  and (_11188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_11189_, _11188_, _11187_);
  and (_39048_[3], _11189_, _38997_);
  and (_11190_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _10952_);
  and (_11191_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_11192_, _11191_, _11190_);
  and (_39048_[4], _11192_, _38997_);
  and (_11193_, _10925_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_39048_[5], _11193_, _11137_);
  and (_11194_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_11195_, _11194_, _11154_);
  and (_39048_[6], _11195_, _38997_);
  nor (_11196_, _11038_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_11197_, _11196_, _11063_);
  and (_39055_[0], _11197_, _11049_);
  nor (_11198_, _11063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_11199_, _11198_, _11064_);
  and (_39055_[1], _11199_, _11049_);
  nor (_11200_, _11064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_11201_, _11200_, _11065_);
  and (_39055_[2], _11201_, _11049_);
  or (_11202_, _11039_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_11203_, _11040_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_11204_, _11203_, _11202_);
  and (_11205_, _11204_, _11017_);
  and (_11206_, _11028_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_11207_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_11208_, _11207_, _11016_);
  or (_11209_, _11208_, _11205_);
  and (_11210_, _11209_, _11049_);
  nor (_11211_, _10916_, _34148_);
  and (_11212_, _11211_, _11014_);
  or (_39056_[0], _11212_, _11210_);
  not (_11213_, _11069_);
  and (_11214_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_11215_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_11216_, _11215_, _11214_);
  and (_11217_, _11216_, _11049_);
  or (_11218_, _10916_, _34122_);
  nand (_11219_, _10916_, _34148_);
  and (_11220_, _11219_, _11014_);
  and (_11221_, _11220_, _11218_);
  or (_39056_[1], _11221_, _11217_);
  nor (_11222_, _11069_, _11023_);
  and (_11223_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or (_11224_, _11223_, _11222_);
  and (_11225_, _11224_, _11049_);
  or (_11226_, _10916_, _34089_);
  or (_11227_, _10915_, _34122_);
  and (_11228_, _11227_, _11014_);
  and (_11229_, _11228_, _11226_);
  or (_39056_[2], _11229_, _11225_);
  nor (_11230_, _11069_, _11019_);
  and (_11231_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_11232_, _11231_, _11230_);
  and (_11233_, _11232_, _11049_);
  or (_11234_, _10915_, _34089_);
  nand (_11235_, _10915_, _34052_);
  and (_11236_, _11235_, _11014_);
  and (_11237_, _11236_, _11234_);
  or (_39056_[3], _11237_, _11233_);
  and (_11238_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_11239_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or (_11240_, _11239_, _11238_);
  and (_11241_, _11240_, _11049_);
  nand (_11242_, _10916_, _34052_);
  nand (_11243_, _10915_, _34017_);
  and (_11244_, _11243_, _11014_);
  and (_11245_, _11244_, _11242_);
  or (_39056_[4], _11245_, _11241_);
  and (_11246_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_11247_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_11248_, _11247_, _11246_);
  and (_11249_, _11248_, _11049_);
  or (_11250_, _10916_, _33978_);
  nand (_11251_, _10916_, _34017_);
  and (_11252_, _11251_, _11014_);
  and (_11253_, _11252_, _11250_);
  or (_39056_[5], _11253_, _11249_);
  and (_11254_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_11255_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or (_11256_, _11255_, _11254_);
  and (_11257_, _11256_, _11049_);
  or (_11258_, _10915_, _33978_);
  or (_11259_, _10916_, _33942_);
  and (_11260_, _11259_, _11014_);
  and (_11261_, _11260_, _11258_);
  or (_39056_[6], _11261_, _11257_);
  and (_11262_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_11263_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_11264_, _11263_, _11262_);
  and (_11265_, _11264_, _11049_);
  nand (_11266_, _10915_, _34221_);
  or (_11267_, _10915_, _33942_);
  and (_11268_, _11267_, _11014_);
  and (_11269_, _11268_, _11266_);
  or (_39056_[7], _11269_, _11265_);
  or (_11270_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or (_11271_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and (_11272_, _11271_, _38997_);
  and (_11273_, _11272_, _11270_);
  or (_11274_, _11273_, _11014_);
  and (_11275_, _11013_, _10916_);
  nand (_11276_, _11275_, _34221_);
  and (_39056_[8], _11276_, _11274_);
  and (_11277_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_11278_, _11069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_11279_, _11278_, _11277_);
  and (_11280_, _11279_, _11049_);
  not (_11281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_11282_, _11281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_11283_, _11282_, _10916_);
  and (_11284_, _11283_, _11014_);
  or (_39056_[9], _11284_, _11280_);
  nand (_11285_, _11077_, _34148_);
  or (_11286_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_11287_, _11286_, _38997_);
  and (_39057_[0], _11287_, _11285_);
  not (_11288_, _11077_);
  or (_11289_, _11288_, _34122_);
  or (_11290_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_11291_, _11290_, _38997_);
  and (_39057_[1], _11291_, _11289_);
  or (_11292_, _11288_, _34089_);
  or (_11293_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_11294_, _11293_, _38997_);
  and (_39057_[2], _11294_, _11292_);
  nand (_11295_, _11077_, _34052_);
  or (_11296_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_11297_, _11296_, _38997_);
  and (_39057_[3], _11297_, _11295_);
  nand (_11298_, _11077_, _34017_);
  or (_11299_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_11300_, _11299_, _38997_);
  and (_39057_[4], _11300_, _11298_);
  or (_11301_, _11288_, _33978_);
  or (_11302_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_11303_, _11302_, _38997_);
  and (_39057_[5], _11303_, _11301_);
  or (_11304_, _11288_, _33942_);
  or (_11305_, _11077_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_11306_, _11305_, _38997_);
  and (_39057_[6], _11306_, _11304_);
  not (_11307_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_11308_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _11307_);
  or (_11309_, _11308_, _10915_);
  nor (_11310_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_11311_, _11310_, _11309_);
  or (_11312_, _11311_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_11313_, _11312_, _11086_);
  not (_11314_, _34229_);
  nor (_11315_, _35722_, _11314_);
  nand (_11316_, _11314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_11317_, _11316_, _11086_);
  or (_11318_, _11317_, _11315_);
  and (_11319_, _11318_, _11313_);
  or (_11320_, _11319_, _11092_);
  nand (_11321_, _11092_, _34148_);
  and (_11322_, _11321_, _38997_);
  and (_39058_[0], _11322_, _11320_);
  or (_11323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_11324_, _11323_, _11086_);
  not (_11325_, _34253_);
  nor (_11326_, _35722_, _11325_);
  nand (_11327_, _11325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_11328_, _11327_, _11086_);
  or (_11329_, _11328_, _11326_);
  and (_11330_, _11329_, _11324_);
  or (_11331_, _11330_, _11092_);
  or (_11332_, _11093_, _34122_);
  and (_11333_, _11332_, _38997_);
  and (_39058_[1], _11333_, _11331_);
  not (_11334_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not (_11335_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_11336_, _10928_, _11335_);
  nor (_11337_, _11336_, _11334_);
  and (_11338_, _11336_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_11339_, _11338_, _11337_);
  or (_11340_, _11339_, _11086_);
  not (_11341_, _33571_);
  and (_11342_, _11341_, _33558_);
  and (_11343_, _11342_, _33644_);
  not (_11344_, _11343_);
  nor (_11345_, _11344_, _35722_);
  or (_11346_, _11343_, _11334_);
  nand (_11347_, _11346_, _11086_);
  or (_11348_, _11347_, _11345_);
  and (_11349_, _11348_, _11340_);
  or (_11350_, _11349_, _11092_);
  or (_11351_, _11093_, _34089_);
  and (_11352_, _11351_, _38997_);
  and (_39058_[2], _11352_, _11350_);
  nand (_11353_, _11086_, _33644_);
  and (_11354_, _11353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_11355_, _11354_, _11092_);
  and (_11356_, _11074_, _33644_);
  and (_11357_, _11356_, _35723_);
  or (_11358_, _11074_, _11073_);
  not (_11359_, _11358_);
  and (_11360_, _11359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_11361_, _11360_, _11357_);
  and (_11362_, _11361_, _11086_);
  or (_11363_, _11362_, _11355_);
  nand (_11364_, _11092_, _34052_);
  and (_11365_, _11364_, _38997_);
  and (_39058_[3], _11365_, _11363_);
  and (_11366_, _11083_, _34251_);
  and (_11367_, _11366_, _34227_);
  and (_11368_, _11367_, _34706_);
  nand (_11369_, _11368_, _11081_);
  and (_11370_, _34228_, _11073_);
  nor (_11371_, _34228_, _11073_);
  nor (_11372_, _11371_, _11370_);
  or (_11373_, _11372_, _11369_);
  and (_11374_, _11373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_11375_, _11374_, _11092_);
  and (_11376_, _11370_, _35723_);
  and (_11377_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_11378_, _11377_, _11376_);
  and (_11379_, _11378_, _11086_);
  or (_11380_, _11379_, _11375_);
  nand (_11381_, _11092_, _34017_);
  and (_11382_, _11381_, _38997_);
  and (_39058_[4], _11382_, _11380_);
  and (_11383_, _11073_, _33572_);
  and (_11384_, _11086_, _11383_);
  or (_11385_, _11384_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_11386_, _11385_, _11093_);
  nand (_11387_, _11384_, _35722_);
  and (_11388_, _11387_, _11386_);
  and (_11389_, _11092_, _33978_);
  or (_11390_, _11389_, _11388_);
  and (_39058_[5], _11390_, _38997_);
  nor (_11391_, _33644_, _33571_);
  and (_11392_, _11391_, _33558_);
  not (_11393_, _11392_);
  or (_11394_, _11369_, _11393_);
  and (_11395_, _11394_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_11396_, _11395_, _11092_);
  nor (_11397_, _11394_, _35722_);
  or (_11398_, _11397_, _11396_);
  or (_11399_, _11093_, _33942_);
  and (_11400_, _11399_, _38997_);
  and (_39058_[6], _11400_, _11398_);
  and (_39019_, t0_i, _38997_);
  and (_39020_, t1_i, _38997_);
  and (_11401_, _11090_, _11356_);
  and (_11402_, _11401_, _33633_);
  nand (_11403_, _11402_, _34221_);
  not (_11404_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_11405_, _11404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  not (_11406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_11407_, _11406_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_11408_, t1_i);
  and (_11409_, _11408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_11410_, _11409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_11411_, _11410_, _11407_);
  and (_11412_, _11411_, _11405_);
  and (_11413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_11414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_11415_, _11414_, _11413_);
  and (_11416_, _11415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_11417_, _11416_, _11412_);
  and (_11418_, _11417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_11419_, _11418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  not (_11420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_11421_, _11420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_11422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_11423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _11422_);
  nor (_11424_, _11423_, _11421_);
  and (_11425_, _11090_, _11383_);
  and (_11426_, _11425_, _33633_);
  nor (_11427_, _11426_, _11424_);
  and (_11428_, _11427_, _11419_);
  or (_11429_, _11428_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_11430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_11431_, _11430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_11432_, _11431_, _11417_);
  nand (_11433_, _11432_, _11427_);
  and (_11434_, _11433_, _11429_);
  and (_11435_, _11419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_11436_, _11435_, _11421_);
  nand (_11437_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_11438_, _11437_, _11426_);
  or (_11439_, _11438_, _11434_);
  or (_11440_, _11439_, _11402_);
  and (_11441_, _11440_, _38997_);
  and (_39021_[7], _11441_, _11403_);
  not (_11442_, _11402_);
  and (_11443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_11444_, _11443_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_11445_, _11444_, _11417_);
  and (_11446_, _11445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_11447_, _11446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_11448_, _11447_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_11449_, _11448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_11450_, _11449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_11451_, _11450_, _11431_);
  not (_11452_, _11423_);
  nor (_11453_, _11431_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_11454_, _11453_, _11452_);
  nor (_11455_, _11454_, _11451_);
  and (_11456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_11457_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_11458_, _11450_);
  and (_11459_, _11458_, _11457_);
  or (_11460_, _11459_, _11456_);
  or (_11461_, _11460_, _11455_);
  nor (_11462_, _11449_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_11463_, _11462_, _11426_);
  and (_11464_, _11463_, _11461_);
  not (_11465_, _11426_);
  nor (_11466_, _11465_, _34221_);
  or (_11467_, _11466_, _11464_);
  and (_11468_, _11467_, _11442_);
  and (_11469_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_11470_, _11469_, _11468_);
  and (_39022_[7], _11470_, _38997_);
  not (_11471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_11472_, _11412_, _11471_);
  or (_11473_, _11472_, _11451_);
  and (_11474_, _11473_, _11423_);
  or (_11475_, _11472_, _11450_);
  and (_11476_, _11475_, _11457_);
  and (_11477_, _11432_, _11421_);
  nand (_11478_, _11412_, _11420_);
  and (_11479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_11480_, _11479_, _11478_);
  or (_11481_, _11480_, _11477_);
  or (_11482_, _11481_, _11476_);
  or (_11483_, _11482_, _11474_);
  nor (_11484_, _11402_, rst);
  and (_11485_, _11484_, _11465_);
  and (_39023_, _11485_, _11483_);
  and (_11486_, _11090_, _11370_);
  and (_11487_, _11486_, _33633_);
  nor (_11488_, _11487_, rst);
  not (_11489_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_11490_, t0_i);
  and (_11491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _11490_);
  nor (_11492_, _11491_, _11489_);
  not (_11493_, _11492_);
  not (_11494_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_11495_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_11496_, _11495_, _11494_);
  and (_11497_, _11496_, _11493_);
  not (_11498_, _11497_);
  and (_11499_, _11498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_11500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_11501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_11502_, _11501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_11503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_11504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_11505_, _11504_, _11503_);
  and (_11506_, _11505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_11507_, _11506_, _11497_);
  and (_11508_, _11507_, _11502_);
  and (_11509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_11510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_11511_, _11510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11512_, _11511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_11513_, _11512_, _11509_);
  and (_11514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_11515_, _11514_, _11513_);
  or (_11516_, _11515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_11517_, _11516_, _11508_);
  nor (_11518_, _11517_, _11500_);
  and (_11519_, _11513_, _11507_);
  nand (_11520_, _11519_, _11514_);
  and (_11521_, _11520_, _11500_);
  nor (_11522_, _11521_, _11518_);
  nor (_11523_, _11522_, _11499_);
  and (_11524_, _11090_, _11343_);
  and (_11525_, _11524_, _33633_);
  nor (_11526_, _11525_, _11523_);
  and (_39024_, _11526_, _11488_);
  and (_11527_, _11500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_11528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_11529_, _11528_, _11507_);
  or (_11530_, _11529_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_11531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _11531_);
  and (_11533_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_11534_, _11508_, _11500_);
  or (_11535_, _11534_, _11533_);
  or (_11536_, _11535_, _11487_);
  and (_11537_, _11536_, _11530_);
  or (_11538_, _11537_, _11527_);
  not (_11539_, _11525_);
  not (_11540_, _11487_);
  or (_11541_, _11540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_11542_, _11541_, _11539_);
  and (_11543_, _11542_, _11538_);
  nor (_11544_, _11539_, _34221_);
  or (_11545_, _11544_, _11543_);
  and (_39025_[7], _11545_, _38997_);
  nand (_11546_, _11487_, _34221_);
  and (_11547_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _11531_);
  or (_11548_, _11532_, _11547_);
  not (_11549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_11550_, _11506_, _11502_);
  and (_11551_, _11497_, _11531_);
  and (_11552_, _11551_, _11550_);
  and (_11553_, _11552_, _11513_);
  and (_11554_, _11553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_11555_, _11554_, _11549_);
  and (_11556_, _11554_, _11549_);
  or (_11557_, _11556_, _11555_);
  and (_11558_, _11557_, _11548_);
  and (_11559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_11560_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_11561_, _11560_, _11512_);
  and (_11562_, _11561_, _11509_);
  and (_11563_, _11562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_11564_, _11563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_11565_, _11560_, _11515_);
  and (_11566_, _11565_, _11564_);
  and (_11567_, _11566_, _11559_);
  and (_11568_, _11519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_11569_, _11568_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_11570_, _11569_, _11521_);
  or (_11571_, _11570_, _11567_);
  or (_11572_, _11571_, _11558_);
  or (_11573_, _11572_, _11487_);
  and (_11574_, _11573_, _11539_);
  and (_11575_, _11574_, _11546_);
  and (_11576_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_11577_, _11576_, _11575_);
  and (_39026_[7], _11577_, _38997_);
  or (_11578_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_11579_, _11559_, _38997_);
  and (_11580_, _11579_, _11578_);
  not (_11581_, _11560_);
  or (_11582_, _11581_, _11515_);
  nand (_11583_, _11582_, _11580_);
  nor (_11584_, _11583_, _11487_);
  and (_39027_, _11584_, _11539_);
  and (_11585_, _34254_, _33633_);
  and (_11586_, _11585_, _33662_);
  or (_11587_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_11588_, _11587_, _38997_);
  nand (_11589_, _11586_, _34221_);
  and (_39028_[7], _11589_, _11588_);
  and (_11590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_11591_, _11590_, _11426_);
  not (_11592_, _11591_);
  and (_11593_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_11594_, _11431_, _11416_);
  and (_11595_, _11594_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_11596_, _11595_, _11421_);
  not (_11597_, _11590_);
  and (_11598_, _11412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_11599_, _11412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_11600_, _11599_, _11598_);
  and (_11601_, _11600_, _11597_);
  nor (_11602_, _11601_, _11596_);
  nor (_11603_, _11602_, _11426_);
  or (_11604_, _11603_, _11402_);
  or (_11605_, _11604_, _11593_);
  nand (_11606_, _11402_, _34148_);
  and (_11607_, _11606_, _38997_);
  and (_39021_[0], _11607_, _11605_);
  or (_11608_, _11442_, _34122_);
  and (_11609_, _11598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_11610_, _11598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_11611_, _11610_, _11609_);
  and (_11612_, _11611_, _11591_);
  and (_11613_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_11614_, _11477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_11615_, _11614_, _11426_);
  or (_11616_, _11615_, _11613_);
  or (_11617_, _11616_, _11612_);
  or (_11618_, _11617_, _11402_);
  and (_11619_, _11618_, _38997_);
  and (_39021_[1], _11619_, _11608_);
  or (_11620_, _11442_, _34089_);
  and (_11621_, _11598_, _11413_);
  nor (_11622_, _11609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_11623_, _11622_, _11621_);
  and (_11624_, _11623_, _11591_);
  and (_11625_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand (_11626_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_11627_, _11626_, _11426_);
  or (_11628_, _11627_, _11625_);
  or (_11629_, _11628_, _11624_);
  or (_11630_, _11629_, _11402_);
  and (_11631_, _11630_, _38997_);
  and (_39021_[2], _11631_, _11620_);
  nand (_11632_, _11402_, _34052_);
  and (_11633_, _11415_, _11412_);
  nor (_11634_, _11621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_11635_, _11634_, _11633_);
  and (_11636_, _11635_, _11591_);
  and (_11637_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_11638_, _11477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_11639_, _11638_, _11426_);
  or (_11640_, _11639_, _11637_);
  or (_11641_, _11640_, _11636_);
  or (_11642_, _11641_, _11402_);
  and (_11643_, _11642_, _38997_);
  and (_39021_[3], _11643_, _11632_);
  nand (_11644_, _11402_, _34017_);
  and (_11645_, _11592_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_11646_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_11647_, _11633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_11648_, _11647_, _11417_);
  and (_11649_, _11648_, _11597_);
  nor (_11650_, _11649_, _11646_);
  nor (_11651_, _11650_, _11426_);
  or (_11652_, _11651_, _11645_);
  or (_11653_, _11652_, _11402_);
  and (_11654_, _11653_, _38997_);
  and (_39021_[4], _11654_, _11644_);
  or (_11655_, _11442_, _33978_);
  not (_11656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_11657_, _11427_, _11656_);
  and (_11658_, _11436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_11659_, _11424_);
  nor (_11660_, _11417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_11661_, _11660_, _11418_);
  and (_11662_, _11661_, _11659_);
  nor (_11663_, _11662_, _11658_);
  nor (_11664_, _11663_, _11426_);
  or (_11665_, _11664_, _11657_);
  or (_11666_, _11665_, _11402_);
  and (_11667_, _11666_, _38997_);
  and (_39021_[5], _11667_, _11655_);
  or (_11668_, _11442_, _33942_);
  not (_11669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_11670_, _11427_, _11669_);
  and (_11671_, _11421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_11672_, _11671_, _11412_);
  and (_11673_, _11672_, _11594_);
  or (_11674_, _11418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_11675_, _11674_, _11659_);
  nor (_11676_, _11675_, _11419_);
  nor (_11677_, _11676_, _11673_);
  nor (_11678_, _11677_, _11426_);
  or (_11679_, _11678_, _11670_);
  or (_11680_, _11679_, _11402_);
  and (_11681_, _11680_, _38997_);
  and (_39021_[6], _11681_, _11668_);
  not (_11682_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_11683_, _11417_, _11422_);
  nor (_11684_, _11431_, _11420_);
  not (_11685_, _11684_);
  and (_11686_, _11685_, _11683_);
  and (_11687_, _11686_, _11682_);
  nor (_11688_, _11686_, _11682_);
  or (_11689_, _11688_, _11687_);
  or (_11690_, _11689_, _11426_);
  nand (_11691_, _11426_, _34148_);
  and (_11692_, _11691_, _11690_);
  or (_11693_, _11692_, _11402_);
  nand (_11694_, _11402_, _11682_);
  and (_11695_, _11694_, _38997_);
  and (_39022_[0], _11695_, _11693_);
  or (_11696_, _11465_, _34122_);
  not (_11697_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_11698_, _11432_, _11452_);
  not (_11699_, _11698_);
  nor (_11700_, _11683_, _11423_);
  nor (_11701_, _11700_, _11682_);
  and (_11702_, _11701_, _11699_);
  nor (_11703_, _11702_, _11697_);
  and (_11704_, _11702_, _11697_);
  or (_11705_, _11704_, _11703_);
  or (_11706_, _11705_, _11426_);
  and (_11707_, _11706_, _11442_);
  and (_11708_, _11707_, _11696_);
  and (_11709_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_11710_, _11709_, _11708_);
  and (_39022_[1], _11710_, _38997_);
  or (_11711_, _11465_, _34089_);
  and (_11712_, _11445_, _11422_);
  and (_11713_, _11685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_11714_, _11713_, _11712_);
  or (_11715_, _11684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_11716_, _11715_);
  and (_11717_, _11443_, _11417_);
  and (_11718_, _11717_, _11716_);
  or (_11719_, _11718_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_11720_, _11719_, _11714_);
  or (_11721_, _11720_, _11426_);
  and (_11722_, _11721_, _11442_);
  and (_11723_, _11722_, _11711_);
  and (_11724_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_11725_, _11724_, _11723_);
  and (_39022_[2], _11725_, _38997_);
  nand (_11726_, _11426_, _34052_);
  or (_11727_, _11712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_11728_, _11712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_11729_, _11728_, _11727_);
  or (_11730_, _11729_, _11423_);
  and (_11731_, _11443_, _11594_);
  and (_11732_, _11731_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_11733_, _11732_, _11412_);
  nor (_11734_, _11733_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_11735_, _11733_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_11736_, _11735_, _11734_);
  or (_11737_, _11736_, _11452_);
  and (_11738_, _11737_, _11730_);
  or (_11739_, _11738_, _11426_);
  and (_11740_, _11739_, _11442_);
  and (_11741_, _11740_, _11726_);
  and (_11742_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_11743_, _11742_, _11741_);
  and (_39022_[3], _11743_, _38997_);
  nand (_11744_, _11426_, _34017_);
  or (_11745_, _11735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_11746_, _11447_, _11431_);
  and (_11747_, _11746_, _11423_);
  and (_11748_, _11747_, _11745_);
  and (_11749_, _11443_, _11416_);
  and (_11750_, _11749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_11751_, _11750_, _11412_);
  and (_11752_, _11751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_11753_, _11752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_11754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not (_11755_, _11447_);
  and (_11756_, _11755_, _11457_);
  or (_11757_, _11756_, _11754_);
  and (_11758_, _11757_, _11753_);
  or (_11759_, _11758_, _11748_);
  or (_11760_, _11759_, _11426_);
  and (_11761_, _11760_, _11442_);
  and (_11762_, _11761_, _11744_);
  and (_11763_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_11764_, _11763_, _11762_);
  and (_39022_[4], _11764_, _38997_);
  or (_11765_, _11465_, _33978_);
  not (_11766_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_11767_, _11716_, _11447_);
  nor (_11768_, _11767_, _11766_);
  and (_11769_, _11767_, _11766_);
  or (_11770_, _11769_, _11768_);
  or (_11771_, _11770_, _11426_);
  and (_11772_, _11771_, _11442_);
  and (_11773_, _11772_, _11765_);
  and (_11774_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_11775_, _11774_, _11773_);
  and (_39022_[5], _11775_, _38997_);
  or (_11776_, _11465_, _33942_);
  not (_11777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_11778_, _11716_, _11448_);
  nor (_11779_, _11778_, _11777_);
  and (_11780_, _11778_, _11777_);
  or (_11781_, _11780_, _11779_);
  or (_11782_, _11781_, _11426_);
  and (_11783_, _11782_, _11442_);
  and (_11784_, _11783_, _11776_);
  and (_11785_, _11402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_11786_, _11785_, _11784_);
  and (_39022_[6], _11786_, _38997_);
  nor (_11787_, _11498_, _11487_);
  or (_11788_, _11787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_11789_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_11790_, _11789_, _11550_);
  and (_11791_, _11497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_11792_, _11791_, _11790_);
  or (_11793_, _11792_, _11487_);
  and (_11794_, _11793_, _11788_);
  or (_11795_, _11794_, _11525_);
  nand (_11796_, _11525_, _34148_);
  and (_11797_, _11796_, _38997_);
  and (_39025_[0], _11797_, _11795_);
  or (_11798_, _11539_, _34122_);
  and (_11799_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_11800_, _11799_, _11525_);
  and (_11801_, _11800_, _38997_);
  nor (_11802_, _11791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_11803_, _11791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_11804_, _11803_, _11802_);
  and (_11805_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_11806_, _11805_, _11508_);
  or (_11807_, _11806_, _11804_);
  and (_11808_, _11807_, _11488_);
  or (_11809_, _11808_, _11801_);
  and (_39025_[1], _11809_, _11798_);
  or (_11810_, _11539_, _34089_);
  nor (_11811_, _11803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_11812_, _11791_, _11503_);
  nor (_11813_, _11812_, _11811_);
  and (_11814_, _11532_, _11508_);
  and (_11815_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_11816_, _11815_, _11813_);
  nor (_11817_, _11816_, _11487_);
  and (_11818_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_11819_, _11818_, _11817_);
  or (_11820_, _11819_, _11525_);
  and (_11821_, _11820_, _38997_);
  and (_39025_[2], _11821_, _11810_);
  and (_11822_, _11505_, _11497_);
  nor (_11823_, _11812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_11824_, _11823_, _11822_);
  and (_11825_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_11826_, _11825_, _11824_);
  nor (_11827_, _11826_, _11487_);
  and (_11828_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_11829_, _11828_, _11827_);
  and (_11830_, _11829_, _11539_);
  nor (_11831_, _11539_, _34052_);
  or (_11832_, _11831_, _11830_);
  and (_39025_[3], _11832_, _38997_);
  nor (_11833_, _11822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_11834_, _11833_, _11507_);
  and (_11835_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_11836_, _11835_, _11834_);
  nor (_11837_, _11836_, _11487_);
  and (_11838_, _11487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_11839_, _11838_, _11837_);
  and (_11840_, _11839_, _11539_);
  nor (_11841_, _11539_, _34017_);
  or (_11842_, _11841_, _11840_);
  and (_39025_[4], _11842_, _38997_);
  or (_11843_, _11539_, _33978_);
  nand (_11844_, _11814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_11845_, _11500_);
  nand (_11846_, _11507_, _11845_);
  or (_11847_, _11846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_11848_, _11847_, _11844_);
  nor (_11849_, _11848_, _11487_);
  not (_11850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_11851_, _11846_, _11850_);
  or (_11852_, _11851_, _11487_);
  and (_11853_, _11852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_11854_, _11853_, _11849_);
  or (_11855_, _11854_, _11525_);
  and (_11856_, _11855_, _38997_);
  and (_39025_[5], _11856_, _11843_);
  and (_11857_, _11852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_11858_, _11532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_11859_, _11858_, _11497_);
  and (_11860_, _11859_, _11550_);
  nor (_11861_, _11851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_11862_, _11861_, _11860_);
  nor (_11863_, _11862_, _11487_);
  or (_11864_, _11863_, _11857_);
  and (_11865_, _11864_, _11539_);
  and (_11866_, _11525_, _33942_);
  or (_11867_, _11866_, _11865_);
  and (_39025_[6], _11867_, _38997_);
  or (_11868_, _11552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_11869_, _11552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not (_11870_, _11869_);
  and (_11871_, _11870_, _11548_);
  and (_11872_, _11871_, _11868_);
  and (_11873_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_11874_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_11875_, _11874_, _11559_);
  nor (_11876_, _11875_, _11873_);
  and (_11877_, _11507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_11878_, _11507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_11879_, _11878_, _11500_);
  nor (_11880_, _11879_, _11877_);
  or (_11881_, _11880_, _11876_);
  nor (_11882_, _11881_, _11872_);
  nand (_11883_, _11882_, _11540_);
  nand (_11884_, _11487_, _34148_);
  and (_11885_, _11884_, _11539_);
  and (_11886_, _11885_, _11883_);
  and (_11887_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_11888_, _11887_, _11886_);
  and (_39026_[0], _11888_, _38997_);
  or (_11889_, _11540_, _34122_);
  or (_11890_, _11869_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_11891_, _11550_, _11497_);
  and (_11892_, _11891_, _11510_);
  not (_11893_, _11892_);
  or (_11894_, _11893_, _11532_);
  and (_11895_, _11894_, _11548_);
  and (_11896_, _11895_, _11890_);
  and (_11897_, _11560_, _11510_);
  or (_11898_, _11873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_11899_, _11898_, _11559_);
  nor (_11900_, _11899_, _11897_);
  and (_11901_, _11877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_11902_, _11877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_11903_, _11902_, _11500_);
  nor (_11904_, _11903_, _11901_);
  or (_11905_, _11904_, _11900_);
  or (_11906_, _11905_, _11896_);
  or (_11907_, _11906_, _11487_);
  and (_11908_, _11907_, _11539_);
  and (_11909_, _11908_, _11889_);
  and (_11910_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_11911_, _11910_, _11909_);
  and (_39026_[1], _11911_, _38997_);
  or (_11912_, _11540_, _34089_);
  or (_11913_, _11892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11914_, _11891_, _11511_);
  not (_11915_, _11914_);
  and (_11916_, _11915_, _11547_);
  and (_11917_, _11916_, _11913_);
  and (_11918_, _11510_, _11497_);
  and (_11919_, _11918_, _11506_);
  or (_11920_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11921_, _11511_, _11507_);
  nor (_11922_, _11921_, _11845_);
  and (_11923_, _11922_, _11920_);
  and (_11924_, _11897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_11925_, _11924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11926_, _11560_, _11511_);
  nand (_11927_, _11926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_11928_, _11927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_11929_, _11928_, _11925_);
  or (_11930_, _11929_, _11923_);
  or (_11931_, _11930_, _11917_);
  or (_11932_, _11931_, _11487_);
  and (_11933_, _11932_, _11539_);
  and (_11934_, _11933_, _11912_);
  and (_11935_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_11936_, _11935_, _11934_);
  and (_39026_[2], _11936_, _38997_);
  nand (_11937_, _11487_, _34052_);
  not (_11938_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_11939_, _11914_, _11531_);
  nor (_11940_, _11939_, _11938_);
  and (_11941_, _11939_, _11938_);
  or (_11942_, _11941_, _11940_);
  and (_11943_, _11942_, _11548_);
  or (_11944_, _11926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_11945_, _11561_);
  and (_11946_, _11945_, _11559_);
  and (_11947_, _11946_, _11944_);
  or (_11948_, _11921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_11949_, _11512_, _11507_);
  nor (_11950_, _11949_, _11845_);
  and (_11951_, _11950_, _11948_);
  or (_11952_, _11951_, _11947_);
  or (_11953_, _11952_, _11943_);
  or (_11954_, _11953_, _11487_);
  and (_11955_, _11954_, _11539_);
  and (_11956_, _11955_, _11937_);
  and (_11957_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_11958_, _11957_, _11956_);
  and (_39026_[3], _11958_, _38997_);
  nand (_11959_, _11487_, _34017_);
  or (_11960_, _11949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_11961_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11962_, _11961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_11963_, _11962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_11964_, _11963_, _11845_);
  and (_11965_, _11964_, _11960_);
  and (_11966_, _11512_, _11497_);
  and (_11967_, _11966_, _11550_);
  or (_11968_, _11967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_11969_, _11967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_11970_, _11969_);
  and (_11971_, _11970_, _11547_);
  and (_11972_, _11971_, _11968_);
  and (_11973_, _11561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_11974_, _11973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_11975_, _11561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_11976_, _11975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_11977_, _11976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_11978_, _11977_, _11974_);
  or (_11979_, _11978_, _11972_);
  or (_11980_, _11979_, _11965_);
  or (_11981_, _11980_, _11487_);
  and (_11982_, _11981_, _11539_);
  and (_11983_, _11982_, _11959_);
  and (_11984_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_11985_, _11984_, _11983_);
  and (_39026_[4], _11985_, _38997_);
  or (_11986_, _11540_, _33978_);
  not (_11987_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_11988_, _11963_, _11987_);
  nor (_11989_, _11963_, _11987_);
  or (_11990_, _11989_, _11988_);
  and (_11991_, _11990_, _11500_);
  not (_11992_, _11562_);
  and (_11993_, _11992_, _11559_);
  or (_11994_, _11973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_11995_, _11994_, _11993_);
  and (_11996_, _11969_, _11531_);
  nand (_11997_, _11996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_11998_, _11996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_11999_, _11998_, _11997_);
  and (_12000_, _11999_, _11548_);
  or (_12001_, _12000_, _11995_);
  or (_12002_, _12001_, _11991_);
  or (_12003_, _12002_, _11487_);
  and (_12004_, _12003_, _11539_);
  and (_12005_, _12004_, _11986_);
  and (_12006_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_12007_, _12006_, _12005_);
  and (_39026_[5], _12007_, _38997_);
  or (_12008_, _11540_, _33942_);
  or (_12009_, _11553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_12010_, _12009_, _11548_);
  nor (_12011_, _12010_, _11554_);
  or (_12012_, _11562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_12013_, _11563_);
  and (_12014_, _12013_, _11559_);
  and (_12015_, _12014_, _12012_);
  or (_12016_, _11519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_12017_, _11568_, _11845_);
  and (_12018_, _12017_, _12016_);
  or (_12019_, _12018_, _12015_);
  or (_12020_, _12019_, _12011_);
  or (_12021_, _12020_, _11487_);
  and (_12022_, _12021_, _11539_);
  and (_12023_, _12022_, _12008_);
  and (_12024_, _11525_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_12025_, _12024_, _12023_);
  and (_39026_[6], _12025_, _38997_);
  nand (_12026_, _11586_, _34148_);
  or (_12027_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_12028_, _12027_, _38997_);
  and (_39028_[0], _12028_, _12026_);
  or (_12029_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_12030_, _12029_, _38997_);
  not (_12031_, _11586_);
  or (_12032_, _12031_, _34122_);
  and (_39028_[1], _12032_, _12030_);
  or (_12033_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_12034_, _12033_, _38997_);
  or (_12035_, _12031_, _34089_);
  and (_39028_[2], _12035_, _12034_);
  or (_12036_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_12037_, _12036_, _38997_);
  nand (_12038_, _11586_, _34052_);
  and (_39028_[3], _12038_, _12037_);
  or (_12039_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_12040_, _12039_, _38997_);
  nand (_12041_, _11586_, _34017_);
  and (_39028_[4], _12041_, _12040_);
  or (_12042_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_12043_, _12042_, _38997_);
  or (_12044_, _12031_, _33978_);
  and (_39028_[5], _12044_, _12043_);
  or (_12045_, _11586_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_12046_, _12045_, _38997_);
  or (_12047_, _12031_, _33942_);
  and (_39028_[6], _12047_, _12046_);
  and (_12048_, _33630_, _34232_);
  and (_12049_, _12048_, _11085_);
  and (_12050_, _12049_, _11075_);
  or (_12051_, _12050_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor (_12052_, _33604_, _33591_);
  and (_12053_, _12052_, _33632_);
  and (_12054_, _12053_, _11076_);
  not (_12055_, _12054_);
  and (_12056_, _12055_, _12051_);
  nand (_12057_, _12050_, _35722_);
  and (_12058_, _12057_, _12056_);
  nor (_12059_, _12055_, _34221_);
  or (_12060_, _12059_, _12058_);
  and (_39011_[7], _12060_, _38997_);
  and (_12061_, _34251_, _33604_);
  and (_12062_, _12061_, _11084_);
  and (_12063_, _12062_, _12048_);
  and (_12064_, _12063_, _11075_);
  or (_12065_, _12064_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_12066_, _33604_, _34232_);
  and (_12067_, _12066_, _33632_);
  and (_12068_, _12067_, _11091_);
  not (_12069_, _12068_);
  and (_12070_, _12069_, _12065_);
  nand (_12071_, _12064_, _35722_);
  and (_12072_, _12071_, _12070_);
  nor (_12073_, _12069_, _34221_);
  or (_12074_, _12073_, _12072_);
  and (_39010_[7], _12074_, _38997_);
  and (_12075_, _12062_, _11081_);
  nand (_12076_, _12075_, _33558_);
  and (_12077_, _12076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_12078_, _11091_, _33633_);
  or (_12079_, _12078_, _12077_);
  nor (_12080_, _11393_, _35722_);
  nand (_12081_, _33558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_12082_, _12081_, _11391_);
  or (_12083_, _12082_, _12080_);
  and (_12084_, _12083_, _12075_);
  or (_12085_, _12084_, _12079_);
  not (_12086_, _12078_);
  or (_12087_, _12086_, _33942_);
  and (_12088_, _12087_, _38997_);
  and (_39009_[3], _12088_, _12085_);
  nor (_12089_, _10898_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not (_12090_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_12091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_12093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _12092_);
  and (_12094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_12095_, _12094_, _12093_);
  nor (_12096_, _12095_, _12091_);
  or (_12097_, _12096_, _12090_);
  and (_12098_, _12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_12099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_12100_, _12099_, _12098_);
  nor (_12101_, _12100_, _12091_);
  and (_12102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _12092_);
  and (_12103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_12104_, _12103_, _12102_);
  nand (_12105_, _12104_, _12101_);
  or (_12106_, _12105_, _12097_);
  and (_12107_, _12106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_12108_, _12107_, _12089_);
  and (_12109_, _11366_, _33633_);
  and (_12110_, _12109_, _11075_);
  or (_12111_, _12110_, _12108_);
  and (_12112_, _12111_, _12086_);
  nand (_12113_, _12110_, _35722_);
  and (_12114_, _12113_, _12112_);
  nor (_12115_, _12086_, _34221_);
  or (_12116_, _12115_, _12114_);
  and (_39008_, _12116_, _38997_);
  not (_12117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and (_12118_, _12117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_12119_, _12104_, _12091_);
  not (_12120_, _12119_);
  or (_12121_, _12120_, _12101_);
  or (_12122_, _12121_, _12097_);
  and (_12123_, _12122_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_12124_, _12123_, _12118_);
  and (_12125_, _12109_, _11383_);
  or (_12126_, _12125_, _12124_);
  and (_12127_, _12126_, _12086_);
  nand (_12128_, _12125_, _35722_);
  and (_12129_, _12128_, _12127_);
  and (_12130_, _12078_, _33978_);
  or (_12131_, _12130_, _12129_);
  and (_39007_, _12131_, _38997_);
  not (_12132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_12133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _12132_);
  nand (_12134_, _12096_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_12135_, _12119_, _12101_);
  or (_12136_, _12135_, _12134_);
  and (_12137_, _12136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_12138_, _12137_, _12133_);
  and (_12139_, _11585_, _11083_);
  or (_12140_, _12139_, _12138_);
  and (_12141_, _12140_, _12086_);
  nand (_12142_, _12139_, _35722_);
  and (_12143_, _12142_, _12141_);
  and (_12144_, _12078_, _34122_);
  or (_12145_, _12144_, _12143_);
  and (_39006_, _12145_, _38997_);
  nand (_12146_, _12109_, _11356_);
  nor (_12147_, _12146_, _35722_);
  and (_12148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_12149_, _12134_, _12121_);
  and (_12150_, _12149_, _12148_);
  and (_12151_, _12150_, _12146_);
  or (_12152_, _12151_, _12078_);
  or (_12153_, _12152_, _12147_);
  nand (_12154_, _12078_, _34052_);
  and (_12155_, _12154_, _38997_);
  and (_39005_, _12155_, _12153_);
  nand (_12156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_12157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _12092_);
  and (_12158_, _12157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_12159_, _12158_, _12156_);
  or (_12160_, _12159_, _12091_);
  and (_12161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_12162_, _12161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_12163_, _12162_);
  and (_12164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_12165_, _12164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_12166_, _12165_);
  and (_12167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_12168_, _12167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_12169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_12170_, _12169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_12171_, _12170_, _12168_);
  and (_12172_, _12171_, _12166_);
  and (_12173_, _12172_, _12163_);
  not (_12174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_12175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_12176_, _12175_, _12174_);
  nand (_12177_, _12176_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_12178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_12179_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_12180_, _12179_, _12178_);
  and (_12181_, _12180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_12182_, _12181_);
  and (_12183_, _12182_, _12177_);
  nand (_12184_, _12183_, _12173_);
  and (_12185_, _12184_, _12160_);
  and (_12186_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_12187_, _12186_, _12092_);
  and (_12188_, _12187_, _12185_);
  not (_12189_, _12188_);
  not (_12190_, _12187_);
  and (_12191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _12091_);
  not (_12192_, _12191_);
  not (_12193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_12194_, _12164_, _12193_);
  not (_12195_, _12194_);
  not (_12196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_12197_, _12167_, _12196_);
  not (_12198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_12199_, _12169_, _12198_);
  nor (_12200_, _12199_, _12197_);
  and (_12201_, _12200_, _12195_);
  nor (_12202_, _12201_, _12192_);
  not (_12203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_12204_, _12176_, _12203_);
  not (_12205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_12206_, _12180_, _12205_);
  nor (_12207_, _12206_, _12204_);
  not (_12208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_12209_, _12161_, _12208_);
  not (_12210_, _12209_);
  and (_12211_, _12210_, _12207_);
  nor (_12212_, _12211_, _12192_);
  nor (_12213_, _12212_, _12202_);
  or (_12214_, _12213_, _12190_);
  and (_12215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _38997_);
  and (_12216_, _12215_, _12214_);
  and (_39004_[1], _12216_, _12189_);
  nor (_12217_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_12218_, _12217_);
  not (_12219_, _12185_);
  and (_12220_, _12213_, _12219_);
  nor (_12221_, _12220_, _12218_);
  nand (_12222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _38997_);
  nor (_39003_[1], _12222_, _12221_);
  and (_12223_, _12183_, _12163_);
  nand (_12224_, _12223_, _12185_);
  or (_12225_, _12212_, _12185_);
  and (_12226_, _12225_, _12187_);
  and (_12227_, _12226_, _12224_);
  or (_12228_, _12227_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_12229_, _12189_, _12172_);
  nor (_12230_, _12190_, _12185_);
  nand (_12231_, _12230_, _12202_);
  and (_12232_, _12231_, _38997_);
  and (_12233_, _12232_, _12229_);
  and (_39002_[2], _12233_, _12228_);
  and (_12234_, _12224_, _12217_);
  or (_12235_, _12234_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_12236_, _12217_, _12185_);
  not (_12237_, _12236_);
  or (_12238_, _12237_, _12172_);
  or (_12239_, _12212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand (_12240_, _12217_, _12202_);
  and (_12241_, _12240_, _12239_);
  or (_12242_, _12241_, _12185_);
  and (_12243_, _12242_, _38997_);
  and (_12244_, _12243_, _12238_);
  and (_39001_[2], _12244_, _12235_);
  nand (_12245_, _12220_, _12091_);
  nor (_12246_, _12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand (_12247_, _12246_, _12186_);
  and (_12248_, _12247_, _38997_);
  and (_39000_, _12248_, _12245_);
  and (_12249_, _12220_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_12250_, _12092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_12251_, _12250_, _12246_);
  nor (_12252_, _12251_, _12219_);
  or (_12253_, _12252_, _12186_);
  or (_12254_, _12253_, _12249_);
  not (_12255_, _12186_);
  or (_12256_, _12251_, _12255_);
  and (_12257_, _12256_, _38997_);
  and (_38999_[1], _12257_, _12254_);
  and (_12258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _38997_);
  and (_38998_[7], _12258_, _12186_);
  and (_38995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _38997_);
  nor (_12259_, _12220_, _12186_);
  and (_12260_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_12261_, _12260_, _12259_);
  and (_38998_[0], _12261_, _38997_);
  and (_12262_, _12186_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_12263_, _12262_, _12259_);
  and (_38998_[1], _12263_, _38997_);
  and (_12264_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _38997_);
  and (_38998_[2], _12264_, _12186_);
  not (_12265_, _12199_);
  nor (_12266_, _12206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_12267_, _12266_, _12204_);
  or (_12268_, _12267_, _12209_);
  and (_12269_, _12268_, _12265_);
  or (_12270_, _12269_, _12197_);
  nor (_12271_, _12213_, _12185_);
  and (_12272_, _12271_, _12195_);
  and (_12273_, _12272_, _12270_);
  not (_12274_, _12170_);
  or (_12275_, _12181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_12276_, _12275_, _12177_);
  or (_12277_, _12276_, _12162_);
  and (_12278_, _12277_, _12274_);
  or (_12279_, _12278_, _12168_);
  and (_12280_, _12185_, _12166_);
  and (_12281_, _12280_, _12279_);
  or (_12282_, _12281_, _12186_);
  or (_12283_, _12282_, _12273_);
  or (_12284_, _12255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_12285_, _12284_, _38997_);
  and (_38998_[3], _12285_, _12283_);
  not (_12286_, _12168_);
  or (_12287_, _12170_, _12162_);
  and (_12288_, _12183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_12289_, _12288_, _12287_);
  and (_12290_, _12289_, _12286_);
  and (_12291_, _12290_, _12280_);
  nor (_12292_, _12197_, _12194_);
  or (_12293_, _12209_, _12199_);
  and (_12294_, _12207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_12295_, _12294_, _12293_);
  and (_12296_, _12295_, _12292_);
  and (_12297_, _12296_, _12271_);
  or (_12298_, _12297_, _12186_);
  or (_12299_, _12298_, _12291_);
  or (_12300_, _12255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_12301_, _12300_, _38997_);
  and (_38998_[4], _12301_, _12299_);
  and (_12302_, _12210_, _12191_);
  nand (_12303_, _12302_, _12201_);
  or (_12304_, _12303_, _12207_);
  nor (_12305_, _12304_, _12185_);
  nand (_12306_, _12173_, _12160_);
  nor (_12307_, _12306_, _12183_);
  or (_12308_, _12307_, _12186_);
  or (_12309_, _12308_, _12305_);
  or (_12310_, _12255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_12311_, _12310_, _38997_);
  and (_38998_[5], _12311_, _12309_);
  and (_12312_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _38997_);
  and (_38998_[6], _12312_, _12186_);
  and (_12313_, _12186_, _12092_);
  or (_12314_, _12313_, _12221_);
  or (_12315_, _12314_, _12230_);
  and (_38999_[0], _12315_, _38997_);
  not (_12316_, _12259_);
  and (_12317_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_12318_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_12319_, _12181_, _12092_);
  or (_12320_, _12319_, _12318_);
  nor (_12321_, _12177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_12322_, _12321_, _12162_);
  nand (_12323_, _12322_, _12320_);
  or (_12324_, _12163_, _12094_);
  and (_12325_, _12324_, _12323_);
  or (_12326_, _12325_, _12170_);
  or (_12327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _12092_);
  or (_12328_, _12327_, _12274_);
  and (_12329_, _12328_, _12286_);
  and (_12330_, _12329_, _12326_);
  and (_12331_, _12168_, _12094_);
  or (_12332_, _12331_, _12165_);
  or (_12333_, _12332_, _12330_);
  or (_12334_, _12327_, _12166_);
  and (_12335_, _12334_, _12185_);
  and (_12336_, _12335_, _12333_);
  and (_12337_, _12206_, _12092_);
  or (_12338_, _12337_, _12318_);
  and (_12339_, _12204_, _12092_);
  nor (_12340_, _12339_, _12209_);
  nand (_12341_, _12340_, _12338_);
  or (_12342_, _12210_, _12094_);
  and (_12343_, _12342_, _12341_);
  or (_12344_, _12343_, _12199_);
  not (_12345_, _12197_);
  or (_12346_, _12327_, _12265_);
  and (_12347_, _12346_, _12345_);
  and (_12348_, _12347_, _12344_);
  and (_12349_, _12197_, _12094_);
  or (_12350_, _12349_, _12194_);
  or (_12351_, _12350_, _12348_);
  and (_12352_, _12327_, _12271_);
  or (_12353_, _12352_, _12272_);
  and (_12354_, _12353_, _12351_);
  or (_12355_, _12354_, _12336_);
  and (_12356_, _12355_, _12255_);
  or (_12357_, _12356_, _12317_);
  and (_39001_[0], _12357_, _38997_);
  and (_12358_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_12359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _12092_);
  and (_12360_, _12359_, _12166_);
  or (_12361_, _12360_, _12172_);
  or (_12362_, _12319_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_12363_, _12362_, _12322_);
  nand (_12364_, _12162_, _12103_);
  nand (_12365_, _12364_, _12171_);
  or (_12366_, _12365_, _12363_);
  and (_12367_, _12366_, _12361_);
  and (_12368_, _12165_, _12103_);
  or (_12369_, _12368_, _12367_);
  and (_12370_, _12369_, _12185_);
  and (_12371_, _12194_, _12103_);
  and (_12372_, _12359_, _12195_);
  or (_12373_, _12372_, _12201_);
  and (_12374_, _12209_, _12103_);
  not (_12375_, _12200_);
  or (_12376_, _12337_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_12377_, _12376_, _12340_);
  or (_12378_, _12377_, _12375_);
  or (_12379_, _12378_, _12374_);
  and (_12380_, _12379_, _12373_);
  or (_12381_, _12380_, _12371_);
  and (_12382_, _12381_, _12271_);
  or (_12383_, _12382_, _12370_);
  and (_12384_, _12383_, _12255_);
  or (_12385_, _12384_, _12358_);
  and (_39001_[1], _12385_, _38997_);
  and (_12386_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_12387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_12388_, _12181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_12389_, _12388_, _12387_);
  nor (_12390_, _12177_, _12092_);
  nor (_12391_, _12390_, _12162_);
  nand (_12392_, _12391_, _12389_);
  or (_12393_, _12163_, _12093_);
  and (_12394_, _12393_, _12392_);
  or (_12395_, _12394_, _12170_);
  or (_12396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_12397_, _12396_, _12274_);
  and (_12398_, _12397_, _12286_);
  and (_12399_, _12398_, _12395_);
  and (_12400_, _12168_, _12093_);
  or (_12401_, _12400_, _12165_);
  or (_12402_, _12401_, _12399_);
  or (_12403_, _12396_, _12166_);
  and (_12404_, _12403_, _12185_);
  and (_12405_, _12404_, _12402_);
  and (_12406_, _12206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_12407_, _12406_, _12387_);
  and (_12408_, _12204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_12409_, _12408_, _12209_);
  nand (_12410_, _12409_, _12407_);
  or (_12411_, _12210_, _12093_);
  and (_12412_, _12411_, _12410_);
  or (_12413_, _12412_, _12199_);
  or (_12414_, _12396_, _12265_);
  and (_12415_, _12414_, _12345_);
  and (_12416_, _12415_, _12413_);
  and (_12417_, _12197_, _12093_);
  or (_12418_, _12417_, _12194_);
  or (_12419_, _12418_, _12416_);
  and (_12420_, _12396_, _12271_);
  or (_12421_, _12420_, _12272_);
  and (_12422_, _12421_, _12419_);
  or (_12423_, _12422_, _12405_);
  and (_12424_, _12423_, _12255_);
  or (_12425_, _12424_, _12386_);
  and (_39002_[0], _12425_, _38997_);
  and (_12426_, _12316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_12427_, _12388_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_12428_, _12427_, _12391_);
  and (_12429_, _12162_, _12102_);
  or (_12430_, _12429_, _12428_);
  and (_12431_, _12430_, _12171_);
  not (_12432_, _12171_);
  or (_12433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_12434_, _12433_, _12432_);
  or (_12435_, _12434_, _12165_);
  or (_12436_, _12435_, _12431_);
  or (_12437_, _12166_, _12102_);
  and (_12438_, _12437_, _12185_);
  and (_12439_, _12438_, _12436_);
  and (_12440_, _12194_, _12102_);
  and (_12441_, _12433_, _12195_);
  or (_12442_, _12441_, _12201_);
  and (_12443_, _12209_, _12102_);
  or (_12444_, _12406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_12445_, _12444_, _12409_);
  or (_12446_, _12445_, _12375_);
  or (_12447_, _12446_, _12443_);
  and (_12448_, _12447_, _12442_);
  or (_12449_, _12448_, _12440_);
  and (_12450_, _12449_, _12271_);
  or (_12451_, _12450_, _12439_);
  and (_12452_, _12451_, _12255_);
  or (_12453_, _12452_, _12426_);
  and (_39002_[1], _12453_, _38997_);
  or (_12454_, _12218_, _12213_);
  and (_12455_, _12454_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_12456_, _12455_, _12236_);
  and (_39003_[0], _12456_, _38997_);
  and (_12457_, _12214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_12458_, _12457_, _12188_);
  and (_39004_[0], _12458_, _38997_);
  and (_12459_, _12075_, _34229_);
  or (_12460_, _12459_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_12461_, _12460_, _12086_);
  nand (_12462_, _12459_, _35722_);
  and (_12463_, _12462_, _12461_);
  and (_12464_, _12078_, _34149_);
  or (_12465_, _12464_, _12463_);
  and (_39009_[0], _12465_, _38997_);
  and (_12466_, _12075_, _11343_);
  or (_12467_, _12466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_12468_, _12467_, _12086_);
  nand (_12469_, _12466_, _35722_);
  and (_12470_, _12469_, _12468_);
  and (_12471_, _12078_, _34089_);
  or (_12472_, _12471_, _12470_);
  and (_39009_[1], _12472_, _38997_);
  and (_12473_, _12075_, _11370_);
  or (_12474_, _12473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_12475_, _12474_, _12086_);
  nand (_12476_, _12473_, _35722_);
  and (_12477_, _12476_, _12475_);
  nor (_12478_, _12086_, _34017_);
  or (_12479_, _12478_, _12477_);
  and (_39009_[2], _12479_, _38997_);
  and (_12480_, _11366_, _33604_);
  and (_12481_, _12480_, _34706_);
  and (_12482_, _12481_, _12048_);
  and (_12483_, _12482_, _34229_);
  or (_12484_, _12483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_12485_, _12484_, _12069_);
  nand (_12486_, _12483_, _35722_);
  and (_12487_, _12486_, _12485_);
  and (_12488_, _12068_, _34149_);
  or (_12489_, _12488_, _12487_);
  and (_39010_[0], _12489_, _38997_);
  not (_12490_, _33572_);
  nand (_12491_, _12482_, _33644_);
  or (_12492_, _12491_, _12490_);
  nor (_12493_, _12492_, _35722_);
  and (_12494_, _12492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_12495_, _12494_, _12068_);
  or (_12496_, _12495_, _12493_);
  or (_12497_, _12069_, _34122_);
  and (_12498_, _12497_, _38997_);
  and (_39010_[1], _12498_, _12496_);
  nand (_12499_, _12482_, _11359_);
  and (_12500_, _12499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_12501_, _12500_, _12068_);
  and (_12502_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_12503_, _12502_, _11345_);
  and (_12504_, _12503_, _12063_);
  or (_12505_, _12504_, _12501_);
  or (_12506_, _12069_, _34089_);
  and (_12507_, _12506_, _38997_);
  and (_39010_[2], _12507_, _12505_);
  and (_12508_, _12491_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_12509_, _12508_, _12068_);
  and (_12510_, _11359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_12511_, _12510_, _11357_);
  and (_12512_, _12511_, _12063_);
  or (_12513_, _12512_, _12509_);
  nand (_12514_, _12068_, _34052_);
  and (_12515_, _12514_, _38997_);
  and (_39010_[3], _12515_, _12513_);
  not (_12516_, _12482_);
  or (_12517_, _12516_, _11372_);
  and (_12518_, _12517_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_12519_, _12518_, _12068_);
  and (_12520_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_12521_, _12520_, _11376_);
  and (_12522_, _12521_, _12063_);
  or (_12523_, _12522_, _12519_);
  nand (_12524_, _12068_, _34017_);
  and (_12525_, _12524_, _38997_);
  and (_39010_[4], _12525_, _12523_);
  nand (_12526_, _12482_, _11383_);
  nor (_12527_, _12526_, _35722_);
  and (_12528_, _12526_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_12529_, _12528_, _12068_);
  or (_12530_, _12529_, _12527_);
  or (_12531_, _12069_, _33978_);
  and (_12532_, _12531_, _38997_);
  and (_39010_[5], _12532_, _12530_);
  nand (_12533_, _12482_, _11392_);
  and (_12534_, _12533_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_12535_, _12534_, _12068_);
  nor (_12536_, _12533_, _35722_);
  or (_12537_, _12536_, _12535_);
  or (_12538_, _12069_, _33942_);
  and (_12539_, _12538_, _38997_);
  and (_39010_[6], _12539_, _12537_);
  and (_12540_, _12048_, _11368_);
  and (_12541_, _12540_, _34229_);
  or (_12542_, _12541_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_12543_, _12542_, _12055_);
  nand (_12544_, _12541_, _35722_);
  and (_12545_, _12544_, _12543_);
  and (_12546_, _12054_, _34149_);
  or (_12547_, _12546_, _12545_);
  and (_39011_[0], _12547_, _38997_);
  nand (_12548_, _12540_, _33644_);
  or (_12549_, _12548_, _12490_);
  nor (_12550_, _12549_, _35722_);
  and (_12551_, _12052_, _11076_);
  and (_12552_, _12551_, _33632_);
  and (_12553_, _12549_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_12554_, _12553_, _12552_);
  or (_12555_, _12554_, _12550_);
  or (_12556_, _12055_, _34122_);
  and (_12557_, _12556_, _38997_);
  and (_39011_[1], _12557_, _12555_);
  nand (_12558_, _12049_, _11359_);
  and (_12559_, _12558_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_12560_, _12559_, _12054_);
  and (_12561_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_12562_, _12561_, _11345_);
  and (_12563_, _12562_, _12049_);
  or (_12564_, _12563_, _12560_);
  or (_12565_, _12055_, _34089_);
  and (_12566_, _12565_, _38997_);
  and (_39011_[2], _12566_, _12564_);
  and (_12567_, _12540_, _11357_);
  not (_12568_, _11074_);
  or (_12569_, _12548_, _12568_);
  and (_12570_, _12569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_12571_, _12570_, _12552_);
  or (_12572_, _12571_, _12567_);
  nand (_12573_, _12054_, _34052_);
  and (_12574_, _12573_, _38997_);
  and (_39011_[3], _12574_, _12572_);
  not (_12575_, _12049_);
  or (_12576_, _12575_, _11372_);
  and (_12577_, _12576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_12578_, _12577_, _12054_);
  and (_12579_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_12580_, _12579_, _11376_);
  and (_12581_, _12580_, _12049_);
  or (_12582_, _12581_, _12578_);
  nand (_12583_, _12054_, _34017_);
  and (_12584_, _12583_, _38997_);
  and (_39011_[4], _12584_, _12582_);
  and (_12585_, _12049_, _11383_);
  or (_12586_, _12585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_12587_, _12586_, _12055_);
  nand (_12588_, _12585_, _35722_);
  and (_12589_, _12588_, _12587_);
  and (_12590_, _12054_, _33978_);
  or (_12591_, _12590_, _12589_);
  and (_39011_[5], _12591_, _38997_);
  nand (_12592_, _12540_, _11392_);
  and (_12593_, _12592_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_12594_, _12593_, _12054_);
  nor (_12595_, _12592_, _35722_);
  or (_12596_, _12595_, _12594_);
  or (_12597_, _12055_, _33942_);
  and (_12598_, _12597_, _38997_);
  and (_39011_[6], _12598_, _12596_);
  and (_39029_, t2_i, _38997_);
  nor (_12599_, t2_i, rst);
  and (_39030_, _12599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand (_12600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _38997_);
  nor (_39031_, _12600_, t2ex_i);
  and (_39032_, t2ex_i, _38997_);
  and (_12601_, _34231_, _33605_);
  and (_12602_, _12601_, _11524_);
  nand (_12603_, _12602_, _34221_);
  and (_12604_, _12601_, _11401_);
  not (_12605_, _12604_);
  and (_12606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_12607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_12608_, _12607_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_12609_, _12608_, _12606_);
  not (_12610_, _12609_);
  and (_12611_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_12612_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_12613_, _12612_, _12611_);
  or (_12614_, _12613_, _12602_);
  and (_12615_, _12614_, _12605_);
  and (_12616_, _12615_, _12603_);
  and (_12617_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_12618_, _12617_, _12616_);
  and (_39033_[7], _12618_, _38997_);
  nand (_12619_, _12604_, _34221_);
  nor (_12620_, _12610_, _12602_);
  or (_12621_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_12622_, _12620_);
  or (_12623_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_12624_, _12623_, _12621_);
  or (_12625_, _12624_, _12604_);
  and (_12626_, _12625_, _38997_);
  and (_39034_[7], _12626_, _12619_);
  not (_12627_, _12607_);
  or (_12628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_12629_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_12630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _12629_);
  and (_12631_, _12630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_12632_, _12631_, _12628_);
  and (_12633_, _12601_, _11425_);
  and (_12634_, _12601_, _11486_);
  nor (_12635_, _12634_, _12633_);
  and (_12636_, _12635_, _12632_);
  and (_12637_, _12636_, _12627_);
  or (_12638_, _12637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_12639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12640_, _12639_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_12641_, _12640_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_12642_, _12641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_12643_, _12642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_12644_, _12643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12645_, _12644_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_12646_, _12645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_12647_, _12646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_12648_, _12647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_12649_, _12648_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_12650_, _12649_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_12651_, _12650_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_12652_, _12651_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_12653_, _12652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_12654_, _12653_);
  nand (_12655_, _12654_, _12637_);
  and (_12656_, _12655_, _38997_);
  and (_39035_, _12656_, _12638_);
  not (_12657_, _12634_);
  nor (_12658_, _12657_, _34221_);
  not (_12659_, _12608_);
  and (_12660_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_12661_, _12660_, _12632_);
  and (_12662_, _12661_, _12653_);
  nand (_12663_, _12644_, _12632_);
  nor (_12664_, _12663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  not (_12665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_12666_, _12606_, _12665_);
  nor (_12667_, _12666_, _12627_);
  and (_12668_, _12663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_12669_, _12668_, _12667_);
  or (_12670_, _12669_, _12664_);
  or (_12671_, _12670_, _12662_);
  not (_12672_, _12667_);
  or (_12673_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_12674_, _12673_, _12635_);
  and (_12675_, _12674_, _12671_);
  and (_12676_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_12677_, _12676_, _12675_);
  or (_12678_, _12677_, _12658_);
  and (_39036_[7], _12678_, _38997_);
  nand (_12679_, _12633_, _34221_);
  and (_12680_, _12667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_12681_, _12652_, _12632_);
  or (_12682_, _12681_, _12680_);
  and (_12683_, _12682_, _12657_);
  or (_12684_, _12683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_12685_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_12686_, _12685_, _12632_);
  nand (_12687_, _12686_, _12653_);
  and (_12688_, _12687_, _12672_);
  or (_12689_, _12680_, _12634_);
  or (_12690_, _12689_, _12688_);
  and (_12691_, _12690_, _12684_);
  or (_12692_, _12691_, _12633_);
  and (_12693_, _12692_, _38997_);
  and (_39037_[7], _12693_, _12679_);
  not (_12694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_12695_, _12635_, _12694_);
  and (_12696_, _12666_, _12607_);
  and (_12697_, _12696_, _12653_);
  and (_12698_, _12697_, _12636_);
  or (_12699_, _12698_, _12695_);
  and (_39038_, _12699_, _38997_);
  or (_12700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_12701_, _33630_, _34232_);
  and (_12702_, _12701_, _12062_);
  or (_12703_, _12702_, _12700_);
  not (_12704_, _11075_);
  nor (_12705_, _12704_, _35722_);
  nand (_12706_, _12704_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_12707_, _12706_, _12702_);
  or (_12708_, _12707_, _12705_);
  and (_12709_, _12708_, _12703_);
  and (_12710_, _12601_, _11091_);
  or (_12711_, _12710_, _12709_);
  nand (_12712_, _12710_, _34221_);
  and (_12713_, _12712_, _38997_);
  and (_39039_[7], _12713_, _12711_);
  or (_12714_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_12715_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12716_, _12715_, _12714_);
  or (_12717_, _12716_, _12602_);
  nand (_12718_, _12602_, _34148_);
  and (_12719_, _12718_, _12717_);
  or (_12720_, _12719_, _12604_);
  or (_12721_, _12605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_12722_, _12721_, _38997_);
  and (_39033_[0], _12722_, _12720_);
  not (_12723_, _12602_);
  or (_12724_, _12723_, _34122_);
  and (_12725_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_12726_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_12727_, _12726_, _12725_);
  or (_12728_, _12727_, _12602_);
  and (_12729_, _12728_, _12605_);
  and (_12730_, _12729_, _12724_);
  and (_12731_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_12732_, _12731_, _12730_);
  and (_39033_[1], _12732_, _38997_);
  or (_12733_, _12723_, _34089_);
  and (_12734_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_12735_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_12736_, _12735_, _12734_);
  or (_12737_, _12736_, _12602_);
  and (_12738_, _12737_, _12605_);
  and (_12739_, _12738_, _12733_);
  and (_12740_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_12741_, _12740_, _12739_);
  and (_39033_[2], _12741_, _38997_);
  nand (_12742_, _12602_, _34052_);
  and (_12743_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_12744_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_12745_, _12744_, _12743_);
  or (_12746_, _12745_, _12602_);
  and (_12747_, _12746_, _12605_);
  and (_12748_, _12747_, _12742_);
  and (_12749_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_12750_, _12749_, _12748_);
  and (_39033_[3], _12750_, _38997_);
  nand (_12751_, _12602_, _34017_);
  and (_12752_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12753_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_12754_, _12753_, _12752_);
  or (_12755_, _12754_, _12602_);
  and (_12756_, _12755_, _12605_);
  and (_12757_, _12756_, _12751_);
  and (_12758_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_12759_, _12758_, _12757_);
  and (_39033_[4], _12759_, _38997_);
  or (_12760_, _12723_, _33978_);
  and (_12761_, _12610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_12762_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_12763_, _12762_, _12761_);
  or (_12764_, _12763_, _12602_);
  and (_12765_, _12764_, _12605_);
  and (_12766_, _12765_, _12760_);
  and (_12767_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_12768_, _12767_, _12766_);
  and (_39033_[5], _12768_, _38997_);
  or (_12769_, _12723_, _33942_);
  not (_12770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_12771_, _12609_, _12770_);
  and (_12772_, _12609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_12773_, _12772_, _12771_);
  or (_12774_, _12773_, _12602_);
  and (_12775_, _12774_, _12605_);
  and (_12776_, _12775_, _12769_);
  and (_12777_, _12604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_12778_, _12777_, _12776_);
  and (_39033_[6], _12778_, _38997_);
  and (_12779_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_12780_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_12781_, _12780_, _12779_);
  or (_12782_, _12781_, _12604_);
  nand (_12783_, _12604_, _34148_);
  and (_12784_, _12783_, _38997_);
  and (_39034_[0], _12784_, _12782_);
  or (_12785_, _12605_, _34122_);
  and (_12786_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_12787_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_12788_, _12787_, _12786_);
  or (_12789_, _12788_, _12604_);
  and (_12790_, _12789_, _38997_);
  and (_39034_[1], _12790_, _12785_);
  or (_12791_, _12605_, _34089_);
  and (_12792_, _12622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_12793_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_12794_, _12793_, _12792_);
  or (_12795_, _12794_, _12604_);
  and (_12796_, _12795_, _38997_);
  and (_39034_[2], _12796_, _12791_);
  nand (_12797_, _12604_, _34052_);
  not (_12798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_12799_, _12620_, _12798_);
  and (_12800_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_12801_, _12800_, _12799_);
  or (_12802_, _12801_, _12604_);
  and (_12803_, _12802_, _38997_);
  and (_39034_[3], _12803_, _12797_);
  nand (_12804_, _12604_, _34017_);
  not (_12805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_12806_, _12620_, _12805_);
  and (_12807_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_12808_, _12807_, _12806_);
  or (_12809_, _12808_, _12604_);
  and (_12810_, _12809_, _38997_);
  and (_39034_[4], _12810_, _12804_);
  or (_12811_, _12605_, _33978_);
  or (_12812_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  not (_12813_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand (_12814_, _12620_, _12813_);
  and (_12815_, _12814_, _12812_);
  or (_12816_, _12815_, _12604_);
  and (_12817_, _12816_, _38997_);
  and (_39034_[5], _12817_, _12811_);
  or (_12818_, _12605_, _33942_);
  not (_12819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_12820_, _12620_, _12819_);
  and (_12821_, _12620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_12822_, _12821_, _12820_);
  or (_12823_, _12822_, _12604_);
  and (_12824_, _12823_, _38997_);
  and (_39034_[6], _12824_, _12818_);
  or (_12825_, _12632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12826_, _12632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  not (_12827_, _12826_);
  and (_12828_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_12829_, _12828_, _12653_);
  or (_12830_, _12829_, _12827_);
  and (_12831_, _12830_, _12825_);
  or (_12832_, _12831_, _12667_);
  or (_12833_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_12834_, _12833_, _12635_);
  and (_12835_, _12834_, _12832_);
  and (_12836_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12837_, _12634_, _34149_);
  or (_12838_, _12837_, _12836_);
  or (_12839_, _12838_, _12835_);
  and (_39036_[0], _12839_, _38997_);
  nor (_12840_, _12827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_12841_, _12827_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_12842_, _12841_, _12667_);
  or (_12843_, _12842_, _12840_);
  and (_12844_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_12845_, _12844_, _12632_);
  and (_12846_, _12845_, _12653_);
  or (_12847_, _12846_, _12843_);
  or (_12848_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_12849_, _12848_, _12635_);
  and (_12850_, _12849_, _12847_);
  and (_12851_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_12852_, _12634_, _34122_);
  or (_12853_, _12852_, _12851_);
  or (_12854_, _12853_, _12850_);
  and (_39036_[1], _12854_, _38997_);
  and (_12855_, _12634_, _34089_);
  and (_12856_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_12857_, _12653_, _12632_);
  and (_12858_, _12857_, _12856_);
  nand (_12859_, _12639_, _12632_);
  and (_12860_, _12859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_12861_, _12859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_12862_, _12861_, _12667_);
  or (_12863_, _12862_, _12860_);
  or (_12864_, _12863_, _12858_);
  or (_12865_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_12866_, _12865_, _12635_);
  and (_12867_, _12866_, _12864_);
  and (_12868_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_12869_, _12868_, _12867_);
  or (_12870_, _12869_, _12855_);
  and (_39036_[2], _12870_, _38997_);
  nor (_12871_, _12657_, _34052_);
  and (_12872_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_12873_, _12872_, _12857_);
  nand (_12874_, _12640_, _12632_);
  and (_12875_, _12874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_12876_, _12874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_12877_, _12876_, _12667_);
  or (_12878_, _12877_, _12875_);
  or (_12879_, _12878_, _12873_);
  or (_12880_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_12881_, _12880_, _12635_);
  and (_12882_, _12881_, _12879_);
  and (_12883_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_12884_, _12883_, _12882_);
  or (_12885_, _12884_, _12871_);
  and (_39036_[3], _12885_, _38997_);
  nor (_12886_, _12657_, _34017_);
  and (_12887_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12888_, _12887_, _12857_);
  nand (_12889_, _12641_, _12632_);
  and (_12890_, _12889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_12891_, _12889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_12892_, _12891_, _12667_);
  or (_12893_, _12892_, _12890_);
  or (_12894_, _12893_, _12888_);
  or (_12895_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12896_, _12895_, _12635_);
  and (_12897_, _12896_, _12894_);
  and (_12898_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_12899_, _12898_, _12897_);
  or (_12900_, _12899_, _12886_);
  and (_39036_[4], _12900_, _38997_);
  and (_12901_, _12634_, _33978_);
  and (_12902_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_12903_, _12902_, _12857_);
  nand (_12904_, _12642_, _12632_);
  and (_12905_, _12904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_12906_, _12904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_12907_, _12906_, _12667_);
  or (_12908_, _12907_, _12905_);
  or (_12909_, _12908_, _12903_);
  or (_12910_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_12911_, _12910_, _12635_);
  and (_12912_, _12911_, _12909_);
  and (_12913_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_12914_, _12913_, _12912_);
  or (_12915_, _12914_, _12901_);
  and (_39036_[5], _12915_, _38997_);
  and (_12916_, _12634_, _33942_);
  nor (_12917_, _12608_, _12770_);
  and (_12918_, _12917_, _12857_);
  and (_12919_, _12643_, _12632_);
  or (_12920_, _12919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12921_, _12920_, _12663_);
  or (_12922_, _12921_, _12667_);
  or (_12923_, _12922_, _12918_);
  nand (_12924_, _12667_, _12770_);
  and (_12925_, _12924_, _12635_);
  and (_12926_, _12925_, _12923_);
  and (_12927_, _12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_12928_, _12927_, _12926_);
  or (_12929_, _12928_, _12916_);
  and (_39036_[6], _12929_, _38997_);
  and (_12930_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_12931_, _12930_, _12857_);
  and (_12932_, _12645_, _12632_);
  or (_12933_, _12932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_12934_, _12932_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_12935_, _12934_, _12933_);
  or (_12936_, _12935_, _12667_);
  or (_12937_, _12936_, _12931_);
  or (_12938_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_12939_, _12938_, _12635_);
  and (_12940_, _12939_, _12937_);
  and (_12941_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_12942_, _12633_, _34149_);
  or (_12943_, _12942_, _12941_);
  or (_12944_, _12943_, _12940_);
  and (_39037_[0], _12944_, _38997_);
  nor (_12945_, _33657_, _33644_);
  and (_12946_, _12945_, _33572_);
  and (_12947_, _12601_, _12946_);
  and (_12948_, _12947_, _33662_);
  not (_12949_, _12948_);
  and (_12950_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_12951_, _12950_, _12857_);
  and (_12952_, _12646_, _12632_);
  or (_12953_, _12952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_12954_, _12952_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_12955_, _12954_, _12953_);
  or (_12956_, _12955_, _12667_);
  or (_12957_, _12956_, _12951_);
  nor (_12958_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_12959_, _12958_, _12634_);
  and (_12960_, _12959_, _12957_);
  and (_12961_, _12945_, _34228_);
  and (_12962_, _12601_, _12961_);
  and (_12963_, _12962_, _33662_);
  and (_12964_, _12963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_12965_, _12964_, _12960_);
  and (_12966_, _12965_, _12949_);
  and (_12967_, _12948_, _34122_);
  or (_12968_, _12967_, _12966_);
  and (_39037_[1], _12968_, _38997_);
  and (_12969_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_12970_, _12969_, _12857_);
  and (_12971_, _12647_, _12632_);
  or (_12972_, _12971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_12973_, _12971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_12974_, _12973_, _12972_);
  or (_12975_, _12974_, _12667_);
  or (_12976_, _12975_, _12970_);
  nor (_12977_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_12978_, _12977_, _12634_);
  and (_12979_, _12978_, _12976_);
  and (_12980_, _12963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_12981_, _12980_, _12979_);
  and (_12982_, _12981_, _12949_);
  and (_12983_, _12948_, _34089_);
  or (_12984_, _12983_, _12982_);
  and (_39037_[2], _12984_, _38997_);
  nor (_12985_, _12608_, _12798_);
  and (_12986_, _12985_, _12857_);
  nor (_12987_, _12973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_12988_, _12973_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_12989_, _12988_, _12667_);
  or (_12990_, _12989_, _12987_);
  or (_12991_, _12990_, _12986_);
  not (_12992_, _12635_);
  and (_12993_, _12667_, _12798_);
  nor (_12994_, _12993_, _12992_);
  and (_12995_, _12994_, _12991_);
  and (_12996_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_12997_, _12996_, _12995_);
  nor (_12998_, _12949_, _34052_);
  or (_12999_, _12998_, _12997_);
  and (_39037_[3], _12999_, _38997_);
  nor (_13000_, _12608_, _12805_);
  and (_13001_, _13000_, _12857_);
  nand (_13002_, _12649_, _12632_);
  nor (_13003_, _13002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_13004_, _13002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_13005_, _13004_, _12667_);
  or (_13006_, _13005_, _13003_);
  or (_13007_, _13006_, _13001_);
  nand (_13008_, _12667_, _12805_);
  and (_13009_, _13008_, _12635_);
  and (_13010_, _13009_, _13007_);
  and (_13011_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_13012_, _13011_, _13010_);
  nor (_13013_, _12949_, _34017_);
  or (_13014_, _13013_, _13012_);
  and (_39037_[4], _13014_, _38997_);
  and (_13015_, _12659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_13016_, _13015_, _12857_);
  and (_13017_, _12650_, _12632_);
  nor (_13018_, _13017_, _12813_);
  and (_13019_, _13017_, _12813_);
  or (_13020_, _13019_, _12667_);
  or (_13021_, _13020_, _13018_);
  or (_13022_, _13021_, _13016_);
  or (_13023_, _12672_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_13024_, _13023_, _12635_);
  and (_13025_, _13024_, _13022_);
  and (_13026_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_13027_, _13026_, _13025_);
  and (_13028_, _12633_, _33978_);
  or (_13029_, _13028_, _13027_);
  and (_39037_[5], _13029_, _38997_);
  and (_13030_, _12634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_13031_, _12608_, _12819_);
  and (_13032_, _13031_, _12857_);
  and (_13033_, _12651_, _12632_);
  nor (_13034_, _13033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_13035_, _13034_, _12681_);
  or (_13036_, _13035_, _12667_);
  or (_13037_, _13036_, _13032_);
  and (_13038_, _12667_, _12819_);
  nor (_13039_, _13038_, _12992_);
  and (_13040_, _13039_, _13037_);
  or (_13041_, _13040_, _13030_);
  and (_13042_, _12633_, _33942_);
  or (_13043_, _13042_, _13041_);
  and (_39037_[6], _13043_, _38997_);
  nand (_13044_, _12701_, _12481_);
  or (_13045_, _13044_, _11314_);
  nor (_13046_, _13045_, _35722_);
  and (_13047_, _13045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_13048_, _13047_, _12710_);
  or (_13049_, _13048_, _13046_);
  nand (_13050_, _12710_, _34148_);
  and (_13051_, _13050_, _38997_);
  and (_39039_[0], _13051_, _13049_);
  not (_13052_, _12710_);
  and (_13053_, _12702_, _34253_);
  or (_13054_, _13053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_13055_, _13054_, _13052_);
  nand (_13056_, _13053_, _35722_);
  and (_13057_, _13056_, _13055_);
  and (_13058_, _12710_, _34122_);
  or (_13059_, _13058_, _13057_);
  and (_39039_[1], _13059_, _38997_);
  or (_13060_, _13044_, _11358_);
  and (_13061_, _13060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_13062_, _13061_, _12710_);
  and (_13063_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_13064_, _13063_, _11345_);
  and (_13065_, _13064_, _12702_);
  or (_13066_, _13065_, _13062_);
  or (_13067_, _13052_, _34089_);
  and (_13068_, _13067_, _38997_);
  and (_39039_[2], _13068_, _13066_);
  or (_13069_, _13044_, _11073_);
  and (_13070_, _13069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_13071_, _13070_, _12710_);
  and (_13072_, _11359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_13073_, _13072_, _11357_);
  and (_13074_, _13073_, _12702_);
  or (_13075_, _13074_, _13071_);
  nand (_13076_, _12710_, _34052_);
  and (_13077_, _13076_, _38997_);
  and (_39039_[3], _13077_, _13075_);
  or (_13078_, _13044_, _11372_);
  and (_13079_, _13078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_13080_, _13079_, _12710_);
  and (_13081_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_13082_, _13081_, _11376_);
  and (_13083_, _13082_, _12702_);
  or (_13084_, _13083_, _13080_);
  nand (_13085_, _12710_, _34017_);
  and (_13086_, _13085_, _38997_);
  and (_39039_[4], _13086_, _13084_);
  and (_13087_, _12702_, _11383_);
  or (_13088_, _13087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_13089_, _13088_, _13052_);
  nand (_13090_, _13087_, _35722_);
  and (_13091_, _13090_, _13089_);
  and (_13092_, _12710_, _33978_);
  or (_13093_, _13092_, _13091_);
  and (_39039_[5], _13093_, _38997_);
  and (_13094_, _12606_, _12694_);
  or (_13095_, _13094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_13096_, _13095_, _12702_);
  not (_13097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_13098_, _11392_, _13097_);
  nand (_13099_, _13098_, _12702_);
  or (_13100_, _13099_, _12080_);
  and (_13101_, _13100_, _13096_);
  or (_13102_, _13101_, _12710_);
  or (_13103_, _13052_, _33942_);
  and (_13104_, _13103_, _38997_);
  and (_39039_[6], _13104_, _13102_);
  and (_13105_, _33657_, _33604_);
  and (_13106_, _13105_, _34706_);
  and (_13107_, _13106_, _11081_);
  and (_13108_, _11075_, _13107_);
  nand (_13109_, _13108_, _35722_);
  or (_13110_, _13108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_13111_, _13110_, _11083_);
  and (_13112_, _13111_, _13109_);
  and (_13113_, _34257_, _33633_);
  nand (_13114_, _13113_, _34221_);
  or (_13115_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_13116_, _13115_, _33662_);
  and (_13117_, _13116_, _13114_);
  not (_13118_, _33661_);
  and (_13119_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_13120_, _13119_, rst);
  or (_13121_, _13120_, _13117_);
  or (_39012_[7], _13121_, _13112_);
  nor (_13122_, _34251_, _33604_);
  and (_13123_, _13122_, _34706_);
  and (_13124_, _13123_, _11081_);
  and (_13125_, _13124_, _11075_);
  nand (_13126_, _13125_, _35722_);
  or (_13127_, _13125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_13128_, _13127_, _11083_);
  and (_13129_, _13128_, _13126_);
  and (_13130_, _11011_, _34257_);
  nand (_13131_, _13130_, _34221_);
  or (_13132_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_13133_, _13132_, _33662_);
  and (_13134_, _13133_, _13131_);
  and (_13135_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_13136_, _13135_, rst);
  or (_13137_, _13136_, _13134_);
  or (_39013_[7], _13137_, _13129_);
  and (_13138_, _12048_, _13106_);
  and (_13139_, _13138_, _11075_);
  nand (_13140_, _13139_, _35722_);
  or (_13141_, _13139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_13142_, _13141_, _11083_);
  and (_13143_, _13142_, _13140_);
  and (_13144_, _12067_, _34257_);
  nand (_13145_, _13144_, _34221_);
  or (_13146_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_13147_, _13146_, _33662_);
  and (_13148_, _13147_, _13145_);
  and (_13149_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_13150_, _13149_, rst);
  or (_13151_, _13150_, _13148_);
  or (_39014_[7], _13151_, _13143_);
  and (_13152_, _13123_, _12048_);
  and (_13153_, _13152_, _11075_);
  nand (_13154_, _13153_, _35722_);
  or (_13155_, _13153_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_13156_, _13155_, _11083_);
  and (_13157_, _13156_, _13154_);
  and (_13158_, _12052_, _34257_);
  and (_13159_, _13158_, _33632_);
  nand (_13160_, _13159_, _34221_);
  or (_13161_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_13162_, _13161_, _33662_);
  and (_13163_, _13162_, _13160_);
  and (_13164_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_13165_, _13164_, rst);
  or (_13166_, _13165_, _13163_);
  or (_39015_[7], _13166_, _13157_);
  nand (_13167_, _13113_, _35722_);
  or (_13168_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_13169_, _13168_, _11083_);
  and (_13170_, _13169_, _13167_);
  nand (_13171_, _13113_, _34148_);
  and (_13172_, _13168_, _33662_);
  and (_13173_, _13172_, _13171_);
  and (_13174_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_13175_, _13174_, rst);
  or (_13176_, _13175_, _13173_);
  or (_39012_[0], _13176_, _13170_);
  and (_13177_, _34259_, _33633_);
  nand (_13178_, _35722_, _13177_);
  or (_13179_, _13177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_13180_, _13179_, _11083_);
  and (_13181_, _13180_, _13178_);
  not (_13182_, _13113_);
  or (_13183_, _13182_, _34122_);
  or (_13184_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_13185_, _13184_, _33662_);
  and (_13186_, _13185_, _13183_);
  and (_13187_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_13188_, _13187_, rst);
  or (_13189_, _13188_, _13186_);
  or (_39012_[1], _13189_, _13181_);
  not (_13190_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_13191_, _11359_, _13107_);
  nor (_13192_, _13191_, _13190_);
  and (_13193_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_13194_, _13193_, _11345_);
  and (_13195_, _13194_, _13107_);
  or (_13196_, _13195_, _13192_);
  and (_13197_, _13196_, _11083_);
  or (_13198_, _13182_, _34089_);
  or (_13199_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_13200_, _13199_, _33662_);
  and (_13201_, _13200_, _13198_);
  nor (_13202_, _33661_, _13190_);
  or (_13203_, _13202_, rst);
  or (_13204_, _13203_, _13201_);
  or (_39012_[2], _13204_, _13197_);
  and (_13205_, _11356_, _13107_);
  nand (_13206_, _13205_, _35722_);
  or (_13207_, _13205_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_13208_, _13207_, _11083_);
  and (_13209_, _13208_, _13206_);
  nand (_13210_, _13113_, _34052_);
  or (_13211_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_13212_, _13211_, _33662_);
  and (_13213_, _13212_, _13210_);
  and (_13214_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_13215_, _13214_, rst);
  or (_13216_, _13215_, _13213_);
  or (_39012_[3], _13216_, _13209_);
  not (_13217_, _13107_);
  or (_13218_, _11372_, _13217_);
  and (_13219_, _13218_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_13220_, _11371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_13221_, _13220_, _11376_);
  and (_13222_, _13221_, _13107_);
  or (_13223_, _13222_, _13219_);
  and (_13224_, _13223_, _11083_);
  nand (_13225_, _13113_, _34017_);
  or (_13226_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_13227_, _13226_, _33662_);
  and (_13228_, _13227_, _13225_);
  and (_13229_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_13230_, _13229_, rst);
  or (_13231_, _13230_, _13228_);
  or (_39012_[4], _13231_, _13224_);
  and (_13232_, _11383_, _13107_);
  nand (_13233_, _13232_, _35722_);
  or (_13234_, _13232_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_13235_, _13234_, _11083_);
  and (_13236_, _13235_, _13233_);
  or (_13237_, _13182_, _33978_);
  or (_13238_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_13239_, _13238_, _33662_);
  and (_13240_, _13239_, _13237_);
  and (_13241_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_13242_, _13241_, rst);
  or (_13243_, _13242_, _13240_);
  or (_39012_[5], _13243_, _13236_);
  nand (_13244_, _11392_, _13107_);
  or (_13245_, _13244_, _35723_);
  not (_13246_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nand (_13247_, _13244_, _13246_);
  and (_13248_, _13247_, _11083_);
  and (_13249_, _13248_, _13245_);
  or (_13250_, _13182_, _33942_);
  or (_13251_, _13113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_13252_, _13251_, _33662_);
  and (_13253_, _13252_, _13250_);
  nor (_13254_, _33661_, _13246_);
  or (_13255_, _13254_, rst);
  or (_13256_, _13255_, _13253_);
  or (_39012_[6], _13256_, _13249_);
  nand (_13257_, _13130_, _35722_);
  or (_13258_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_13259_, _13258_, _11083_);
  and (_13260_, _13259_, _13257_);
  nand (_13261_, _13130_, _34148_);
  and (_13262_, _13258_, _33662_);
  and (_13263_, _13262_, _13261_);
  and (_13264_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_13265_, _13264_, rst);
  or (_13266_, _13265_, _13263_);
  or (_39013_[0], _13266_, _13260_);
  and (_13267_, _13124_, _34253_);
  nand (_13268_, _13267_, _35722_);
  or (_13269_, _13267_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_13270_, _13269_, _11083_);
  and (_13271_, _13270_, _13268_);
  not (_13272_, _13130_);
  or (_13273_, _13272_, _34122_);
  or (_13274_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_13275_, _13274_, _33662_);
  and (_13276_, _13275_, _13273_);
  and (_13277_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_13278_, _13277_, rst);
  or (_13279_, _13278_, _13276_);
  or (_39013_[1], _13279_, _13271_);
  and (_13280_, _13124_, _11343_);
  nand (_13281_, _13280_, _35722_);
  or (_13282_, _13280_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_13283_, _13282_, _11083_);
  and (_13284_, _13283_, _13281_);
  or (_13285_, _13272_, _34089_);
  or (_13286_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_13287_, _13286_, _33662_);
  and (_13288_, _13287_, _13285_);
  and (_13289_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_13290_, _13289_, rst);
  or (_13291_, _13290_, _13288_);
  or (_39013_[2], _13291_, _13284_);
  and (_13292_, _13124_, _11356_);
  nand (_13293_, _13292_, _35722_);
  or (_13294_, _13292_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_13295_, _13294_, _11083_);
  and (_13296_, _13295_, _13293_);
  nand (_13297_, _13130_, _34052_);
  or (_13298_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_13299_, _13298_, _33662_);
  and (_13300_, _13299_, _13297_);
  and (_13301_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_13302_, _13301_, rst);
  or (_13303_, _13302_, _13300_);
  or (_39013_[3], _13303_, _13296_);
  and (_13304_, _13124_, _11370_);
  nand (_13305_, _13304_, _35722_);
  or (_13306_, _13304_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_13307_, _13306_, _11083_);
  and (_13308_, _13307_, _13305_);
  nand (_13309_, _13130_, _34017_);
  or (_13310_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_13311_, _13310_, _33662_);
  and (_13312_, _13311_, _13309_);
  and (_13313_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_13314_, _13313_, rst);
  or (_13315_, _13314_, _13312_);
  or (_39013_[4], _13315_, _13308_);
  and (_13316_, _13124_, _11383_);
  nand (_13317_, _13316_, _35722_);
  or (_13318_, _13316_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_13319_, _13318_, _11083_);
  and (_13320_, _13319_, _13317_);
  or (_13321_, _13272_, _33978_);
  or (_13322_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_13323_, _13322_, _33662_);
  and (_13324_, _13323_, _13321_);
  and (_13325_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_13326_, _13325_, rst);
  or (_13327_, _13326_, _13324_);
  or (_39013_[5], _13327_, _13320_);
  nand (_13328_, _13124_, _11392_);
  or (_13329_, _13328_, _35723_);
  not (_13330_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nand (_13331_, _13328_, _13330_);
  and (_13332_, _13331_, _11083_);
  and (_13333_, _13332_, _13329_);
  or (_13334_, _13272_, _33942_);
  or (_13335_, _13130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_13336_, _13335_, _33662_);
  and (_13337_, _13336_, _13334_);
  nor (_13338_, _33661_, _13330_);
  or (_13339_, _13338_, rst);
  or (_13340_, _13339_, _13337_);
  or (_39013_[6], _13340_, _13333_);
  and (_13341_, _13138_, _34229_);
  nand (_13342_, _13341_, _35722_);
  or (_13343_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_13344_, _13343_, _11083_);
  and (_13345_, _13344_, _13342_);
  nand (_13346_, _13144_, _34148_);
  and (_13347_, _13343_, _33662_);
  and (_13348_, _13347_, _13346_);
  and (_13349_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_13350_, _13349_, rst);
  or (_13351_, _13350_, _13348_);
  or (_39014_[0], _13351_, _13345_);
  and (_13352_, _13138_, _34253_);
  nand (_13353_, _13352_, _35722_);
  or (_13354_, _13352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_13355_, _13354_, _11083_);
  and (_13356_, _13355_, _13353_);
  not (_13357_, _13144_);
  or (_13358_, _13357_, _34122_);
  or (_13359_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_13360_, _13359_, _33662_);
  and (_13361_, _13360_, _13358_);
  and (_13362_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_13363_, _13362_, rst);
  or (_13364_, _13363_, _13361_);
  or (_39014_[1], _13364_, _13356_);
  and (_13365_, _13138_, _11343_);
  nand (_13366_, _13365_, _35722_);
  or (_13367_, _13365_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_13368_, _13367_, _11083_);
  and (_13369_, _13368_, _13366_);
  or (_13370_, _13357_, _34089_);
  or (_13371_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_13372_, _13371_, _33662_);
  and (_13373_, _13372_, _13370_);
  and (_13374_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_13375_, _13374_, rst);
  or (_13376_, _13375_, _13373_);
  or (_39014_[2], _13376_, _13369_);
  and (_13377_, _13138_, _11356_);
  nand (_13378_, _13377_, _35722_);
  or (_13379_, _13377_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_13380_, _13379_, _11083_);
  and (_13381_, _13380_, _13378_);
  nand (_13382_, _13144_, _34052_);
  or (_13383_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_13384_, _13383_, _33662_);
  and (_13385_, _13384_, _13382_);
  and (_13386_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_13387_, _13386_, rst);
  or (_13388_, _13387_, _13385_);
  or (_39014_[3], _13388_, _13381_);
  and (_13389_, _13138_, _11370_);
  nand (_13390_, _13389_, _35722_);
  or (_13391_, _13389_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_13392_, _13391_, _11083_);
  and (_13393_, _13392_, _13390_);
  nand (_13394_, _13144_, _34017_);
  or (_13395_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_13396_, _13395_, _33662_);
  and (_13397_, _13396_, _13394_);
  and (_13398_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_13399_, _13398_, rst);
  or (_13400_, _13399_, _13397_);
  or (_39014_[4], _13400_, _13393_);
  and (_13401_, _13138_, _11383_);
  nand (_13402_, _13401_, _35722_);
  or (_13403_, _13401_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_13404_, _13403_, _11083_);
  and (_13405_, _13404_, _13402_);
  or (_13406_, _13357_, _33978_);
  or (_13407_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_13408_, _13407_, _33662_);
  and (_13409_, _13408_, _13406_);
  and (_13410_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_13411_, _13410_, rst);
  or (_13412_, _13411_, _13409_);
  or (_39014_[5], _13412_, _13405_);
  nand (_13413_, _13138_, _11392_);
  or (_13414_, _13413_, _35723_);
  not (_13415_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nand (_13416_, _13413_, _13415_);
  and (_13417_, _13416_, _11083_);
  and (_13418_, _13417_, _13414_);
  or (_13419_, _13357_, _33942_);
  or (_13420_, _13144_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_13421_, _13420_, _33662_);
  and (_13422_, _13421_, _13419_);
  nor (_13423_, _33661_, _13415_);
  or (_13424_, _13423_, rst);
  or (_13425_, _13424_, _13422_);
  or (_39014_[6], _13425_, _13418_);
  and (_13426_, _13152_, _34229_);
  nand (_13427_, _13426_, _35722_);
  or (_13428_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_13429_, _13428_, _11083_);
  and (_13430_, _13429_, _13427_);
  nand (_13431_, _13159_, _34148_);
  and (_13432_, _13428_, _33662_);
  and (_13433_, _13432_, _13431_);
  and (_13434_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_13435_, _13434_, rst);
  or (_13436_, _13435_, _13433_);
  or (_39015_[0], _13436_, _13430_);
  and (_13437_, _13152_, _34253_);
  nand (_13438_, _13437_, _35722_);
  or (_13439_, _13437_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_13440_, _13439_, _11083_);
  and (_13441_, _13440_, _13438_);
  not (_13442_, _13159_);
  or (_13443_, _13442_, _34122_);
  or (_13444_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_13445_, _13444_, _33662_);
  and (_13446_, _13445_, _13443_);
  and (_13447_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_13448_, _13447_, rst);
  or (_13449_, _13448_, _13446_);
  or (_39015_[1], _13449_, _13441_);
  and (_13450_, _13152_, _11343_);
  nand (_13451_, _13450_, _35722_);
  or (_13452_, _13450_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_13453_, _13452_, _11083_);
  and (_13454_, _13453_, _13451_);
  or (_13455_, _13442_, _34089_);
  or (_13456_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_13457_, _13456_, _33662_);
  and (_13458_, _13457_, _13455_);
  and (_13459_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_13460_, _13459_, rst);
  or (_13461_, _13460_, _13458_);
  or (_39015_[2], _13461_, _13454_);
  and (_13462_, _13152_, _11356_);
  nand (_13463_, _13462_, _35722_);
  or (_13464_, _13462_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_13465_, _13464_, _11083_);
  and (_13466_, _13465_, _13463_);
  nand (_13467_, _13159_, _34052_);
  or (_13468_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_13469_, _13468_, _33662_);
  and (_13470_, _13469_, _13467_);
  and (_13471_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_13472_, _13471_, rst);
  or (_13473_, _13472_, _13470_);
  or (_39015_[3], _13473_, _13466_);
  and (_13474_, _13152_, _11370_);
  nand (_13475_, _13474_, _35722_);
  or (_13476_, _13474_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_13477_, _13476_, _11083_);
  and (_13478_, _13477_, _13475_);
  nand (_13479_, _13159_, _34017_);
  or (_13480_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_13481_, _13480_, _33662_);
  and (_13482_, _13481_, _13479_);
  and (_13483_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_13484_, _13483_, rst);
  or (_13485_, _13484_, _13482_);
  or (_39015_[4], _13485_, _13478_);
  and (_13486_, _13152_, _11383_);
  nand (_13487_, _13486_, _35722_);
  or (_13488_, _13486_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_13489_, _13488_, _11083_);
  and (_13490_, _13489_, _13487_);
  or (_13491_, _13442_, _33978_);
  or (_13492_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_13493_, _13492_, _33662_);
  and (_13494_, _13493_, _13491_);
  and (_13495_, _13118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_13496_, _13495_, rst);
  or (_13497_, _13496_, _13494_);
  or (_39015_[5], _13497_, _13490_);
  nand (_13498_, _13152_, _11392_);
  or (_13499_, _13498_, _35723_);
  not (_13500_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nand (_13501_, _13498_, _13500_);
  and (_13502_, _13501_, _11083_);
  and (_13503_, _13502_, _13499_);
  or (_13504_, _13442_, _33942_);
  or (_13505_, _13159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_13506_, _13505_, _33662_);
  and (_13507_, _13506_, _13504_);
  nor (_13508_, _33661_, _13500_);
  or (_13509_, _13508_, rst);
  or (_13510_, _13509_, _13507_);
  or (_39015_[6], _13510_, _13503_);
  and (_13511_, _12701_, _11083_);
  and (_13512_, _13511_, _13123_);
  not (_13513_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_13514_, _11075_, _13513_);
  or (_13515_, _13514_, _12705_);
  and (_13516_, _13515_, _13512_);
  nor (_13517_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_13518_, _13517_);
  nand (_13519_, _13518_, _35722_);
  and (_13520_, _13517_, _13513_);
  nor (_13521_, _13520_, _13512_);
  and (_13522_, _13521_, _13519_);
  or (_13523_, _13522_, _34235_);
  or (_13524_, _13523_, _13516_);
  nand (_13525_, _34235_, _34221_);
  and (_13526_, _13525_, _38997_);
  and (_39016_[6], _13526_, _13524_);
  and (_13527_, _34235_, _34122_);
  and (_13528_, _13512_, _34253_);
  nand (_13529_, _13528_, _35722_);
  or (_13530_, _13528_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_13531_, _13530_, _34236_);
  and (_13532_, _13531_, _13529_);
  or (_13533_, _13532_, _13527_);
  and (_39016_[0], _13533_, _38997_);
  and (_13534_, _33930_, _33673_);
  not (_13535_, _13534_);
  nor (_13536_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_13537_, _13536_);
  and (_13538_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_13539_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_13540_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _13539_);
  not (_13541_, _13540_);
  or (_13542_, _13541_, _33987_);
  not (_13543_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_13544_, _13543_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_13545_, _13544_);
  or (_13546_, _13545_, _35601_);
  and (_13547_, _13546_, _13542_);
  nor (_13548_, _13544_, _13540_);
  or (_13549_, _34131_, _13539_);
  nand (_13550_, _13549_, _13548_);
  nand (_13551_, _13550_, _13547_);
  nand (_13552_, _13536_, _33778_);
  and (_13553_, _13552_, _13551_);
  and (_13554_, _13553_, _33815_);
  or (_13555_, _13541_, _33951_);
  or (_13556_, _13545_, _34035_);
  and (_13557_, _13556_, _13555_);
  or (_13558_, _34098_, _13539_);
  nand (_13559_, _13558_, _13548_);
  nand (_13560_, _13559_, _13557_);
  nand (_13561_, _13536_, _34196_);
  and (_13562_, _13561_, _13560_);
  and (_13563_, _13562_, _33884_);
  and (_13564_, _13563_, _13554_);
  and (_13565_, _13553_, _33884_);
  and (_13566_, _13562_, _33798_);
  nand (_13567_, _13566_, _13565_);
  and (_13568_, _13553_, _33798_);
  or (_13569_, _13568_, _13563_);
  and (_13570_, _13569_, _13567_);
  and (_13571_, _13570_, _13564_);
  or (_13572_, _13567_, _33765_);
  and (_13573_, _13553_, _33766_);
  not (_13574_, _13573_);
  nand (_13575_, _13574_, _13567_);
  and (_13576_, _13575_, _13566_);
  nand (_13577_, _13576_, _13572_);
  or (_13578_, _13573_, _13566_);
  and (_13579_, _13578_, _13577_);
  and (_13580_, _13579_, _13571_);
  not (_13581_, _13576_);
  nand (_13582_, _13561_, _13560_);
  or (_13583_, _13582_, _33765_);
  nand (_13584_, _13552_, _13551_);
  or (_13585_, _13584_, _34180_);
  or (_13586_, _13585_, _13583_);
  nand (_13587_, _13585_, _13583_);
  and (_13588_, _13587_, _13586_);
  nand (_13589_, _13588_, _13581_);
  or (_13590_, _13588_, _13581_);
  nand (_13591_, _13590_, _13589_);
  nand (_13592_, _13591_, _13580_);
  not (_13593_, _33831_);
  and (_13594_, _13562_, _13593_);
  and (_13595_, _13553_, _33865_);
  nand (_13596_, _13595_, _13594_);
  or (_13597_, _13584_, _33831_);
  and (_13598_, _13562_, _33865_);
  and (_13599_, _13598_, _13597_);
  nand (_13600_, _13599_, _13554_);
  nand (_13601_, _13600_, _13596_);
  not (_13602_, _13564_);
  and (_13603_, _13562_, _33815_);
  or (_13604_, _13603_, _13565_);
  and (_13605_, _13604_, _13602_);
  nand (_13606_, _13605_, _13601_);
  not (_13607_, _13606_);
  not (_13608_, _13571_);
  or (_13609_, _13570_, _13564_);
  and (_13610_, _13609_, _13608_);
  and (_13611_, _13610_, _13607_);
  nand (_13612_, _13579_, _13571_);
  or (_13613_, _13579_, _13571_);
  and (_13614_, _13613_, _13612_);
  nand (_13615_, _13614_, _13611_);
  not (_13616_, _13615_);
  or (_13617_, _13591_, _13580_);
  and (_13618_, _13617_, _13592_);
  nand (_13619_, _13618_, _13616_);
  and (_13620_, _13619_, _13592_);
  and (_13621_, _13553_, _35711_);
  and (_13622_, _13621_, _13594_);
  or (_13623_, _13595_, _13594_);
  and (_13624_, _13623_, _13596_);
  and (_13625_, _13624_, _13622_);
  or (_13626_, _13599_, _13554_);
  and (_13627_, _13626_, _13600_);
  nand (_13628_, _13627_, _13625_);
  not (_13629_, _13628_);
  or (_13630_, _13605_, _13601_);
  and (_13631_, _13630_, _13606_);
  nand (_13632_, _13631_, _13629_);
  not (_13633_, _13632_);
  nand (_13634_, _13610_, _13607_);
  or (_13635_, _13610_, _13607_);
  and (_13636_, _13635_, _13634_);
  nand (_13637_, _13636_, _13633_);
  not (_13638_, _13637_);
  or (_13639_, _13614_, _13611_);
  and (_13640_, _13639_, _13615_);
  and (_13641_, _13618_, _13640_);
  nand (_13642_, _13641_, _13638_);
  nand (_13643_, _13642_, _13620_);
  and (_13644_, _13562_, _35707_);
  and (_13645_, _13644_, _13574_);
  and (_13646_, _13588_, _13576_);
  and (_13647_, _13646_, _13645_);
  nor (_13648_, _13646_, _13645_);
  nor (_13649_, _13648_, _13647_);
  nand (_13650_, _13649_, _13643_);
  not (_13651_, _13647_);
  and (_13652_, _13651_, _13586_);
  nand (_13653_, _13652_, _13650_);
  nand (_13654_, _13653_, _13538_);
  and (_13655_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  or (_13656_, _13649_, _13643_);
  and (_13657_, _13656_, _13650_);
  nand (_13658_, _13657_, _13655_);
  or (_13659_, _13653_, _13538_);
  nand (_13660_, _13659_, _13654_);
  or (_13661_, _13660_, _13658_);
  nand (_13662_, _13661_, _13654_);
  and (_13663_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_13664_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_13665_, _13664_, _13663_);
  and (_13666_, _13665_, _13662_);
  and (_13667_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_13668_, _13640_, _13638_);
  nand (_13669_, _13668_, _13615_);
  nand (_13670_, _13618_, _13669_);
  or (_13671_, _13618_, _13669_);
  and (_13672_, _13671_, _13670_);
  nand (_13673_, _13672_, _13667_);
  or (_13674_, _13672_, _13667_);
  nand (_13675_, _13674_, _13673_);
  and (_13676_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_13677_, _13640_, _13638_);
  and (_13678_, _13677_, _13668_);
  nand (_13679_, _13678_, _13676_);
  or (_13680_, _13678_, _13676_);
  and (_13681_, _13680_, _13679_);
  and (_13682_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_13683_, _13636_, _13633_);
  and (_13684_, _13683_, _13637_);
  nand (_13685_, _13684_, _13682_);
  or (_13686_, _13684_, _13682_);
  nand (_13687_, _13686_, _13685_);
  and (_13688_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_13689_, _13631_, _13629_);
  and (_13690_, _13689_, _13632_);
  nand (_13691_, _13690_, _13688_);
  and (_13692_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_13693_, _13627_, _13625_);
  and (_13694_, _13693_, _13628_);
  nand (_13695_, _13694_, _13692_);
  and (_13696_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_13697_, _13624_, _13622_);
  or (_13698_, _13624_, _13622_);
  and (_13699_, _13698_, _13697_);
  and (_13700_, _13699_, _13696_);
  not (_13701_, _13700_);
  or (_13702_, _13694_, _13692_);
  nand (_13703_, _13702_, _13695_);
  or (_13704_, _13703_, _13701_);
  and (_13705_, _13704_, _13695_);
  or (_13706_, _13690_, _13688_);
  nand (_13707_, _13706_, _13691_);
  or (_13708_, _13707_, _13705_);
  and (_13709_, _13708_, _13691_);
  or (_13710_, _13709_, _13687_);
  nand (_13711_, _13710_, _13685_);
  nand (_13712_, _13711_, _13681_);
  and (_13713_, _13712_, _13679_);
  or (_13714_, _13713_, _13675_);
  and (_13715_, _13714_, _13673_);
  or (_13716_, _13657_, _13655_);
  and (_13717_, _13716_, _13658_);
  and (_13718_, _13659_, _13654_);
  and (_13719_, _13718_, _13717_);
  nand (_13720_, _13665_, _13719_);
  nor (_13721_, _13720_, _13715_);
  or (_13722_, _13721_, _13666_);
  and (_13723_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_13724_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_13725_, _13724_, _13723_);
  and (_13726_, _13725_, _13722_);
  and (_13727_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_13728_, _13727_, _13726_);
  and (_13729_, _13537_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_13730_, _13729_, _13728_);
  and (_13731_, _13728_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  or (_13732_, _13731_, _13730_);
  or (_13733_, _13732_, _13535_);
  nor (_13734_, _13727_, _13726_);
  nor (_13735_, _13734_, _13728_);
  and (_13736_, _13723_, _13722_);
  nor (_13737_, _13724_, _13736_);
  nor (_13738_, _13737_, _13726_);
  not (_13739_, _13717_);
  or (_13740_, _13739_, _13715_);
  not (_13741_, _13740_);
  and (_13742_, _13739_, _13715_);
  nor (_13743_, _13742_, _13741_);
  and (_13744_, _13740_, _13658_);
  or (_13745_, _13660_, _13744_);
  nand (_13746_, _13660_, _13744_);
  and (_13747_, _13746_, _13745_);
  or (_13748_, _13747_, _13743_);
  nand (_13749_, _13745_, _13654_);
  nand (_13750_, _13749_, _13663_);
  or (_13751_, _13749_, _13663_);
  and (_13752_, _13751_, _13750_);
  or (_13753_, _13752_, _13748_);
  nor (_13754_, _13723_, _13722_);
  nor (_13755_, _13754_, _13736_);
  or (_13756_, _13755_, _13753_);
  or (_13757_, _13756_, _13738_);
  or (_13758_, _13757_, _13735_);
  and (_13759_, _13758_, _13534_);
  or (_13760_, _35634_, _35632_);
  not (_13761_, _35584_);
  nand (_13762_, _35632_, _13761_);
  and (_13763_, _13762_, _35582_);
  and (_13764_, _13763_, _13760_);
  not (_13765_, _35672_);
  nor (_13766_, _13765_, _35670_);
  and (_13767_, _13765_, _35670_);
  or (_13768_, _13767_, _13766_);
  and (_13769_, _13768_, _35637_);
  nor (_13770_, _34131_, _34098_);
  and (_13771_, _35601_, _34035_);
  and (_13772_, _13771_, _13770_);
  and (_13773_, _33778_, _34196_);
  and (_13774_, _33921_, _33913_);
  and (_13775_, _33987_, _33951_);
  and (_13776_, _13775_, _13774_);
  and (_13777_, _13776_, _13773_);
  nand (_13778_, _13777_, _13772_);
  nand (_13779_, _13778_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_13780_, _13779_, _13769_);
  nor (_13781_, _13780_, _13764_);
  not (_13782_, _13664_);
  and (_13783_, _13782_, _13750_);
  nor (_13784_, _13783_, _13722_);
  nand (_13785_, _13784_, _13534_);
  nand (_13786_, _13785_, _13781_);
  nor (_13787_, _13786_, _13759_);
  nand (_13788_, _13787_, _13733_);
  nor (_13789_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_13790_, _13789_, _13512_);
  and (_13791_, _13790_, _13788_);
  and (_13792_, _11344_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_13793_, _13792_, _11345_);
  and (_13794_, _13793_, _13512_);
  or (_13795_, _13794_, _34235_);
  or (_13796_, _13795_, _13791_);
  or (_13797_, _34236_, _34089_);
  and (_13798_, _13797_, _38997_);
  and (_39016_[1], _13798_, _13796_);
  and (_13799_, _13512_, _11356_);
  nand (_13800_, _13799_, _35722_);
  or (_13801_, _13799_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_13802_, _13801_, _34236_);
  and (_13803_, _13802_, _13800_);
  or (_13804_, _13803_, _34282_);
  and (_39016_[2], _13804_, _38997_);
  and (_13805_, _13512_, _11370_);
  nand (_13806_, _13805_, _35722_);
  or (_13807_, _13805_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_13808_, _13807_, _34236_);
  and (_13809_, _13808_, _13806_);
  or (_13810_, _13809_, _34238_);
  and (_39016_[3], _13810_, _38997_);
  and (_13811_, _34235_, _33978_);
  and (_13812_, _13512_, _11383_);
  nand (_13813_, _13812_, _35722_);
  or (_13814_, _13812_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_13815_, _13814_, _34236_);
  and (_13816_, _13815_, _13813_);
  or (_13817_, _13816_, _13811_);
  and (_39016_[4], _13817_, _38997_);
  and (_13818_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_13819_, _13818_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_13820_, _35628_, _35582_);
  and (_13821_, _35658_, _35637_);
  nand (_13822_, _33935_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_13823_, _13822_, _13818_);
  or (_13824_, _13823_, _13821_);
  or (_13825_, _13824_, _13820_);
  and (_13826_, _13825_, _13819_);
  or (_13827_, _13826_, _13512_);
  not (_13828_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_13829_, _11392_, _13828_);
  nand (_13830_, _13829_, _13512_);
  or (_13831_, _13830_, _12080_);
  and (_13832_, _13831_, _13827_);
  or (_13833_, _13832_, _34235_);
  or (_13834_, _34236_, _33942_);
  and (_13835_, _13834_, _38997_);
  and (_39016_[5], _13835_, _13833_);
  nand (_13836_, _11074_, _33665_);
  not (_13837_, _13774_);
  nor (_13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_13839_, _13838_, _34180_);
  nor (_13840_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_13841_, _13840_);
  and (_13842_, _13841_, _13839_);
  not (_13843_, _13842_);
  or (_13844_, _34131_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_13845_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_13846_, _34062_, _13845_);
  and (_13847_, _13846_, _13844_);
  or (_13848_, _13847_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_13849_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_13850_, _34007_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_13851_, _33778_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_13852_, _13851_, _13850_);
  or (_13853_, _13852_, _13849_);
  and (_13854_, _13853_, _13848_);
  nor (_13855_, _13854_, _13843_);
  and (_13856_, _13854_, _13843_);
  nand (_13857_, _13838_, _33765_);
  nor (_13858_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_13859_, _13858_);
  and (_13860_, _13859_, _13857_);
  not (_13861_, _13860_);
  and (_13862_, _34098_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_13863_, _13862_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_13864_, _34035_, _13845_);
  nand (_13865_, _33951_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_13866_, _13865_, _13864_);
  or (_13867_, _13866_, _13849_);
  and (_13868_, _13867_, _13863_);
  or (_13869_, _13868_, _13861_);
  nor (_13870_, _13869_, _13856_);
  nor (_13871_, _13870_, _13855_);
  nor (_13872_, _13856_, _13855_);
  nand (_13873_, _13868_, _13861_);
  and (_13874_, _13873_, _13869_);
  and (_13875_, _13874_, _13872_);
  nand (_13876_, _13838_, _33797_);
  nor (_13877_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_13878_, _13877_);
  and (_13879_, _13878_, _13876_);
  and (_13880_, _34131_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_13881_, _13880_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_13882_, _34062_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_13883_, _34007_, _13845_);
  and (_13884_, _13883_, _13882_);
  or (_13885_, _13884_, _13849_);
  nand (_13886_, _13885_, _13881_);
  and (_13887_, _13886_, _13879_);
  not (_13888_, _13887_);
  or (_13889_, _34098_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_13890_, _34035_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_13891_, _13890_, _13889_);
  and (_13892_, _13891_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_13893_, _13892_);
  nand (_13894_, _13838_, _33883_);
  nor (_13895_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_13896_, _13895_);
  and (_13897_, _13896_, _13894_);
  and (_13898_, _13897_, _13893_);
  not (_13899_, _13898_);
  nor (_13900_, _13886_, _13879_);
  or (_13901_, _13900_, _13887_);
  or (_13902_, _13901_, _13899_);
  nand (_13903_, _13902_, _13888_);
  nand (_13904_, _13903_, _13875_);
  and (_13905_, _13904_, _13871_);
  and (_13906_, _13847_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_13907_, _13906_);
  nor (_13908_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_13909_, _13908_);
  nand (_13910_, _13838_, _33814_);
  and (_13911_, _13910_, _13909_);
  nand (_13912_, _13911_, _13907_);
  or (_13913_, _13911_, _13907_);
  nand (_13914_, _13913_, _13912_);
  and (_13915_, _13862_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_13916_, _13915_);
  not (_13917_, _13838_);
  or (_13918_, _13917_, _33865_);
  nor (_13919_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_13920_, _13919_);
  and (_13921_, _13920_, _13918_);
  nand (_13922_, _13921_, _13916_);
  and (_13923_, _13880_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_13924_, _13923_);
  nand (_13925_, _13838_, _33831_);
  nor (_13926_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_13927_, _13926_);
  and (_13928_, _13927_, _13925_);
  nor (_13929_, _13928_, _13924_);
  or (_13930_, _13921_, _13916_);
  nand (_13931_, _13930_, _13922_);
  or (_13932_, _13931_, _13929_);
  and (_13933_, _13932_, _13922_);
  or (_13934_, _13933_, _13914_);
  nand (_13935_, _13934_, _13912_);
  or (_13936_, _13897_, _13893_);
  and (_13937_, _13936_, _13899_);
  not (_13938_, _13901_);
  and (_13939_, _13938_, _13937_);
  and (_13940_, _13939_, _13875_);
  nand (_13941_, _13940_, _13935_);
  nand (_13942_, _13941_, _13905_);
  nor (_13943_, _13891_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_13944_, _33951_, _13845_);
  and (_13945_, _34196_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_13946_, _13945_, _13944_);
  nor (_13947_, _13946_, _13849_);
  nor (_13948_, _13947_, _13943_);
  not (_13949_, _13948_);
  nor (_13950_, _13773_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_13951_, _13866_, _13852_);
  nor (_13952_, _13946_, _13884_);
  and (_13953_, _13952_, _13951_);
  nor (_13954_, _13953_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_13955_, _13954_, _13950_);
  and (_13956_, _13955_, _13949_);
  and (_13957_, _13956_, _13942_);
  nor (_13958_, _13957_, _13843_);
  not (_13959_, _13874_);
  and (_13960_, _13937_, _13935_);
  nor (_13961_, _13960_, _13898_);
  or (_13962_, _13961_, _13900_);
  and (_13963_, _13962_, _13888_);
  or (_13964_, _13963_, _13959_);
  and (_13965_, _13964_, _13869_);
  nand (_13966_, _13965_, _13872_);
  or (_13967_, _13965_, _13872_);
  nand (_13968_, _13967_, _13966_);
  and (_13969_, _13968_, _13957_);
  nor (_13970_, _13969_, _13958_);
  not (_13971_, _13854_);
  and (_13972_, _13963_, _13959_);
  not (_13973_, _13972_);
  nand (_13974_, _13973_, _13964_);
  nand (_13975_, _13974_, _13957_);
  nor (_13976_, _13957_, _13860_);
  not (_13977_, _13976_);
  and (_13978_, _13977_, _13975_);
  nand (_13979_, _13978_, _13971_);
  or (_13980_, _13978_, _13971_);
  and (_13981_, _13980_, _13979_);
  not (_13982_, _13868_);
  nand (_13983_, _13901_, _13961_);
  or (_13984_, _13901_, _13961_);
  nand (_13985_, _13984_, _13983_);
  nand (_13986_, _13985_, _13957_);
  nor (_13987_, _13957_, _13879_);
  not (_13988_, _13987_);
  and (_13989_, _13988_, _13986_);
  and (_13990_, _13989_, _13982_);
  not (_13991_, _13957_);
  nor (_13992_, _13937_, _13935_);
  nor (_13993_, _13992_, _13960_);
  nor (_13994_, _13993_, _13991_);
  nor (_13995_, _13957_, _13897_);
  nor (_13996_, _13995_, _13994_);
  and (_13997_, _13996_, _13886_);
  not (_13998_, _13997_);
  nor (_13999_, _13989_, _13982_);
  or (_14000_, _13990_, _13999_);
  nor (_14001_, _14000_, _13998_);
  or (_14002_, _14001_, _13990_);
  and (_14003_, _13933_, _13914_);
  not (_14004_, _14003_);
  and (_14005_, _14004_, _13934_);
  or (_14006_, _14005_, _13991_);
  or (_14007_, _13957_, _13911_);
  and (_14008_, _14007_, _14006_);
  nor (_14009_, _14008_, _13893_);
  not (_14010_, _14009_);
  nand (_14011_, _13991_, _13928_);
  nor (_14012_, _13928_, _13923_);
  and (_14013_, _13928_, _13923_);
  nor (_14014_, _14013_, _14012_);
  nand (_14015_, _13957_, _14014_);
  nand (_14016_, _14015_, _14011_);
  nand (_14017_, _14016_, _13916_);
  or (_14018_, _14016_, _13916_);
  nand (_14019_, _14018_, _14017_);
  nor (_14020_, _13838_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_14021_, _13838_, _33848_);
  nor (_14022_, _14021_, _14020_);
  nor (_14023_, _14022_, _13924_);
  or (_14024_, _14023_, _14019_);
  and (_14025_, _14024_, _14017_);
  and (_14026_, _13931_, _13929_);
  not (_14027_, _14026_);
  and (_14028_, _14027_, _13932_);
  or (_14029_, _14028_, _13991_);
  or (_14030_, _13957_, _13921_);
  and (_14031_, _14030_, _14029_);
  nand (_14032_, _14031_, _13907_);
  or (_14033_, _14031_, _13907_);
  and (_14034_, _14033_, _14032_);
  not (_14035_, _14034_);
  or (_14036_, _14035_, _14025_);
  and (_14037_, _14008_, _13893_);
  not (_14038_, _14037_);
  and (_14039_, _14038_, _14032_);
  nand (_14040_, _14039_, _14036_);
  and (_14041_, _14040_, _14010_);
  nor (_14042_, _13996_, _13886_);
  nor (_14043_, _14042_, _13997_);
  not (_14044_, _14000_);
  and (_14045_, _14044_, _14043_);
  and (_14046_, _14045_, _14041_);
  or (_14047_, _14046_, _14002_);
  nand (_14048_, _14047_, _13981_);
  or (_14049_, _13970_, _13948_);
  and (_14050_, _14049_, _13979_);
  nand (_14051_, _14050_, _14048_);
  and (_14052_, _13970_, _13948_);
  not (_14053_, _14052_);
  and (_14054_, _14053_, _13955_);
  and (_14055_, _14054_, _14051_);
  or (_14056_, _14055_, _13970_);
  nand (_14057_, _14054_, _14051_);
  and (_14058_, _14053_, _14049_);
  and (_14059_, _14048_, _13979_);
  or (_14060_, _14059_, _14058_);
  nand (_14061_, _14059_, _14058_);
  and (_14062_, _14061_, _14060_);
  or (_14063_, _14062_, _14057_);
  and (_14064_, _14063_, _14056_);
  or (_14065_, _14064_, _13837_);
  nor (_14066_, _34183_, _34180_);
  nor (_14067_, _14066_, _35691_);
  and (_14068_, _14067_, _33734_);
  nor (_14069_, _14068_, _35693_);
  and (_14070_, _14069_, _34180_);
  nor (_14071_, _14069_, _34180_);
  nor (_14072_, _14071_, _14070_);
  nor (_14073_, _14072_, _35696_);
  and (_14074_, _35712_, _33888_);
  not (_14075_, _14074_);
  and (_14076_, _33935_, _35707_);
  not (_14077_, _14076_);
  and (_14078_, _35681_, _35711_);
  nor (_14079_, _14078_, _33929_);
  and (_14080_, _14079_, _14077_);
  and (_14081_, _14080_, _34212_);
  and (_14082_, _14081_, _34209_);
  and (_14083_, _14082_, _14075_);
  not (_14084_, _14083_);
  nor (_14085_, _14084_, _14073_);
  and (_14086_, _14085_, _34203_);
  and (_14087_, _35632_, _35639_);
  nor (_14088_, _35632_, _35639_);
  nor (_14089_, _14088_, _14087_);
  and (_14090_, _14089_, _35582_);
  and (_14091_, _35670_, _35639_);
  not (_14092_, _14091_);
  nor (_14093_, _35671_, _35638_);
  and (_14094_, _14093_, _14092_);
  nor (_14095_, _14094_, _14090_);
  and (_14096_, _14095_, _14086_);
  and (_14097_, _14096_, _13733_);
  and (_14098_, _14097_, _14065_);
  nor (_14099_, _14098_, _13836_);
  and (_14100_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _33129_);
  and (_14101_, _14100_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_14102_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_14103_, _14102_, _14101_);
  or (_14104_, _14103_, _14099_);
  nor (_14105_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_14106_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_14107_, _14106_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14108_, _14107_, _14105_);
  nor (_14109_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_14110_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_14111_, _14110_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14112_, _14111_, _14109_);
  not (_14113_, _14112_);
  nor (_14114_, _14113_, _35672_);
  nor (_14115_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_14116_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_14117_, _14116_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14118_, _14117_, _14115_);
  and (_14119_, _14118_, _14114_);
  nor (_14120_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_14121_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_14122_, _14121_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14123_, _14122_, _14120_);
  and (_14124_, _14123_, _14119_);
  and (_14125_, _14124_, _14108_);
  nor (_14126_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_14127_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_14128_, _14127_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14129_, _14128_, _14126_);
  and (_14130_, _14129_, _14125_);
  nor (_14131_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_14132_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_14133_, _14132_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14134_, _14133_, _14131_);
  and (_14135_, _14134_, _14130_);
  nor (_14136_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_14137_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_14138_, _14137_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14139_, _14138_, _14136_);
  nand (_14140_, _14139_, _14135_);
  nor (_14141_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_14142_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_14143_, _14142_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_14144_, _14143_, _14141_);
  and (_14145_, _14144_, _14140_);
  nor (_14146_, _14144_, _14140_);
  or (_14147_, _14146_, _14145_);
  nand (_14148_, _14147_, _35637_);
  and (_14149_, _13713_, _13675_);
  not (_14150_, _14149_);
  and (_14151_, _14150_, _13714_);
  and (_14152_, _14151_, _13534_);
  nor (_14153_, _34132_, _34180_);
  and (_14154_, _14153_, _34181_);
  and (_14155_, _14154_, _34098_);
  and (_14156_, _14155_, _34062_);
  and (_14157_, _35623_, _33734_);
  and (_14158_, _14157_, _14156_);
  nor (_14159_, _35587_, _33734_);
  and (_14160_, _34184_, _34180_);
  and (_14161_, _13772_, _14160_);
  and (_14162_, _14161_, _33987_);
  and (_14163_, _14162_, _14159_);
  or (_14164_, _14163_, _14158_);
  and (_14165_, _33951_, _33734_);
  and (_14166_, _33987_, _33734_);
  nor (_14167_, _14166_, _14165_);
  and (_14168_, _14167_, _14164_);
  and (_14169_, _33778_, _33734_);
  nor (_14170_, _14169_, _33779_);
  and (_14171_, _14170_, _14168_);
  and (_14172_, _14171_, _34197_);
  nor (_14173_, _14171_, _34197_);
  nor (_14174_, _14173_, _14172_);
  and (_14175_, _14174_, _33899_);
  and (_14176_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_14177_, _34197_, _33734_);
  nor (_14178_, _14177_, _35697_);
  nor (_14179_, _14178_, _34006_);
  and (_14180_, _35708_, _33815_);
  and (_14181_, _33935_, _34197_);
  or (_14182_, _14181_, _14180_);
  or (_14183_, _14182_, _14179_);
  nor (_14184_, _14183_, _14176_);
  not (_14185_, _14184_);
  nor (_14186_, _14185_, _14175_);
  not (_14187_, _14186_);
  nor (_14188_, _14187_, _14152_);
  and (_14189_, _14188_, _14148_);
  nand (_14190_, _14189_, _14101_);
  and (_14191_, _14190_, _38997_);
  and (_38993_[7], _14191_, _14104_);
  and (_14192_, _11342_, _33665_);
  nor (_14193_, _14192_, _14101_);
  not (_14194_, _14193_);
  nand (_14195_, _14194_, _14098_);
  or (_14196_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_14197_, _14196_, _38997_);
  and (_38994_[7], _14197_, _14195_);
  not (_14198_, _14022_);
  and (_14199_, _14055_, _13923_);
  nor (_14200_, _14199_, _14198_);
  and (_14201_, _14199_, _14198_);
  or (_14202_, _14201_, _14200_);
  nand (_14203_, _14202_, _13774_);
  and (_14204_, _13743_, _13534_);
  and (_14205_, _35648_, _33734_);
  nor (_14206_, _14205_, _35649_);
  nand (_14207_, _14206_, _35582_);
  nor (_14208_, _35696_, _33848_);
  and (_14209_, _35708_, _33888_);
  nor (_14210_, _14209_, _14208_);
  nand (_14211_, _14206_, _35637_);
  and (_14212_, _35675_, _35707_);
  or (_14213_, _34213_, _33831_);
  nand (_14214_, _33935_, _35711_);
  nand (_14215_, _14214_, _14213_);
  nor (_14216_, _14215_, _14212_);
  and (_14217_, _14216_, _34145_);
  and (_14218_, _14217_, _14211_);
  and (_14219_, _14218_, _14210_);
  and (_14220_, _14219_, _14207_);
  not (_14221_, _14220_);
  nor (_14222_, _14221_, _14204_);
  nand (_14223_, _14222_, _14203_);
  not (_14224_, _14223_);
  nor (_14225_, _14224_, _13836_);
  and (_14226_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_14227_, _14226_, _14101_);
  or (_14228_, _14227_, _14225_);
  not (_14229_, _14101_);
  and (_14230_, _34131_, _33935_);
  and (_14231_, _35708_, _33884_);
  nor (_14232_, _35697_, _34200_);
  not (_14233_, _14232_);
  nor (_14234_, _14233_, _34186_);
  nor (_14235_, _14234_, _34131_);
  and (_14236_, _14234_, _34131_);
  or (_14237_, _14236_, _34100_);
  nor (_14238_, _14237_, _14235_);
  nor (_14239_, _34006_, _33848_);
  or (_14240_, _14239_, _14238_);
  or (_14241_, _14240_, _14231_);
  and (_14242_, _14055_, _13774_);
  and (_14243_, _14113_, _35672_);
  nor (_14244_, _14243_, _14114_);
  and (_14245_, _14244_, _35637_);
  and (_14246_, _13621_, _13534_);
  or (_14247_, _14246_, _14245_);
  or (_14248_, _14247_, _14242_);
  or (_14249_, _14248_, _14241_);
  or (_14250_, _14249_, _14230_);
  or (_14251_, _14250_, _14229_);
  and (_14252_, _14251_, _38997_);
  and (_38993_[0], _14252_, _14228_);
  nand (_14253_, _13747_, _13534_);
  and (_14254_, _14023_, _14019_);
  not (_14255_, _14254_);
  and (_14256_, _14255_, _14024_);
  or (_14257_, _14256_, _14057_);
  or (_14258_, _14055_, _14016_);
  and (_14259_, _14258_, _14257_);
  nand (_14260_, _14259_, _13774_);
  nor (_14261_, _34134_, _34111_);
  or (_14262_, _14261_, _35641_);
  and (_14263_, _14262_, _35649_);
  nor (_14264_, _14262_, _35649_);
  or (_14265_, _14264_, _14263_);
  and (_14266_, _14265_, _35637_);
  nor (_14267_, _35619_, _35618_);
  nor (_14268_, _14267_, _35620_);
  nor (_14269_, _14268_, _35583_);
  nor (_14270_, _14269_, _14266_);
  nor (_14271_, _35690_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_14272_, _14271_, _13593_);
  nor (_14273_, _14271_, _13593_);
  nor (_14274_, _14273_, _14272_);
  nor (_14275_, _14274_, _35696_);
  or (_14276_, _33928_, _33848_);
  nand (_14277_, _33934_, _33865_);
  not (_14278_, _14277_);
  and (_14279_, _33935_, _13593_);
  nor (_14280_, _14279_, _14278_);
  and (_14281_, _14280_, _14276_);
  and (_14282_, _14281_, _34116_);
  and (_14283_, _14282_, _34113_);
  not (_14284_, _14283_);
  nor (_14285_, _14284_, _14275_);
  and (_14286_, _14285_, _34106_);
  and (_14287_, _14286_, _14270_);
  and (_14288_, _14287_, _14260_);
  nand (_14289_, _14288_, _14253_);
  not (_14290_, _14289_);
  nor (_14291_, _14290_, _13836_);
  and (_14292_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_14293_, _14292_, _14101_);
  or (_14294_, _14293_, _14291_);
  nor (_14295_, _14118_, _14114_);
  nor (_14296_, _14295_, _14119_);
  and (_14297_, _14296_, _35637_);
  not (_14298_, _14297_);
  and (_14299_, _13957_, _13774_);
  not (_14300_, _14299_);
  and (_14301_, _14154_, _33734_);
  and (_14302_, _34132_, _14160_);
  and (_14303_, _14302_, _33888_);
  nor (_14304_, _14303_, _14301_);
  nor (_14305_, _14304_, _34098_);
  and (_14306_, _14304_, _34098_);
  nor (_14307_, _14306_, _14305_);
  nor (_14308_, _14307_, _34100_);
  and (_14309_, _34098_, _33935_);
  and (_14310_, _13562_, _35711_);
  not (_14311_, _14310_);
  and (_14312_, _14311_, _13597_);
  nor (_14313_, _14312_, _13622_);
  and (_14314_, _14313_, _13534_);
  and (_14315_, _35708_, _33798_);
  nor (_14316_, _34006_, _33831_);
  or (_14317_, _14316_, _14315_);
  or (_14318_, _14317_, _14314_);
  nor (_14319_, _14318_, _14309_);
  not (_14320_, _14319_);
  nor (_14321_, _14320_, _14308_);
  and (_14322_, _14321_, _14300_);
  and (_14323_, _14322_, _14298_);
  nand (_14324_, _14323_, _14101_);
  and (_14325_, _14324_, _38997_);
  and (_38993_[1], _14325_, _14294_);
  nand (_14326_, _13752_, _13534_);
  not (_14327_, _14036_);
  and (_14328_, _14035_, _14025_);
  nor (_14329_, _14328_, _14327_);
  or (_14330_, _14329_, _14057_);
  or (_14331_, _14055_, _14031_);
  and (_14332_, _14331_, _14330_);
  nand (_14333_, _14332_, _13774_);
  nor (_14334_, _35620_, _35615_);
  nor (_14335_, _14334_, _35621_);
  nor (_14336_, _14335_, _35583_);
  or (_14337_, _34213_, _33814_);
  and (_14338_, _33935_, _33865_);
  nor (_14339_, _34117_, _14338_);
  and (_14340_, _14339_, _14337_);
  and (_14341_, _14340_, _34082_);
  and (_14342_, _14341_, _34079_);
  not (_14343_, _14342_);
  nor (_14344_, _14343_, _14336_);
  nor (_14345_, _35652_, _35650_);
  nor (_14346_, _14345_, _35638_);
  and (_14347_, _14346_, _35654_);
  and (_14348_, _35689_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_14349_, _14273_, _34064_);
  nor (_14350_, _14349_, _14348_);
  nor (_14351_, _14350_, _35696_);
  nor (_14352_, _14351_, _14347_);
  and (_14353_, _14352_, _14344_);
  and (_14354_, _14353_, _34073_);
  and (_14355_, _14354_, _14333_);
  and (_14356_, _14355_, _14326_);
  nor (_14357_, _14356_, _13836_);
  and (_14358_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_14359_, _14358_, _14101_);
  or (_14360_, _14359_, _14357_);
  nor (_14361_, _14123_, _14119_);
  nor (_14362_, _14361_, _14124_);
  and (_14363_, _14362_, _35637_);
  not (_14364_, _14363_);
  and (_14365_, _14302_, _34107_);
  and (_14366_, _14365_, _33888_);
  and (_14367_, _14155_, _33734_);
  nor (_14368_, _14367_, _14366_);
  and (_14369_, _14368_, _35601_);
  nor (_14370_, _14368_, _35601_);
  or (_14371_, _14370_, _34100_);
  nor (_14372_, _14371_, _14369_);
  nor (_14373_, _13699_, _13696_);
  nor (_14374_, _14373_, _13700_);
  and (_14375_, _14374_, _13534_);
  and (_14376_, _34062_, _33935_);
  and (_14377_, _35708_, _33766_);
  and (_14378_, _33674_, _33865_);
  and (_14379_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_14380_, _14379_, _14378_);
  or (_14381_, _14380_, _14377_);
  nor (_14382_, _14381_, _14376_);
  not (_14383_, _14382_);
  nor (_14384_, _14383_, _14375_);
  not (_14385_, _14384_);
  nor (_14386_, _14385_, _14372_);
  and (_14387_, _14386_, _14364_);
  nand (_14388_, _14387_, _14101_);
  and (_14389_, _14388_, _38997_);
  and (_38993_[2], _14389_, _14360_);
  not (_14390_, _14008_);
  or (_14391_, _14055_, _14390_);
  or (_14392_, _14037_, _14009_);
  and (_14393_, _14036_, _14032_);
  and (_14394_, _14393_, _14392_);
  nor (_14395_, _14393_, _14392_);
  or (_14396_, _14395_, _14394_);
  or (_14397_, _14396_, _14057_);
  nand (_14398_, _14397_, _14391_);
  nand (_14399_, _14398_, _13774_);
  nor (_14400_, _35621_, _35612_);
  nor (_14401_, _14400_, _35622_);
  nor (_14402_, _14401_, _35583_);
  not (_14403_, _14402_);
  and (_14404_, _35654_, _35647_);
  or (_14405_, _14404_, _35638_);
  nor (_14406_, _14405_, _35655_);
  not (_14407_, _14406_);
  nor (_14408_, _35689_, _13828_);
  nor (_14409_, _14408_, _33815_);
  and (_14410_, _33935_, _33815_);
  nor (_14411_, _35690_, _35696_);
  nor (_14412_, _14411_, _14410_);
  nor (_14413_, _14412_, _14409_);
  or (_14414_, _34213_, _33883_);
  not (_14415_, _34083_);
  and (_14416_, _14415_, _14414_);
  not (_14417_, _14416_);
  nor (_14418_, _14417_, _14413_);
  and (_14419_, _14418_, _34051_);
  and (_14420_, _14419_, _14407_);
  and (_14421_, _14420_, _14403_);
  and (_14422_, _14421_, _14399_);
  and (_14423_, _14422_, _13785_);
  nor (_14424_, _14423_, _13836_);
  and (_14425_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_14426_, _14425_, _14101_);
  or (_14427_, _14426_, _14424_);
  nor (_14428_, _14124_, _14108_);
  not (_14429_, _14428_);
  nor (_14430_, _14125_, _35638_);
  and (_14431_, _14430_, _14429_);
  not (_14432_, _14431_);
  and (_14433_, _13703_, _13701_);
  not (_14434_, _14433_);
  and (_14435_, _14434_, _13704_);
  and (_14436_, _14435_, _13534_);
  not (_14437_, _14436_);
  and (_14438_, _14156_, _33734_);
  and (_14439_, _14365_, _35601_);
  and (_14440_, _14439_, _33888_);
  nor (_14441_, _14440_, _14438_);
  nor (_14442_, _14441_, _34035_);
  not (_14443_, _14442_);
  and (_14444_, _14441_, _34035_);
  nor (_14445_, _14444_, _34100_);
  and (_14446_, _14445_, _14443_);
  and (_14447_, _35623_, _33935_);
  nor (_14448_, _34006_, _33814_);
  and (_14449_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_14450_, _14449_, _14448_);
  or (_14451_, _14450_, _35709_);
  nor (_14452_, _14451_, _14447_);
  not (_14453_, _14452_);
  nor (_14454_, _14453_, _14446_);
  and (_14455_, _14454_, _14437_);
  and (_14456_, _14455_, _14432_);
  nand (_14457_, _14456_, _14101_);
  and (_14458_, _14457_, _38997_);
  and (_38993_[3], _14458_, _14427_);
  nand (_14459_, _14043_, _14041_);
  or (_14460_, _14043_, _14041_);
  and (_14461_, _14460_, _14459_);
  and (_14462_, _14461_, _14055_);
  and (_14463_, _14057_, _13996_);
  or (_14464_, _14463_, _14462_);
  nand (_14465_, _14464_, _13774_);
  nand (_14466_, _13755_, _13534_);
  nor (_14467_, _35628_, _33991_);
  and (_14468_, _35628_, _33991_);
  nor (_14469_, _14468_, _14467_);
  and (_14470_, _14469_, _35582_);
  not (_14471_, _14470_);
  not (_14472_, _35659_);
  nor (_14473_, _35658_, _33991_);
  nor (_14474_, _14473_, _35638_);
  and (_14475_, _14474_, _14472_);
  nor (_14476_, _35691_, _33884_);
  not (_14477_, _14476_);
  nor (_14478_, _35692_, _35696_);
  and (_14479_, _14478_, _14477_);
  and (_14480_, _33935_, _33884_);
  not (_14481_, _14480_);
  or (_14482_, _34213_, _33797_);
  not (_14483_, _34020_);
  and (_14484_, _14483_, _14482_);
  and (_14485_, _14484_, _14481_);
  and (_14486_, _14485_, _33993_);
  not (_14487_, _14486_);
  nor (_14488_, _14487_, _14479_);
  and (_14489_, _14488_, _34016_);
  not (_14490_, _14489_);
  nor (_14491_, _14490_, _14475_);
  and (_14492_, _14491_, _14471_);
  and (_14493_, _14492_, _14466_);
  nand (_14494_, _14493_, _14465_);
  not (_14495_, _14494_);
  nor (_14496_, _14495_, _13836_);
  and (_14497_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_14498_, _14497_, _14101_);
  or (_14499_, _14498_, _14496_);
  nor (_14500_, _14129_, _14125_);
  nor (_14501_, _14500_, _14130_);
  and (_14502_, _14501_, _35637_);
  not (_14503_, _14502_);
  and (_14504_, _13707_, _13705_);
  not (_14505_, _14504_);
  and (_14506_, _14505_, _13708_);
  and (_14507_, _14506_, _13534_);
  and (_14508_, _14161_, _33888_);
  nor (_14509_, _14508_, _14158_);
  and (_14510_, _14509_, _33987_);
  nor (_14511_, _14509_, _33987_);
  nor (_14512_, _14511_, _14510_);
  and (_14513_, _14512_, _33899_);
  nor (_14514_, _33884_, _33734_);
  not (_14515_, _14514_);
  nor (_14516_, _14166_, _34006_);
  and (_14517_, _14516_, _14515_);
  and (_14518_, _34007_, _33935_);
  and (_14519_, _35708_, _35711_);
  and (_14520_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_14521_, _14520_, _14519_);
  nor (_14522_, _14521_, _14518_);
  not (_14523_, _14522_);
  nor (_14524_, _14523_, _14517_);
  not (_14525_, _14524_);
  nor (_14526_, _14525_, _14513_);
  not (_14527_, _14526_);
  nor (_14528_, _14527_, _14507_);
  and (_14529_, _14528_, _14503_);
  nand (_14530_, _14529_, _14101_);
  and (_14531_, _14530_, _38997_);
  and (_38993_[4], _14531_, _14499_);
  nand (_14532_, _14057_, _13989_);
  and (_14533_, _14459_, _13998_);
  nand (_14534_, _14533_, _14044_);
  or (_14535_, _14533_, _14044_);
  nand (_14536_, _14535_, _14534_);
  nand (_14537_, _14536_, _14055_);
  nand (_14538_, _14537_, _14532_);
  nand (_14539_, _14538_, _13774_);
  nand (_14540_, _13738_, _13534_);
  nor (_14541_, _35629_, _35599_);
  nor (_14542_, _14541_, _35630_);
  nor (_14543_, _14542_, _35583_);
  not (_14544_, _14543_);
  nor (_14545_, _33990_, _33967_);
  or (_14546_, _14545_, _35662_);
  and (_14547_, _14546_, _14472_);
  or (_14548_, _14547_, _35638_);
  nor (_14549_, _14548_, _35660_);
  nor (_14550_, _14068_, _35692_);
  and (_14551_, _14550_, _33797_);
  nor (_14552_, _14550_, _33797_);
  nor (_14553_, _14552_, _14551_);
  nor (_14554_, _14553_, _35696_);
  and (_14555_, _33935_, _33798_);
  not (_14556_, _14555_);
  or (_14557_, _34213_, _33765_);
  not (_14558_, _33994_);
  and (_14559_, _14558_, _14557_);
  and (_14560_, _14559_, _14556_);
  and (_14561_, _14560_, _33972_);
  and (_14562_, _14561_, _33969_);
  not (_14563_, _14562_);
  nor (_14564_, _14563_, _14554_);
  and (_14565_, _14564_, _33963_);
  not (_14566_, _14565_);
  nor (_14567_, _14566_, _14549_);
  and (_14568_, _14567_, _14544_);
  and (_14569_, _14568_, _14540_);
  and (_14570_, _14569_, _14539_);
  nor (_14571_, _14570_, _13836_);
  and (_14572_, _13836_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_14573_, _14572_, _14101_);
  or (_14574_, _14573_, _14571_);
  nor (_14575_, _14134_, _14130_);
  nor (_14576_, _14575_, _14135_);
  and (_14577_, _14576_, _35637_);
  not (_14578_, _14577_);
  and (_14579_, _13709_, _13687_);
  not (_14580_, _14579_);
  and (_14581_, _14580_, _13710_);
  and (_14582_, _14581_, _13534_);
  nor (_14583_, _14162_, _14158_);
  nor (_14584_, _14583_, _14166_);
  and (_14585_, _14584_, _33951_);
  nor (_14586_, _14584_, _33951_);
  or (_14587_, _14586_, _14585_);
  and (_14588_, _14587_, _33899_);
  and (_14589_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_14590_, _33798_, _33734_);
  or (_14591_, _14590_, _34006_);
  nor (_14592_, _14591_, _14165_);
  and (_14593_, _35708_, _13593_);
  and (_14594_, _35587_, _33935_);
  or (_14595_, _14594_, _14593_);
  or (_14596_, _14595_, _14592_);
  nor (_14597_, _14596_, _14589_);
  not (_14598_, _14597_);
  nor (_14599_, _14598_, _14588_);
  not (_14600_, _14599_);
  nor (_14601_, _14600_, _14582_);
  and (_14602_, _14601_, _14578_);
  nand (_14603_, _14602_, _14101_);
  and (_14604_, _14603_, _38997_);
  and (_38993_[5], _14604_, _14574_);
  or (_14605_, _14047_, _13981_);
  and (_14606_, _14605_, _14048_);
  or (_14607_, _14606_, _14057_);
  or (_14608_, _14055_, _13978_);
  and (_14609_, _14608_, _14607_);
  and (_14610_, _14609_, _13774_);
  and (_14611_, _13735_, _13534_);
  or (_14612_, _35666_, _35660_);
  nor (_14613_, _35667_, _35638_);
  and (_14614_, _14613_, _14612_);
  nor (_14615_, _35630_, _35596_);
  nor (_14616_, _14615_, _35631_);
  nor (_14617_, _14616_, _35583_);
  nor (_14618_, _14551_, _33765_);
  and (_14619_, _14551_, _33765_);
  or (_14620_, _14619_, _14618_);
  and (_14621_, _14620_, _35688_);
  and (_14622_, _33935_, _33766_);
  or (_14623_, _33973_, _34214_);
  nor (_14624_, _14623_, _14622_);
  and (_14625_, _14624_, _33926_);
  nand (_14626_, _14625_, _33918_);
  nor (_14627_, _14626_, _14621_);
  nand (_14628_, _14627_, _33903_);
  or (_14629_, _14628_, _14617_);
  or (_14630_, _14629_, _14614_);
  or (_14631_, _14630_, _14611_);
  or (_14632_, _14631_, _14610_);
  or (_14633_, _14632_, _13836_);
  not (_14634_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand (_14635_, _13836_, _14634_);
  and (_14636_, _14635_, _14633_);
  or (_14637_, _14636_, _14101_);
  or (_14638_, _14139_, _14135_);
  and (_14639_, _14638_, _14140_);
  and (_14640_, _14639_, _35637_);
  or (_14641_, _13711_, _13681_);
  and (_14642_, _14641_, _13712_);
  and (_14643_, _14642_, _13534_);
  and (_14644_, _14168_, _33778_);
  nor (_14645_, _14168_, _33778_);
  or (_14646_, _14645_, _14644_);
  and (_14647_, _14646_, _33899_);
  or (_14648_, _33766_, _33734_);
  nor (_14649_, _14169_, _34006_);
  and (_14650_, _14649_, _14648_);
  and (_14651_, _35708_, _33865_);
  and (_14652_, _35585_, _33935_);
  and (_14653_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_14654_, _14653_, _14652_);
  or (_14655_, _14654_, _14651_);
  or (_14656_, _14655_, _14650_);
  or (_14657_, _14656_, _14647_);
  or (_14658_, _14657_, _14643_);
  or (_14659_, _14658_, _14640_);
  or (_14660_, _14659_, _14229_);
  and (_14661_, _14660_, _38997_);
  and (_38993_[6], _14661_, _14637_);
  or (_14662_, _14223_, _14193_);
  or (_14663_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_14664_, _14663_, _38997_);
  and (_38994_[0], _14664_, _14662_);
  or (_14665_, _14289_, _14193_);
  or (_14666_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_14667_, _14666_, _38997_);
  and (_38994_[1], _14667_, _14665_);
  nand (_14668_, _14356_, _14194_);
  or (_14669_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_14670_, _14669_, _38997_);
  and (_38994_[2], _14670_, _14668_);
  nand (_14671_, _14423_, _14194_);
  or (_14672_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_14673_, _14672_, _38997_);
  and (_38994_[3], _14673_, _14671_);
  or (_14674_, _14494_, _14193_);
  or (_14675_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_14676_, _14675_, _38997_);
  and (_38994_[4], _14676_, _14674_);
  nand (_14677_, _14570_, _14194_);
  or (_14678_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_14679_, _14678_, _38997_);
  and (_38994_[5], _14679_, _14677_);
  or (_14680_, _14632_, _14193_);
  or (_14681_, _14194_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_14682_, _14681_, _38997_);
  and (_38994_[6], _14682_, _14680_);
  and (_36923_, _33533_, _38997_);
  and (_39017_, _36923_, _33475_);
  and (_39018_[7], _34223_, _38997_);
  nand (_39018_[0], _34466_, _38997_);
  nand (_39018_[1], _34557_, _38997_);
  nand (_39018_[2], _34766_, _38997_);
  and (_39018_[3], _34401_, _38997_);
  and (_39018_[4], _34525_, _38997_);
  nor (_39018_[5], _34615_, rst);
  nor (_39018_[6], _34649_, rst);
  not (_14683_, _14098_);
  nand (_14684_, _13158_, _34231_);
  or (_14685_, _14684_, _14683_);
  not (_14686_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_14687_, _14684_, _14686_);
  and (_14688_, _14687_, _33662_);
  and (_14689_, _14688_, _14685_);
  nor (_14690_, _33661_, _14686_);
  nor (_14691_, _33630_, _33591_);
  and (_14692_, _14691_, _13123_);
  and (_14693_, _14692_, _11075_);
  nand (_14694_, _14693_, _35722_);
  or (_14695_, _14693_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_14696_, _14695_, _11083_);
  and (_14697_, _14696_, _14694_);
  or (_14698_, _14697_, _14690_);
  or (_14699_, _14698_, _14689_);
  and (_38992_[7], _14699_, _38997_);
  or (_14700_, _14684_, _14223_);
  not (_14701_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_14702_, _14684_, _14701_);
  and (_14703_, _14702_, _33662_);
  and (_14704_, _14703_, _14700_);
  nor (_14705_, _33661_, _14701_);
  or (_14706_, _14684_, _35723_);
  and (_14707_, _14702_, _11083_);
  and (_14708_, _14707_, _14706_);
  or (_14709_, _14708_, _14705_);
  or (_14710_, _14709_, _14704_);
  and (_38992_[0], _14710_, _38997_);
  or (_14711_, _14684_, _14289_);
  not (_14712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_14713_, _14684_, _14712_);
  and (_14714_, _14713_, _33662_);
  and (_14715_, _14714_, _14711_);
  nor (_14716_, _33661_, _14712_);
  and (_14717_, _14692_, _34253_);
  nand (_14718_, _14717_, _35722_);
  or (_14719_, _14717_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_14720_, _14719_, _11083_);
  and (_14721_, _14720_, _14718_);
  or (_14722_, _14721_, _14716_);
  or (_14723_, _14722_, _14715_);
  and (_38992_[1], _14723_, _38997_);
  not (_14724_, _14356_);
  or (_14725_, _14684_, _14724_);
  not (_14726_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_14727_, _14684_, _14726_);
  and (_14728_, _14727_, _33662_);
  and (_14729_, _14728_, _14725_);
  nor (_14730_, _33661_, _14726_);
  nand (_14731_, _14692_, _11359_);
  and (_14732_, _14731_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_14733_, _34252_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_14734_, _14733_, _11345_);
  and (_14735_, _14734_, _14692_);
  or (_14736_, _14735_, _14732_);
  and (_14737_, _14736_, _11083_);
  or (_14738_, _14737_, _14730_);
  or (_14739_, _14738_, _14729_);
  and (_38992_[2], _14739_, _38997_);
  not (_14740_, _14423_);
  or (_14741_, _14684_, _14740_);
  not (_14742_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_14743_, _14684_, _14742_);
  and (_14744_, _14743_, _33662_);
  and (_14745_, _14744_, _14741_);
  nor (_14746_, _33661_, _14742_);
  and (_14747_, _14692_, _11356_);
  nand (_14748_, _14747_, _35722_);
  or (_14749_, _14747_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_14750_, _14749_, _11083_);
  and (_14751_, _14750_, _14748_);
  or (_14752_, _14751_, _14746_);
  or (_14753_, _14752_, _14745_);
  and (_38992_[3], _14753_, _38997_);
  or (_14754_, _14684_, _14494_);
  not (_14755_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_14756_, _14684_, _14755_);
  and (_14757_, _14756_, _33662_);
  and (_14758_, _14757_, _14754_);
  nor (_14759_, _33661_, _14755_);
  and (_14760_, _14692_, _11370_);
  nand (_14761_, _14760_, _35722_);
  or (_14762_, _14760_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_14763_, _14762_, _11083_);
  and (_14764_, _14763_, _14761_);
  or (_14765_, _14764_, _14759_);
  or (_14766_, _14765_, _14758_);
  and (_38992_[4], _14766_, _38997_);
  not (_14767_, _14570_);
  or (_14768_, _14684_, _14767_);
  not (_14769_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_14770_, _14684_, _14769_);
  and (_14771_, _14770_, _33662_);
  and (_14772_, _14771_, _14768_);
  nor (_14773_, _33661_, _14769_);
  and (_14774_, _14692_, _11383_);
  nand (_14775_, _14774_, _35722_);
  or (_14776_, _14774_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_14777_, _14776_, _11083_);
  and (_14778_, _14777_, _14775_);
  or (_14779_, _14778_, _14773_);
  or (_14780_, _14779_, _14772_);
  and (_38992_[5], _14780_, _38997_);
  or (_14781_, _14684_, _14632_);
  not (_14782_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_14783_, _14684_, _14782_);
  and (_14784_, _14783_, _33662_);
  and (_14785_, _14784_, _14781_);
  nor (_14786_, _33661_, _14782_);
  nand (_14787_, _14692_, _11392_);
  or (_14788_, _14787_, _35723_);
  nand (_14789_, _14787_, _14782_);
  and (_14790_, _14789_, _11083_);
  and (_14791_, _14790_, _14788_);
  or (_14792_, _14791_, _14786_);
  or (_14793_, _14792_, _14785_);
  and (_38992_[6], _14793_, _38997_);
  nor (_14794_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_14795_, _14794_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_14796_, _12066_, _34231_);
  and (_14797_, _14796_, _34257_);
  and (_14798_, _14797_, _33662_);
  nor (_14799_, _14798_, _14795_);
  or (_14800_, _14799_, _14098_);
  not (_14801_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_14802_, _14100_, _14801_);
  not (_14803_, _14802_);
  and (_14804_, _14691_, _11083_);
  and (_14805_, _14804_, _13106_);
  and (_14806_, _14805_, _11075_);
  and (_14807_, _14806_, _35722_);
  nor (_14808_, _14806_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_14809_, _14808_);
  nand (_14810_, _14809_, _14799_);
  or (_14811_, _14810_, _14807_);
  and (_14812_, _14811_, _14803_);
  and (_14813_, _14812_, _14800_);
  and (_14814_, _14802_, _14189_);
  or (_14815_, _14814_, _14813_);
  nor (_38991_[7], _14815_, rst);
  or (_14816_, _14799_, _14223_);
  nor (_14817_, _34229_, _34128_);
  nor (_14818_, _14817_, _11315_);
  or (_14819_, _14802_, _14795_);
  nor (_14820_, _14819_, _14798_);
  and (_14821_, _14820_, _14805_);
  not (_14822_, _14821_);
  nor (_14823_, _14822_, _14818_);
  not (_14824_, _14799_);
  nor (_14825_, _14805_, _34128_);
  nor (_14826_, _14825_, _14824_);
  not (_14827_, _14826_);
  nor (_14828_, _14827_, _14823_);
  nor (_14829_, _14828_, _14802_);
  nand (_14830_, _14829_, _14816_);
  nand (_14831_, _14802_, _14250_);
  nand (_14832_, _14831_, _14830_);
  and (_38991_[0], _14832_, _38997_);
  nor (_14833_, _14803_, _14323_);
  not (_14834_, _14833_);
  or (_14835_, _14799_, _14289_);
  not (_14836_, _14805_);
  nor (_14837_, _34253_, _34095_);
  nor (_14838_, _14837_, _11326_);
  nor (_14839_, _14838_, _14836_);
  nor (_14840_, _14805_, _34095_);
  nor (_14841_, _14840_, _14824_);
  not (_14842_, _14841_);
  nor (_14843_, _14842_, _14839_);
  nor (_14844_, _14843_, _14802_);
  nand (_14845_, _14844_, _14835_);
  nand (_14846_, _14845_, _14834_);
  and (_38991_[1], _14846_, _38997_);
  or (_14847_, _14799_, _14356_);
  and (_14848_, _14805_, _11343_);
  and (_14849_, _14848_, _35722_);
  nor (_14850_, _14848_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_14851_, _14850_);
  nand (_14852_, _14851_, _14799_);
  or (_14853_, _14852_, _14849_);
  and (_14854_, _14853_, _14803_);
  nand (_14855_, _14854_, _14847_);
  and (_14856_, _14802_, _14387_);
  not (_14857_, _14856_);
  and (_14858_, _14857_, _14855_);
  and (_38991_[2], _14858_, _38997_);
  or (_14859_, _14799_, _14423_);
  and (_14860_, _14821_, _11357_);
  and (_14861_, _14805_, _11356_);
  nand (_14862_, _14799_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_14863_, _14862_, _14861_);
  or (_14864_, _14863_, _14802_);
  nor (_14865_, _14864_, _14860_);
  nand (_14866_, _14865_, _14859_);
  and (_14867_, _14802_, _14456_);
  not (_14868_, _14867_);
  and (_14869_, _14868_, _14866_);
  and (_38991_[3], _14869_, _38997_);
  nor (_14870_, _14803_, _14529_);
  not (_14871_, _14870_);
  or (_14872_, _14799_, _14494_);
  nor (_14873_, _11370_, _33984_);
  nor (_14874_, _14873_, _11376_);
  nor (_14875_, _14874_, _14822_);
  nor (_14876_, _14805_, _33984_);
  nor (_14877_, _14876_, _14824_);
  not (_14878_, _14877_);
  nor (_14879_, _14878_, _14875_);
  nor (_14880_, _14879_, _14802_);
  nand (_14881_, _14880_, _14872_);
  nand (_14882_, _14881_, _14871_);
  and (_38991_[4], _14882_, _38997_);
  or (_14883_, _14799_, _14570_);
  nand (_14884_, _14821_, _11383_);
  or (_14885_, _14884_, _35722_);
  and (_14886_, _14805_, _11383_);
  nand (_14887_, _14799_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_14888_, _14887_, _14886_);
  and (_14889_, _14888_, _14803_);
  and (_14890_, _14889_, _14885_);
  nand (_14891_, _14890_, _14883_);
  and (_14892_, _14802_, _14602_);
  not (_14893_, _14892_);
  and (_14894_, _14893_, _14891_);
  and (_38991_[5], _14894_, _38997_);
  and (_14895_, _14824_, _14632_);
  and (_14896_, _14821_, _12080_);
  nand (_14897_, _14805_, _11392_);
  and (_14898_, _14799_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_14899_, _14898_, _14897_);
  or (_14900_, _14899_, _14802_);
  or (_14901_, _14900_, _14896_);
  or (_14902_, _14901_, _14895_);
  or (_14903_, _14803_, _14659_);
  and (_14904_, _14903_, _14902_);
  and (_38991_[6], _14904_, _38997_);
  and (_14905_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_14906_, _14905_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_14907_, _14905_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_14908_, _14907_, _14906_);
  and (_36859_[1], _14908_, _38997_);
  and (_36860_[5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _38997_);
  nor (_36861_[7], _14064_, rst);
  and (_36860_[0], _14055_, _38997_);
  and (_36860_[1], _13957_, _38997_);
  and (_36860_[2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _38997_);
  and (_36860_[3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _38997_);
  and (_36860_[4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _38997_);
  or (_14909_, _13774_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_14910_, _14905_, rst);
  and (_36859_[0], _14910_, _14909_);
  and (_36861_[0], _14202_, _38997_);
  and (_36861_[1], _14259_, _38997_);
  and (_36861_[2], _14332_, _38997_);
  and (_36861_[3], _14398_, _38997_);
  and (_36861_[4], _14464_, _38997_);
  and (_36861_[5], _14538_, _38997_);
  and (_36861_[6], _14609_, _38997_);
  nand (_14911_, _13548_, _13534_);
  or (_14912_, _13534_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_14913_, _14912_, _38997_);
  and (_36862_[1], _14913_, _14911_);
  nor (_36863_[15], _13732_, rst);
  nor (_14914_, _13534_, _13543_);
  and (_14915_, _13534_, _13543_);
  or (_14916_, _14915_, _14914_);
  and (_36862_[0], _14916_, _38997_);
  and (_36863_[0], _13621_, _38997_);
  and (_36863_[1], _14313_, _38997_);
  and (_36863_[2], _14374_, _38997_);
  and (_36863_[3], _14435_, _38997_);
  and (_36863_[4], _14506_, _38997_);
  and (_36863_[5], _14581_, _38997_);
  and (_36863_[6], _14642_, _38997_);
  and (_36863_[7], _14151_, _38997_);
  and (_36863_[8], _13743_, _38997_);
  and (_36863_[9], _13747_, _38997_);
  and (_36863_[10], _13752_, _38997_);
  and (_36863_[11], _13784_, _38997_);
  and (_36863_[12], _13755_, _38997_);
  and (_36863_[13], _13738_, _38997_);
  and (_36863_[14], _13735_, _38997_);
  nor (_36867_[2], _33497_, rst);
  and (_14917_, _33387_, _33410_);
  and (_14918_, _33371_, _33252_);
  nor (_14919_, _14918_, _14917_);
  and (_14920_, _33371_, _33385_);
  not (_14921_, _14920_);
  and (_14922_, _14921_, _14919_);
  and (_14923_, _33135_, _38997_);
  not (_14924_, _14923_);
  or (_14925_, _14924_, _14917_);
  or (_36868_[2], _14925_, _14922_);
  and (_14926_, _33197_, _33172_);
  not (_14927_, _33222_);
  nor (_14928_, _33246_, _14927_);
  and (_14929_, _14928_, _14926_);
  not (_14930_, _33295_);
  not (_14931_, _33319_);
  and (_14932_, _33344_, _14931_);
  and (_14933_, _14932_, _14930_);
  and (_14934_, _14933_, _14929_);
  not (_14935_, _33271_);
  nor (_14936_, _33197_, _14935_);
  and (_14937_, _14932_, _33295_);
  and (_14938_, _14937_, _14936_);
  not (_14939_, _33246_);
  not (_14940_, _33172_);
  and (_14941_, _33197_, _14940_);
  and (_14942_, _14941_, _14939_);
  nor (_14943_, _33344_, _33319_);
  nor (_14944_, _33295_, _14935_);
  and (_14945_, _14944_, _14943_);
  and (_14946_, _14945_, _14942_);
  or (_14947_, _14946_, _14938_);
  nor (_14948_, _14947_, _14934_);
  and (_14949_, _14943_, _14930_);
  and (_14950_, _33246_, _33271_);
  and (_14951_, _14950_, _14941_);
  or (_14952_, _14951_, _14936_);
  and (_14953_, _14952_, _14949_);
  and (_14954_, _33344_, _33319_);
  and (_14955_, _14954_, _33271_);
  and (_14956_, _14955_, _14929_);
  nor (_14957_, _14956_, _14953_);
  nand (_14958_, _14957_, _14948_);
  and (_14959_, _14941_, _14928_);
  and (_14960_, _14959_, _14935_);
  and (_14961_, _14960_, _14943_);
  and (_14962_, _33295_, _14935_);
  and (_14963_, _14962_, _14943_);
  and (_14964_, _14963_, _14929_);
  and (_14965_, _14926_, _33246_);
  and (_14966_, _14965_, _33222_);
  nor (_14967_, _33344_, _14931_);
  and (_14968_, _14967_, _33295_);
  and (_14969_, _14968_, _14966_);
  nor (_14970_, _14969_, _14964_);
  not (_14971_, _14970_);
  or (_14972_, _14971_, _14961_);
  or (_14973_, _14972_, _14958_);
  and (_14974_, _33295_, _33271_);
  and (_14975_, _14967_, _14974_);
  nor (_14976_, _33295_, _33271_);
  and (_14977_, _14967_, _14976_);
  or (_14978_, _14977_, _14975_);
  and (_14979_, _14978_, _14929_);
  and (_14980_, _14974_, _14932_);
  and (_14981_, _14942_, _14927_);
  and (_14982_, _14981_, _14980_);
  nor (_14983_, _14982_, _14979_);
  and (_14984_, _14926_, _14939_);
  not (_14985_, _14984_);
  and (_14986_, _14976_, _14954_);
  nor (_14987_, _14986_, _14927_);
  nor (_14988_, _14987_, _14985_);
  not (_14989_, _14988_);
  and (_14990_, _14962_, _14954_);
  and (_14991_, _14990_, _14929_);
  and (_14992_, _14967_, _14944_);
  and (_14993_, _14992_, _14929_);
  nor (_14994_, _14993_, _14991_);
  and (_14995_, _14994_, _14989_);
  and (_14996_, _14954_, _14944_);
  and (_14997_, _14965_, _14927_);
  and (_14998_, _14997_, _14996_);
  and (_14999_, _14967_, _14930_);
  and (_15000_, _14999_, _14966_);
  or (_15001_, _15000_, _14998_);
  and (_15002_, _14943_, _33295_);
  and (_15003_, _14997_, _15002_);
  and (_15004_, _14965_, _14933_);
  or (_15005_, _15004_, _15003_);
  nor (_15006_, _15005_, _15001_);
  and (_15007_, _15006_, _14995_);
  nand (_15008_, _15007_, _14983_);
  or (_15009_, _15008_, _14973_);
  and (_15010_, _15009_, _33136_);
  not (_15011_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_15012_, _33134_, _33129_);
  and (_15013_, _15012_, _33456_);
  nor (_15014_, _15013_, _15011_);
  or (_15015_, _15014_, rst);
  or (_36869_[1], _15015_, _15010_);
  nand (_15016_, _33319_, _33130_);
  or (_15017_, _33130_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_15018_, _15017_, _38997_);
  and (_36870_[7], _15018_, _15016_);
  and (_15019_, \oc8051_top_1.oc8051_sfr1.wait_data , _38997_);
  and (_15020_, _15019_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_15021_, _33252_, _33381_);
  nor (_15022_, _15021_, _33459_);
  and (_15023_, _33423_, _33410_);
  nor (_15024_, _15023_, _34354_);
  nand (_15025_, _15024_, _15022_);
  and (_15026_, _33388_, _33410_);
  and (_15027_, _33478_, _33372_);
  or (_15028_, _15027_, _15026_);
  and (_15029_, _33388_, _33252_);
  nor (_15030_, _15029_, _34349_);
  nand (_15031_, _15030_, _33362_);
  or (_15032_, _15031_, _15028_);
  or (_15033_, _15032_, _15025_);
  and (_15034_, _15033_, _14923_);
  or (_36871_, _15034_, _15020_);
  not (_15035_, _33485_);
  and (_15036_, _33437_, _33252_);
  or (_15037_, _15036_, _15035_);
  and (_15038_, _33443_, _33417_);
  or (_15039_, _15038_, _33521_);
  and (_15040_, _33365_, _33366_);
  and (_15041_, _15040_, _33423_);
  or (_15042_, _15041_, _15039_);
  or (_15043_, _15042_, _15037_);
  and (_15044_, _15043_, _33135_);
  and (_15045_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15046_, _33467_, _15011_);
  not (_15047_, _33481_);
  and (_15048_, _15047_, _15046_);
  or (_15049_, _15048_, _15045_);
  or (_15050_, _15049_, _15044_);
  and (_36872_[1], _15050_, _38997_);
  and (_15051_, _15019_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15052_, _33478_, _33395_);
  or (_15053_, _33395_, _33418_);
  and (_15054_, _15053_, _33368_);
  or (_15055_, _15054_, _15052_);
  and (_15056_, _15040_, _33359_);
  or (_15057_, _15056_, _15055_);
  and (_15058_, _15053_, _33201_);
  and (_15059_, _33201_, _33275_);
  and (_15060_, _15059_, _33358_);
  or (_15061_, _15060_, _15058_);
  and (_15062_, _15059_, _33375_);
  nor (_15063_, _15062_, _33504_);
  not (_15064_, _15063_);
  and (_15065_, _33374_, _33275_);
  and (_15066_, _33478_, _15065_);
  or (_15067_, _15066_, _33506_);
  or (_15068_, _15067_, _15064_);
  or (_15069_, _15068_, _15037_);
  or (_15070_, _15069_, _15061_);
  or (_15071_, _15070_, _15057_);
  and (_15072_, _15071_, _14923_);
  or (_36873_[1], _15072_, _15051_);
  and (_15073_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15074_, _33436_, _33135_);
  or (_15075_, _15074_, _15073_);
  or (_15076_, _15075_, _15048_);
  and (_36874_[2], _15076_, _38997_);
  and (_15077_, _33367_, _33202_);
  and (_15078_, _33391_, _33358_);
  nor (_15079_, _15078_, _15077_);
  nor (_15080_, _15079_, _33354_);
  and (_15081_, _15026_, _33131_);
  nor (_15082_, _15081_, _15080_);
  nor (_15083_, _15082_, _33467_);
  nor (_15084_, _14917_, _33354_);
  nor (_15085_, _15084_, _14922_);
  and (_15086_, _15085_, _15046_);
  or (_15087_, _15086_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15088_, _15087_, _15083_);
  or (_15089_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _33129_);
  and (_15090_, _15089_, _38997_);
  and (_36875_[2], _15090_, _15088_);
  and (_15091_, _15019_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_15092_, _15060_, _15035_);
  and (_15093_, _33418_, _33201_);
  or (_15094_, _15093_, _33419_);
  or (_15095_, _15094_, _15092_);
  or (_15096_, _34356_, _34354_);
  or (_15097_, _15096_, _33434_);
  or (_15098_, _33359_, _33423_);
  and (_15099_, _15098_, _33398_);
  or (_15100_, _15056_, _15038_);
  or (_15101_, _15100_, _34348_);
  or (_15102_, _15101_, _15099_);
  or (_15103_, _15102_, _15097_);
  or (_15104_, _15103_, _15095_);
  and (_15105_, _15104_, _14923_);
  or (_36876_[1], _15105_, _15091_);
  and (_15106_, _15019_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_15107_, _33398_, _33418_);
  not (_15108_, _33511_);
  and (_15109_, _33515_, _33380_);
  or (_15110_, _15109_, _15108_);
  or (_15111_, _15110_, _15107_);
  and (_15112_, _15040_, _33429_);
  and (_15113_, _33349_, _33410_);
  or (_15114_, _15113_, _15041_);
  or (_15115_, _15114_, _15112_);
  or (_15116_, _15115_, _15061_);
  or (_15117_, _15116_, _15111_);
  and (_15118_, _33403_, _33465_);
  or (_15119_, _15118_, _33411_);
  or (_15120_, _15119_, _34359_);
  and (_15121_, _33478_, _33403_);
  or (_15122_, _15121_, _15120_);
  and (_15123_, _33443_, _33380_);
  and (_15124_, _33443_, _33407_);
  or (_15125_, _15124_, _15123_);
  or (_15126_, _33506_, _33430_);
  or (_15127_, _33416_, _33406_);
  or (_15128_, _15127_, _15126_);
  or (_15129_, _15128_, _15125_);
  or (_15130_, _15129_, _15057_);
  or (_15131_, _15130_, _15122_);
  or (_15132_, _15131_, _15117_);
  and (_15133_, _15132_, _14923_);
  or (_36877_[3], _15133_, _15106_);
  and (_15134_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_15135_, _33481_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15136_, _15135_, _15134_);
  and (_15137_, _15136_, _38997_);
  and (_15138_, _33398_, _33350_);
  and (_15139_, _15059_, _33387_);
  or (_15140_, _15139_, _15138_);
  and (_15141_, _15040_, _33350_);
  or (_15142_, _15141_, _15140_);
  and (_15143_, _15040_, _33437_);
  and (_15144_, _33350_, _33201_);
  or (_15145_, _15144_, _33522_);
  or (_15146_, _15145_, _15143_);
  or (_15147_, _15146_, _15142_);
  and (_15148_, _15147_, _14923_);
  or (_36878_[1], _15148_, _15137_);
  or (_15149_, _34351_, _33436_);
  or (_15150_, _15149_, _34350_);
  or (_15151_, _15054_, _33432_);
  or (_15152_, _15151_, _15150_);
  or (_15153_, _34355_, _33434_);
  and (_15154_, _33359_, _33465_);
  and (_15155_, _33370_, _33275_);
  and (_15156_, _15155_, _33368_);
  or (_15157_, _15156_, _33420_);
  or (_15158_, _15157_, _15154_);
  or (_15159_, _15158_, _15119_);
  or (_15160_, _15159_, _15153_);
  or (_15161_, _15160_, _15152_);
  and (_15162_, _33397_, _33201_);
  and (_15163_, _15059_, _33370_);
  or (_15164_, _15163_, _15162_);
  or (_15165_, _15164_, _15039_);
  or (_15166_, _15165_, _15061_);
  and (_15167_, _33398_, _33275_);
  and (_15168_, _15167_, _33370_);
  or (_15169_, _15168_, _33506_);
  or (_15170_, _15169_, _33399_);
  and (_15171_, _33388_, _33201_);
  and (_15172_, _15077_, _33275_);
  or (_15173_, _15172_, _33507_);
  or (_15174_, _15173_, _15171_);
  or (_15175_, _15174_, _33386_);
  or (_15176_, _15175_, _15170_);
  or (_15177_, _15176_, _15166_);
  or (_15178_, _15177_, _15161_);
  and (_15179_, _15178_, _33135_);
  and (_15180_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15181_, _33461_, _33359_);
  and (_15182_, _15080_, _33458_);
  or (_15183_, _15182_, _15048_);
  or (_15184_, _15183_, _15181_);
  or (_15185_, _15184_, _15180_);
  or (_15186_, _15185_, _15179_);
  and (_36879_, _15186_, _38997_);
  and (_36867_[0], _33530_, _38997_);
  and (_36867_[1], _33472_, _38997_);
  nand (_36868_[0], _15085_, _14923_);
  or (_36868_[1], _14924_, _14919_);
  or (_15187_, _15000_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_15188_, _15187_, _15003_);
  or (_15189_, _15188_, _14961_);
  and (_15190_, _15189_, _15013_);
  nor (_15191_, _15012_, _33456_);
  or (_15192_, _15191_, rst);
  or (_36869_[0], _15192_, _15190_);
  nand (_15193_, _33222_, _33130_);
  or (_15194_, _33130_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_15195_, _15194_, _38997_);
  and (_36870_[0], _15195_, _15193_);
  or (_15196_, _33246_, _33490_);
  or (_15197_, _33130_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_15198_, _15197_, _38997_);
  and (_36870_[1], _15198_, _15196_);
  nand (_15199_, _33172_, _33130_);
  or (_15200_, _33130_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_15201_, _15200_, _38997_);
  and (_36870_[2], _15201_, _15199_);
  nand (_15202_, _33197_, _33130_);
  or (_15203_, _33130_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_15204_, _15203_, _38997_);
  and (_36870_[3], _15204_, _15202_);
  or (_15205_, _33271_, _33490_);
  or (_15206_, _33130_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_15207_, _15206_, _38997_);
  and (_36870_[4], _15207_, _15205_);
  nand (_15208_, _33295_, _33130_);
  or (_15209_, _33130_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_15210_, _15209_, _38997_);
  and (_36870_[5], _15210_, _15208_);
  or (_15211_, _33344_, _33490_);
  or (_15212_, _33130_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_15213_, _15212_, _38997_);
  and (_36870_[6], _15213_, _15211_);
  and (_15214_, _15059_, _33381_);
  or (_15215_, _15214_, _15144_);
  or (_15216_, _15215_, _15143_);
  or (_15217_, _33359_, _33418_);
  and (_15218_, _15217_, _33478_);
  or (_15219_, _15218_, _15052_);
  and (_15220_, _33478_, _33408_);
  and (_15221_, _33371_, _33275_);
  and (_15222_, _15221_, _33478_);
  and (_15223_, _15040_, _33382_);
  or (_15224_, _15223_, _15222_);
  or (_15225_, _15224_, _15220_);
  or (_15226_, _15225_, _15219_);
  or (_15227_, _15226_, _15216_);
  and (_15228_, _15040_, _33403_);
  or (_15229_, _15228_, _15036_);
  and (_15230_, _33443_, _33371_);
  and (_15231_, _33443_, _33381_);
  or (_15232_, _15231_, _33522_);
  or (_15233_, _15232_, _15230_);
  or (_15234_, _15233_, _15142_);
  or (_15235_, _15234_, _15229_);
  or (_15236_, _15124_, _15112_);
  and (_15237_, _15167_, _33381_);
  and (_15238_, _15040_, _33372_);
  or (_15239_, _15238_, _15237_);
  or (_15240_, _15239_, _15236_);
  nand (_15241_, _33511_, _33485_);
  not (_15242_, _33518_);
  or (_15243_, _15113_, _15242_);
  or (_15244_, _15243_, _15241_);
  or (_15245_, _15244_, _15240_);
  or (_15246_, _15245_, _15235_);
  or (_15247_, _15246_, _15227_);
  and (_15248_, _15247_, _33135_);
  and (_15249_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15250_, _15249_, _15086_);
  or (_15251_, _15250_, _15248_);
  and (_36872_[0], _15251_, _38997_);
  and (_15252_, _15019_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_15253_, _15125_, _15028_);
  and (_15254_, _33478_, _33383_);
  or (_15255_, _15254_, _15229_);
  or (_15256_, _15255_, _15253_);
  and (_15257_, _33429_, _33465_);
  and (_15258_, _33478_, _33429_);
  or (_15259_, _15258_, _15064_);
  or (_15260_, _15259_, _15257_);
  or (_15261_, _15066_, _15118_);
  or (_15262_, _15261_, _33435_);
  or (_15263_, _15262_, _15260_);
  or (_15264_, _15263_, _15111_);
  or (_15265_, _15264_, _15256_);
  and (_15266_, _15265_, _14923_);
  or (_36873_[0], _15266_, _15252_);
  or (_15267_, _15175_, _15161_);
  and (_15268_, _15267_, _33135_);
  and (_15269_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15270_, _15269_, _15184_);
  or (_15271_, _15270_, _15268_);
  and (_36874_[0], _15271_, _38997_);
  and (_15272_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15273_, _15272_, _15183_);
  nand (_15274_, _33431_, _33354_);
  nand (_15275_, _15274_, _33520_);
  or (_15276_, _15275_, _15080_);
  or (_15277_, _15276_, _15170_);
  and (_15278_, _15277_, _33135_);
  or (_15279_, _15278_, _15273_);
  and (_36874_[1], _15279_, _38997_);
  or (_15280_, _14917_, _33480_);
  and (_15281_, _15141_, _33275_);
  or (_15282_, _15281_, _15223_);
  or (_15283_, _15282_, _15280_);
  or (_15284_, _15220_, _15258_);
  and (_15285_, _15221_, _33368_);
  and (_15286_, _15141_, _33354_);
  or (_15287_, _15286_, _15285_);
  or (_15288_, _15287_, _15284_);
  or (_15289_, _15288_, _15080_);
  or (_15290_, _15289_, _15283_);
  and (_15291_, _15040_, _33376_);
  or (_15292_, _15291_, _15027_);
  or (_15293_, _15222_, _33479_);
  or (_15294_, _15293_, _15292_);
  or (_15295_, _15294_, _15219_);
  and (_15296_, _33478_, _33423_);
  or (_15297_, _15113_, _15296_);
  or (_15298_, _15297_, _15216_);
  nor (_15299_, _15163_, _33522_);
  nand (_15300_, _15299_, _33484_);
  or (_15301_, _15168_, _15121_);
  or (_15302_, _15301_, _15300_);
  or (_15303_, _15140_, _15237_);
  and (_15304_, _33386_, _33464_);
  or (_15305_, _15304_, _15303_);
  or (_15306_, _15305_, _15302_);
  or (_15307_, _15306_, _15298_);
  or (_15308_, _15307_, _15295_);
  or (_15309_, _15308_, _15290_);
  and (_15310_, _15309_, _33135_);
  and (_15311_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_15312_, _33481_, _33131_);
  and (_15313_, _33372_, _33252_);
  or (_15314_, _15026_, _33482_);
  nor (_15315_, _33201_, _33275_);
  and (_15316_, _33371_, _33389_);
  and (_15317_, _15316_, _15315_);
  or (_15318_, _15317_, _15314_);
  or (_15319_, _15318_, _15313_);
  and (_15320_, _15319_, _15046_);
  or (_15321_, _15320_, _15312_);
  or (_15322_, _15321_, _15311_);
  or (_15323_, _15322_, _15310_);
  and (_36875_[0], _15323_, _38997_);
  and (_15324_, _15059_, _33371_);
  or (_15325_, _15156_, _15036_);
  or (_15326_, _15325_, _15324_);
  or (_15327_, _15326_, _33384_);
  or (_15328_, _15327_, _15303_);
  and (_15329_, _33429_, _33410_);
  and (_15330_, _15221_, _33398_);
  or (_15331_, _15330_, _33386_);
  or (_15332_, _15331_, _15329_);
  or (_15333_, _33522_, _33480_);
  or (_15334_, _15333_, _33482_);
  not (_15335_, _33484_);
  or (_15336_, _15335_, _33411_);
  or (_15337_, _15336_, _15334_);
  or (_15338_, _15337_, _15332_);
  or (_15339_, _15338_, _15328_);
  or (_15340_, _15298_, _15295_);
  or (_15341_, _15340_, _15339_);
  and (_15342_, _15341_, _33135_);
  and (_15343_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15344_, _15343_, _15321_);
  or (_15345_, _15344_, _15342_);
  and (_36875_[1], _15345_, _38997_);
  and (_15346_, _15019_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_15347_, _15095_, _34362_);
  or (_15348_, _15347_, _15153_);
  or (_15349_, _33410_, _33201_);
  and (_15350_, _15349_, _33351_);
  and (_15351_, _33478_, _33418_);
  and (_15352_, _33376_, _33410_);
  or (_15353_, _15352_, _15351_);
  and (_15354_, _15217_, _33410_);
  or (_15355_, _15354_, _15353_);
  or (_15356_, _15355_, _15350_);
  and (_15357_, _15167_, _33350_);
  or (_15358_, _15281_, _15357_);
  or (_15359_, _15139_, _15038_);
  or (_15360_, _15143_, _15056_);
  or (_15361_, _15360_, _15359_);
  or (_15362_, _15361_, _15358_);
  or (_15363_, _33522_, _34351_);
  or (_15364_, _15363_, _15099_);
  or (_15365_, _15364_, _15362_);
  or (_15366_, _15365_, _15356_);
  or (_15367_, _15366_, _15348_);
  and (_15368_, _15367_, _14923_);
  or (_36876_[0], _15368_, _15346_);
  or (_15369_, _15109_, _15041_);
  or (_15370_, _15286_, _15107_);
  or (_15371_, _15370_, _15369_);
  nor (_15372_, _15123_, _33404_);
  nand (_15373_, _15372_, _33486_);
  or (_15374_, _15373_, _15371_);
  and (_15375_, _33359_, _33410_);
  and (_15376_, _33351_, _33410_);
  or (_15377_, _15351_, _15376_);
  or (_15378_, _15377_, _15375_);
  or (_15379_, _15378_, _15283_);
  or (_15380_, _15379_, _15374_);
  nor (_15381_, _34358_, _33386_);
  not (_15382_, _15381_);
  or (_15383_, _33503_, _15382_);
  or (_15384_, _15383_, _15215_);
  or (_15385_, _15384_, _15122_);
  or (_15386_, _15385_, _15380_);
  and (_15387_, _15386_, _14923_);
  and (_15388_, _15019_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_15389_, _33492_, _38997_);
  or (_15390_, _15389_, _15388_);
  or (_36877_[0], _15390_, _15387_);
  and (_15391_, _33350_, _33410_);
  or (_15392_, _15391_, _15361_);
  or (_15393_, _33504_, _33405_);
  or (_15394_, _15393_, _15062_);
  not (_15395_, _33523_);
  or (_15396_, _15041_, _15395_);
  or (_15397_, _15396_, _15394_);
  or (_15398_, _15397_, _15392_);
  not (_15399_, _15223_);
  and (_15400_, _15399_, _15381_);
  not (_15401_, _15400_);
  or (_15402_, _15401_, _15055_);
  or (_15403_, _15402_, _15398_);
  or (_15404_, _15214_, _15061_);
  or (_15405_, _15222_, _34347_);
  or (_15406_, _15405_, _15292_);
  nor (_15407_, _33506_, _15237_);
  not (_15408_, _15407_);
  or (_15409_, _15408_, _15406_);
  or (_15410_, _15409_, _15404_);
  or (_15411_, _15410_, _15403_);
  and (_15412_, _15411_, _33135_);
  and (_15413_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15414_, _15413_, _33491_);
  or (_15415_, _15414_, _15412_);
  and (_36877_[1], _15415_, _38997_);
  and (_15416_, _33358_, _33410_);
  or (_15417_, _15039_, _33434_);
  or (_15418_, _15417_, _15416_);
  or (_15419_, _15418_, _15055_);
  or (_15420_, _15419_, _15401_);
  or (_15421_, _33479_, _33416_);
  or (_15422_, _15421_, _33420_);
  or (_15423_, _15422_, _15218_);
  or (_15424_, _15408_, _15405_);
  or (_15425_, _15424_, _15423_);
  or (_15426_, _15425_, _15404_);
  or (_15427_, _15426_, _15420_);
  and (_15428_, _15427_, _14923_);
  and (_15429_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_15430_, _15429_, _33493_);
  and (_15431_, _15430_, _38997_);
  or (_36877_[2], _15431_, _15428_);
  and (_15432_, _15019_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_15433_, _33202_);
  and (_15434_, _33376_, _15433_);
  or (_15435_, _15434_, _34356_);
  or (_15436_, _15376_, _15023_);
  or (_15437_, _15436_, _15435_);
  or (_15438_, _15437_, _15355_);
  or (_15439_, _15147_, _34362_);
  or (_15440_, _15439_, _15438_);
  and (_15441_, _15440_, _14923_);
  or (_36878_[0], _15441_, _15432_);
  nor (_36864_[7], _33319_, rst);
  nor (_36865_[7], _34342_, rst);
  and (_15442_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_15443_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_15444_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_15445_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_15446_, _15445_, _15444_);
  and (_15447_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_15448_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_15449_, _15448_, _15447_);
  and (_15450_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  not (_15451_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_15452_, _33146_, _15451_);
  nor (_15453_, _15452_, _15450_);
  and (_15454_, _15453_, _15449_);
  and (_15455_, _15454_, _15446_);
  nor (_15456_, _15455_, _33140_);
  nor (_15457_, _15456_, _15443_);
  nor (_15458_, _15457_, _34325_);
  nor (_15459_, _15458_, _15442_);
  nor (_36866_[7], _15459_, rst);
  nor (_36864_[0], _33222_, rst);
  and (_36864_[1], _33246_, _38997_);
  nor (_36864_[2], _33172_, rst);
  nor (_36864_[3], _33197_, rst);
  and (_36864_[4], _33271_, _38997_);
  nor (_36864_[5], _33295_, rst);
  and (_36864_[6], _33344_, _38997_);
  nor (_36865_[0], _34457_, rst);
  nor (_36865_[1], _34575_, rst);
  nor (_36865_[2], _34757_, rst);
  nor (_36865_[3], _34417_, rst);
  nor (_36865_[4], _34495_, rst);
  nor (_36865_[5], _34603_, rst);
  nor (_36865_[6], _34685_, rst);
  and (_15460_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_15461_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_15462_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_15463_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_15464_, _15463_, _15462_);
  and (_15465_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_15466_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_15467_, _15466_, _15465_);
  and (_15468_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not (_15469_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_15470_, _33146_, _15469_);
  nor (_15471_, _15470_, _15468_);
  and (_15472_, _15471_, _15467_);
  and (_15473_, _15472_, _15464_);
  nor (_15474_, _15473_, _33140_);
  nor (_15475_, _15474_, _15461_);
  nor (_15476_, _15475_, _34325_);
  nor (_15477_, _15476_, _15460_);
  nor (_36866_[0], _15477_, rst);
  and (_15478_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_15479_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_15480_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_15481_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_15482_, _15481_, _15480_);
  and (_15483_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_15484_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_15485_, _15484_, _15483_);
  and (_15486_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_15487_, _33236_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_15488_, _15487_, _15486_);
  and (_15489_, _15488_, _15485_);
  and (_15490_, _15489_, _15482_);
  nor (_15491_, _15490_, _33140_);
  nor (_15492_, _15491_, _15479_);
  nor (_15493_, _15492_, _34325_);
  nor (_15494_, _15493_, _15478_);
  nor (_36866_[1], _15494_, rst);
  and (_15495_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_15496_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_15497_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_15498_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_15499_, _15498_, _15497_);
  and (_15500_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not (_15501_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_15502_, _33146_, _15501_);
  nor (_15503_, _15502_, _15500_);
  and (_15504_, _15503_, _15499_);
  and (_15505_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_15506_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_15507_, _15506_, _15505_);
  and (_15508_, _15507_, _15504_);
  nor (_15509_, _15508_, _33140_);
  nor (_15510_, _15509_, _15496_);
  nor (_15511_, _15510_, _34325_);
  nor (_15512_, _15511_, _15495_);
  nor (_36866_[2], _15512_, rst);
  and (_15513_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_15514_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_15515_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_15516_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_15517_, _15516_, _15515_);
  and (_15518_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_15519_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_15520_, _15519_, _15518_);
  and (_15521_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not (_15522_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_15523_, _33146_, _15522_);
  nor (_15524_, _15523_, _15521_);
  and (_15525_, _15524_, _15520_);
  and (_15526_, _15525_, _15517_);
  nor (_15527_, _15526_, _33140_);
  nor (_15528_, _15527_, _15514_);
  nor (_15529_, _15528_, _34325_);
  nor (_15530_, _15529_, _15513_);
  nor (_36866_[3], _15530_, rst);
  and (_15531_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_15532_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_15533_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_15534_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_15535_, _15534_, _15533_);
  and (_15536_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_15537_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_15538_, _15537_, _15536_);
  and (_15539_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  not (_15540_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_15541_, _33146_, _15540_);
  nor (_15542_, _15541_, _15539_);
  and (_15543_, _15542_, _15538_);
  and (_15544_, _15543_, _15535_);
  nor (_15545_, _15544_, _33140_);
  nor (_15546_, _15545_, _15532_);
  nor (_15547_, _15546_, _34325_);
  nor (_15548_, _15547_, _15531_);
  nor (_36866_[4], _15548_, rst);
  and (_15549_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_15550_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_15551_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_15552_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_15553_, _15552_, _15551_);
  and (_15554_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  not (_15555_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_15556_, _33146_, _15555_);
  nor (_15557_, _15556_, _15554_);
  and (_15558_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_15559_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_15560_, _15559_, _15558_);
  and (_15561_, _15560_, _15557_);
  and (_15562_, _15561_, _15553_);
  nor (_15563_, _15562_, _33140_);
  nor (_15564_, _15563_, _15550_);
  nor (_15565_, _15564_, _34325_);
  nor (_15566_, _15565_, _15549_);
  nor (_36866_[5], _15566_, rst);
  and (_15567_, _34325_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_15568_, _33140_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_15569_, _33154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_15570_, _33150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_15571_, _15570_, _15569_);
  and (_15572_, _33162_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_15573_, _33159_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_15574_, _15573_, _15572_);
  and (_15575_, _33156_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not (_15576_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_15577_, _33146_, _15576_);
  nor (_15578_, _15577_, _15575_);
  and (_15579_, _15578_, _15574_);
  and (_15580_, _15579_, _15571_);
  nor (_15581_, _15580_, _33140_);
  nor (_15582_, _15581_, _15568_);
  nor (_15583_, _15582_, _34325_);
  nor (_15584_, _15583_, _15567_);
  nor (_36866_[6], _15584_, rst);
  and (_15585_, _33136_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_15586_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_15587_, _15585_, _14142_);
  and (_15588_, _15587_, _38997_);
  and (_36889_[15], _15588_, _15586_);
  not (_15589_, _15585_);
  or (_15590_, _15589_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00006_, _15585_, _38997_);
  and (_15591_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _38997_);
  or (_15592_, _15591_, _00006_);
  and (_36890_[15], _15592_, _15590_);
  and (_36891_, _34346_, _38997_);
  nor (_36892_[4], _34239_, rst);
  and (_36893_[7], _34320_, _38997_);
  nor (_15593_, _34529_, _34227_);
  and (_15594_, _34529_, _34227_);
  nor (_15595_, _15594_, _15593_);
  nor (_15596_, _34637_, _34232_);
  and (_15597_, _34637_, _34232_);
  nor (_15598_, _15597_, _15596_);
  and (_15599_, _15598_, _15595_);
  nor (_15600_, _34421_, _34251_);
  and (_15601_, _34421_, _34251_);
  nor (_15602_, _15601_, _15600_);
  nor (_15603_, _34691_, _33631_);
  and (_15604_, _34691_, _33631_);
  nor (_15605_, _15604_, _15603_);
  and (_15606_, _15605_, _34710_);
  and (_15607_, _15606_, _15602_);
  and (_15608_, _15607_, _15599_);
  and (_15609_, _34579_, _11341_);
  nor (_15610_, _34579_, _11341_);
  or (_15611_, _15610_, _15609_);
  nor (_15612_, _34471_, _33558_);
  and (_15613_, _34471_, _33558_);
  nor (_15614_, _15613_, _15612_);
  nor (_15615_, _15614_, _15611_);
  nor (_15616_, _34770_, _33644_);
  and (_15617_, _34770_, _33644_);
  nor (_15618_, _15617_, _15616_);
  nor (_15619_, _15618_, _13118_);
  and (_15620_, _15619_, _15615_);
  and (_15621_, _15620_, _15608_);
  nor (_15622_, _33618_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_15623_, _15622_, _15621_);
  not (_15624_, _15623_);
  not (_15625_, _33462_);
  and (_15626_, _15625_, _33362_);
  nor (_15627_, _15626_, _33467_);
  and (_15628_, _15627_, _15625_);
  nor (_15629_, _11075_, _11089_);
  and (_15630_, _15629_, _15608_);
  and (_15631_, _15630_, _15628_);
  not (_15632_, _15631_);
  nor (_15633_, _15022_, _33275_);
  not (_15634_, _33361_);
  not (_15635_, _14089_);
  not (_15636_, _15627_);
  and (_15637_, _15636_, _33463_);
  nor (_15638_, _14206_, _35617_);
  and (_15639_, _15638_, _14335_);
  and (_15640_, _15639_, _14401_);
  not (_15641_, _15640_);
  nor (_15642_, _15641_, _14469_);
  and (_15643_, _15642_, _14542_);
  and (_15644_, _15643_, _14616_);
  and (_15645_, _15644_, _15637_);
  and (_15646_, _15645_, _15635_);
  not (_15647_, _15646_);
  and (_15648_, _15628_, _33728_);
  nor (_15649_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_15650_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_15651_, _15650_, _15649_);
  nor (_15652_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_15653_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_15654_, _15653_, _15652_);
  and (_15655_, _15654_, _15651_);
  and (_15656_, _15655_, _33460_);
  and (_15657_, _33462_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_15658_, _15657_, _15656_);
  nor (_15659_, _15658_, _15648_);
  and (_15660_, _15659_, _15647_);
  or (_15661_, _15660_, _15634_);
  nor (_15662_, _15661_, _15633_);
  or (_15663_, _33382_, _33408_);
  and (_15664_, _15663_, _33252_);
  not (_15665_, _15664_);
  and (_15666_, _15063_, _33353_);
  and (_15667_, _15666_, _15665_);
  not (_15668_, _15093_);
  nor (_15669_, _15291_, _33419_);
  and (_15670_, _15669_, _15668_);
  and (_15671_, _15670_, _15667_);
  and (_15672_, _15671_, _15660_);
  nor (_15673_, _15672_, _15662_);
  nor (_15674_, _15029_, _15335_);
  and (_15675_, _15674_, _33510_);
  not (_15676_, _15675_);
  nor (_15677_, _15676_, _15673_);
  nor (_15678_, _15677_, _34367_);
  not (_15679_, _15678_);
  nor (_15680_, _15079_, _33477_);
  nor (_15681_, _15680_, _33469_);
  and (_15682_, _15681_, _15679_);
  and (_15683_, _14820_, _14836_);
  not (_15684_, _15683_);
  and (_15685_, _15684_, _33460_);
  not (_15686_, _13512_);
  nor (_15687_, _13518_, _34235_);
  and (_15688_, _15687_, _15686_);
  not (_15689_, _15688_);
  and (_15690_, _15689_, _33462_);
  nor (_15691_, _15690_, _15685_);
  not (_15692_, _15691_);
  nor (_15693_, _15692_, _15682_);
  and (_15694_, _15693_, _15632_);
  and (_15695_, _15694_, _15624_);
  and (_15696_, _15695_, _33470_);
  and (_36896_, _15696_, _38997_);
  and (_36897_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _38997_);
  and (_36898_[7], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _38997_);
  nor (_15697_, _33161_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_15698_, _15697_, _34325_);
  nor (_15699_, _15698_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_15700_, _15699_);
  and (_15701_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_15702_, _15701_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_15703_, _15702_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_15704_, _15703_, _15700_);
  and (_15705_, _15704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_15706_, _15705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_15707_, _15706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_15708_, _15707_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_15709_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_15710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_15711_, _15710_, _15709_);
  and (_15712_, _15711_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_15713_, _15712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_15714_, _15713_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_15715_, _15713_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_15716_, _15715_, _15714_);
  or (_15717_, _15716_, _15695_);
  and (_15718_, _15717_, _38997_);
  and (_15719_, _15063_, _33362_);
  nand (_15720_, _15719_, _15669_);
  nand (_15721_, _15720_, _33458_);
  and (_15722_, _33358_, _33465_);
  nand (_15723_, _15722_, _33131_);
  and (_15724_, _33350_, _33131_);
  and (_15725_, _15724_, _33252_);
  nor (_15726_, _15725_, _33469_);
  and (_15727_, _15726_, _15723_);
  and (_15728_, _15727_, _15721_);
  and (_15729_, _15728_, _34342_);
  nand (_15730_, _15727_, _15721_);
  and (_15731_, _15730_, _15459_);
  nor (_15732_, _15731_, _15729_);
  and (_15733_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_15734_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_15735_, _15734_);
  and (_15736_, _15728_, _34685_);
  and (_15737_, _15730_, _15584_);
  nor (_15738_, _15737_, _15736_);
  and (_15739_, _15738_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_15740_, _15739_);
  nor (_15741_, _15738_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_15742_, _15741_, _15739_);
  and (_15743_, _15728_, _34603_);
  and (_15744_, _15730_, _15566_);
  nor (_15745_, _15744_, _15743_);
  nor (_15746_, _15745_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_15747_, _15745_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_15748_, _15728_, _34495_);
  and (_15749_, _15730_, _15548_);
  nor (_15750_, _15749_, _15748_);
  nand (_15751_, _15750_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_15752_, _15728_, _34417_);
  and (_15753_, _15730_, _15530_);
  nor (_15754_, _15753_, _15752_);
  nor (_15755_, _15754_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_15756_, _15754_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_15757_, _34757_);
  or (_15758_, _15730_, _15757_);
  not (_15759_, _15512_);
  or (_15760_, _15728_, _15759_);
  and (_15761_, _15760_, _15758_);
  and (_15762_, _15761_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_15763_, _34575_);
  or (_15764_, _15730_, _15763_);
  not (_15765_, _15494_);
  or (_15766_, _15728_, _15765_);
  and (_15767_, _15766_, _15764_);
  nand (_15768_, _15767_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_15769_, _15768_);
  not (_15770_, _34457_);
  or (_15771_, _15730_, _15770_);
  not (_15772_, _15477_);
  or (_15773_, _15728_, _15772_);
  and (_15774_, _15773_, _15771_);
  and (_15775_, _15774_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_15776_, _15767_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_15777_, _15776_, _15768_);
  and (_15778_, _15777_, _15775_);
  or (_15779_, _15778_, _15769_);
  not (_15780_, _15762_);
  or (_15781_, _15761_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_15782_, _15781_, _15780_);
  and (_15783_, _15782_, _15779_);
  or (_15784_, _15783_, _15762_);
  nor (_15785_, _15784_, _15756_);
  nor (_15786_, _15785_, _15755_);
  or (_15787_, _15750_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_15788_, _15787_, _15751_);
  nand (_15789_, _15788_, _15786_);
  nand (_15790_, _15789_, _15751_);
  nor (_15791_, _15790_, _15747_);
  nor (_15792_, _15791_, _15746_);
  nand (_15793_, _15792_, _15742_);
  nand (_15794_, _15793_, _15740_);
  and (_15795_, _15794_, _15735_);
  or (_15796_, _15795_, _15733_);
  and (_15797_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_15798_, _15797_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_15799_, _15798_, _15796_);
  and (_15800_, _15799_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_15801_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_15802_, _15801_, _15800_);
  or (_15803_, _15802_, _15732_);
  not (_15804_, _15732_);
  or (_15805_, _15796_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_15806_, _15805_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_15807_, _15806_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_15808_, _15807_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_15809_, _15808_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_15810_, _15809_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_15811_, _15810_, _15804_);
  nand (_15812_, _15811_, _15803_);
  nor (_15813_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_15814_, _15732_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_15815_, _15814_, _15813_);
  or (_15816_, _15815_, _15812_);
  nor (_15817_, _15816_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_15818_, _15816_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_15819_, _15818_, _15817_);
  and (_15820_, _15063_, _15022_);
  and (_15821_, _15820_, _33362_);
  and (_15822_, _15821_, _15674_);
  and (_15823_, _15822_, _15670_);
  nor (_15824_, _15823_, _34367_);
  nor (_15825_, _15824_, _15725_);
  nor (_15826_, _33484_, _34367_);
  nor (_15827_, _15826_, _15680_);
  not (_15828_, _15827_);
  and (_15829_, _15828_, _15728_);
  nor (_15830_, _15829_, _15825_);
  and (_15831_, _15830_, _15819_);
  nor (_15832_, _14098_, _33470_);
  not (_15833_, _15826_);
  nor (_15834_, _15833_, _14189_);
  not (_15835_, _34342_);
  and (_15836_, _15828_, _15730_);
  and (_15837_, _15836_, _15835_);
  and (_15838_, _33252_, _33131_);
  and (_15839_, _15838_, _33350_);
  not (_15840_, _15839_);
  not (_15841_, _33468_);
  nor (_15842_, _15841_, _33442_);
  and (_15843_, _15078_, _33131_);
  nor (_15844_, _15843_, _15842_);
  and (_15845_, _15844_, _15721_);
  and (_15846_, _15845_, _15840_);
  nor (_15847_, _15828_, _15824_);
  and (_15848_, _15847_, _15846_);
  and (_15849_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_15850_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_15851_, _15850_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_15852_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_15853_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_15854_, _15853_, _15852_);
  and (_15855_, _15854_, _15851_);
  and (_15856_, _15855_, _15798_);
  and (_15857_, _15856_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_15858_, _15857_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_15859_, _15858_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_15860_, _15859_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_15861_, _15860_, _14142_);
  or (_15862_, _15860_, _14142_);
  and (_15863_, _15862_, _15861_);
  not (_15864_, _15824_);
  and (_15865_, _15829_, _15864_);
  and (_15866_, _15865_, _15863_);
  or (_15867_, _15866_, _15849_);
  or (_15868_, _15867_, _15837_);
  nor (_15869_, _15868_, _15834_);
  nand (_15870_, _15869_, _15695_);
  or (_15871_, _15870_, _15832_);
  or (_15872_, _15871_, _15831_);
  and (_36899_[15], _15872_, _15718_);
  and (_15873_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _38997_);
  and (_15874_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_15875_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_15876_, _33135_, _15875_);
  not (_15877_, _15876_);
  not (_15878_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_15879_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_15880_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_15881_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_15882_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_15883_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_15884_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_15885_, _15884_, _15882_);
  and (_15886_, _15885_, _15883_);
  nor (_15887_, _15886_, _15882_);
  nor (_15888_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_15889_, _15888_, _15881_);
  not (_15890_, _15889_);
  nor (_15891_, _15890_, _15887_);
  nor (_15892_, _15891_, _15881_);
  not (_15893_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_15894_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_15895_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_15896_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_15897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_15898_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_15899_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_15900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_15901_, _15900_, _15899_);
  and (_15902_, _15901_, _15898_);
  and (_15903_, _15902_, _15897_);
  and (_15904_, _15903_, _15896_);
  and (_15905_, _15904_, _15895_);
  and (_15906_, _15905_, _15894_);
  and (_15907_, _15906_, _15893_);
  and (_15908_, _15907_, _15892_);
  and (_15909_, _15908_, _15880_);
  and (_15910_, _15909_, _15879_);
  and (_15911_, _15910_, _15878_);
  nor (_15912_, _15911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_15913_, _15911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_15914_, _15913_, _15912_);
  nor (_15915_, _15910_, _15878_);
  nor (_15916_, _15915_, _15911_);
  not (_15917_, _15916_);
  nor (_15918_, _15909_, _15879_);
  nor (_15919_, _15918_, _15910_);
  not (_15920_, _15919_);
  nor (_15921_, _15908_, _15880_);
  nor (_15922_, _15921_, _15909_);
  not (_15923_, _15922_);
  and (_15924_, _15892_, _15906_);
  nor (_15925_, _15924_, _15893_);
  nor (_15926_, _15925_, _15908_);
  not (_15927_, _15926_);
  and (_15928_, _15892_, _15904_);
  and (_15929_, _15928_, _15895_);
  nor (_15930_, _15929_, _15894_);
  or (_15931_, _15930_, _15924_);
  nor (_15932_, _15928_, _15895_);
  nor (_15933_, _15932_, _15929_);
  not (_15934_, _15933_);
  and (_15935_, _15892_, _15902_);
  nor (_15936_, _15935_, _15897_);
  and (_15937_, _15892_, _15903_);
  nor (_15938_, _15937_, _15936_);
  not (_15939_, _15938_);
  and (_15940_, _15892_, _15901_);
  nor (_15941_, _15940_, _15898_);
  nor (_15942_, _15941_, _15935_);
  not (_15943_, _15942_);
  and (_15944_, _15892_, _15900_);
  nor (_15945_, _15944_, _15899_);
  nor (_15946_, _15945_, _15940_);
  not (_15947_, _15946_);
  not (_15948_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_15949_, _15892_, _15948_);
  nor (_15950_, _15892_, _15948_);
  nor (_15951_, _15950_, _15949_);
  not (_15952_, _15951_);
  not (_15953_, _14966_);
  and (_15954_, _14962_, _14932_);
  not (_15955_, _15954_);
  and (_15956_, _14954_, _14974_);
  nor (_15957_, _15956_, _14980_);
  and (_15958_, _15957_, _15955_);
  and (_15959_, _14976_, _14943_);
  and (_15960_, _14943_, _14974_);
  or (_15961_, _15960_, _15959_);
  not (_15962_, _15961_);
  nor (_15963_, _14996_, _14945_);
  and (_15964_, _15963_, _15962_);
  and (_15965_, _15964_, _15958_);
  nor (_15966_, _15965_, _15953_);
  not (_15967_, _15966_);
  not (_15968_, _14967_);
  and (_15969_, _14959_, _14944_);
  nor (_15970_, _15969_, _14981_);
  nor (_15971_, _15970_, _15968_);
  not (_15972_, _15971_);
  and (_15973_, _15972_, _14995_);
  and (_15974_, _15973_, _15967_);
  and (_15975_, _15960_, _14929_);
  and (_15976_, _14966_, _14963_);
  nor (_15977_, _15976_, _15975_);
  nor (_15978_, _14965_, _14942_);
  not (_15979_, _15978_);
  and (_15980_, _15979_, _14986_);
  and (_15981_, _14976_, _14932_);
  and (_15982_, _15981_, _14981_);
  nor (_15983_, _15982_, _15980_);
  and (_15984_, _15983_, _15977_);
  and (_15985_, _14954_, _14930_);
  and (_15986_, _15985_, _14951_);
  not (_15987_, _15986_);
  and (_15988_, _33246_, _14935_);
  and (_15989_, _15988_, _14943_);
  and (_15990_, _15989_, _14941_);
  nor (_15991_, _15990_, _14938_);
  and (_15992_, _15991_, _15987_);
  not (_15993_, _33197_);
  and (_15994_, _14963_, _15993_);
  and (_15995_, _15956_, _14942_);
  nor (_15996_, _15995_, _15994_);
  and (_15997_, _15996_, _15992_);
  and (_15998_, _15997_, _14957_);
  and (_15999_, _15998_, _15984_);
  and (_16000_, _14990_, _33222_);
  and (_16001_, _16000_, _15979_);
  not (_16002_, _16001_);
  and (_16003_, _14997_, _14990_);
  not (_16004_, _14959_);
  nor (_16005_, _15960_, _14996_);
  nor (_16006_, _16005_, _16004_);
  nor (_16007_, _16006_, _16003_);
  and (_16008_, _16007_, _16002_);
  and (_16009_, _14945_, _14929_);
  nor (_16010_, _15959_, _14996_);
  nor (_16011_, _16010_, _33197_);
  nor (_16012_, _16011_, _16009_);
  nor (_16013_, _15959_, _14937_);
  not (_16014_, _16013_);
  and (_16015_, _16014_, _14929_);
  or (_16016_, _14963_, _14996_);
  and (_16017_, _16016_, _14981_);
  nor (_16018_, _16017_, _16015_);
  and (_16019_, _16018_, _16012_);
  and (_16020_, _16019_, _16008_);
  and (_16021_, _16020_, _15999_);
  and (_16022_, _14981_, _14945_);
  and (_16023_, _14997_, _15956_);
  nor (_16024_, _16023_, _16022_);
  and (_16025_, _14959_, _14945_);
  not (_16026_, _16025_);
  and (_16027_, _16026_, _14983_);
  and (_16028_, _16027_, _16024_);
  not (_16029_, _14981_);
  nor (_16030_, _15954_, _15960_);
  and (_16031_, _14944_, _14932_);
  nor (_16032_, _16031_, _14990_);
  and (_16033_, _16032_, _16030_);
  nor (_16034_, _16033_, _16029_);
  not (_16035_, _16034_);
  and (_16036_, _14977_, _14959_);
  nor (_16037_, _16036_, _14971_);
  and (_16038_, _16037_, _16035_);
  and (_16039_, _16038_, _16028_);
  and (_16040_, _16039_, _16021_);
  and (_16041_, _16040_, _15974_);
  nor (_16042_, _15885_, _15883_);
  nor (_16043_, _16042_, _15886_);
  not (_16044_, _16043_);
  nor (_16045_, _16044_, _16041_);
  not (_16046_, _16045_);
  and (_16047_, _14997_, _14986_);
  or (_16048_, _16003_, _16047_);
  or (_16049_, _16017_, _15975_);
  or (_16050_, _14993_, _14969_);
  or (_16051_, _16050_, _16049_);
  or (_16052_, _16051_, _16048_);
  not (_16053_, _14953_);
  nand (_16054_, _16028_, _16053_);
  or (_16055_, _16054_, _16052_);
  nor (_16056_, _16055_, _16041_);
  not (_16057_, _16056_);
  nor (_16058_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_16059_, _16058_, _15883_);
  and (_16060_, _16059_, _16057_);
  and (_16061_, _16044_, _16041_);
  nor (_16062_, _16061_, _16045_);
  nand (_16063_, _16062_, _16060_);
  and (_16064_, _16063_, _16046_);
  not (_16065_, _16064_);
  and (_16066_, _15890_, _15887_);
  nor (_16067_, _16066_, _15891_);
  and (_16068_, _16067_, _16065_);
  and (_16069_, _16068_, _15952_);
  not (_16070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_16071_, _15949_, _16070_);
  or (_16072_, _16071_, _15944_);
  and (_16073_, _16072_, _16069_);
  and (_16074_, _16073_, _15947_);
  and (_16075_, _16074_, _15943_);
  and (_16076_, _16075_, _15939_);
  nor (_16077_, _15937_, _15896_);
  or (_16078_, _16077_, _15928_);
  and (_16079_, _16078_, _16076_);
  and (_16080_, _16079_, _15934_);
  and (_16081_, _16080_, _15931_);
  and (_16082_, _16081_, _15927_);
  and (_16083_, _16082_, _15923_);
  and (_16084_, _16083_, _15920_);
  and (_16085_, _16084_, _15917_);
  or (_16086_, _16085_, _15914_);
  nand (_16087_, _16085_, _15914_);
  and (_16088_, _16087_, _16086_);
  or (_16089_, _16088_, _15877_);
  or (_16090_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_16091_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_16092_, _16091_, _16090_);
  and (_16093_, _16092_, _16089_);
  or (_36900_[15], _16093_, _15874_);
  nor (_16094_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_36901_, _16094_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_36902_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _38997_);
  not (_16095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_16096_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_16097_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_16098_, _16097_, _16096_);
  not (_16099_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_16100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_16101_, _16100_, _16099_);
  and (_16102_, _16101_, _16098_);
  and (_16103_, _16102_, _16095_);
  and (_16104_, \oc8051_top_1.oc8051_rom1.ea_int , _33132_);
  nand (_16105_, _16104_, _33135_);
  nand (_16106_, _16105_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_16107_, _16106_, _16103_);
  and (_36903_, _16107_, _38997_);
  and (_16108_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_16109_, _16108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_36904_[7], _16109_, _38997_);
  nor (_16110_, _15699_, _34325_);
  nor (_16111_, _16041_, _33148_);
  not (_16112_, _16111_);
  nor (_16113_, _16056_, _33144_);
  and (_16114_, _16041_, _33148_);
  nor (_16115_, _16114_, _16111_);
  nand (_16116_, _16115_, _16113_);
  and (_16117_, _16116_, _16112_);
  nor (_16118_, _16117_, _34325_);
  and (_16119_, _16118_, _33143_);
  nor (_16120_, _16118_, _33143_);
  nor (_16121_, _16120_, _16119_);
  nor (_16122_, _16121_, _16110_);
  and (_16123_, _33149_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_16124_, _16123_, _16110_);
  and (_16125_, _16124_, _16055_);
  or (_16126_, _16125_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_16127_, _16126_, _16122_);
  and (_36905_[2], _16127_, _38997_);
  and (_16128_, _33240_, _33265_);
  and (_16129_, _33338_, _33313_);
  and (_16130_, _16129_, _16128_);
  and (_16131_, _33136_, _38997_);
  and (_16132_, _16131_, _33191_);
  and (_16133_, _16132_, _33217_);
  and (_16134_, _33167_, _33290_);
  and (_16135_, _16134_, _16133_);
  and (_36908_, _16135_, _16130_);
  nor (_16136_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_16137_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_16138_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_36910_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _38997_);
  and (_16139_, _36910_, _16138_);
  or (_36909_[7], _16139_, _16137_);
  not (_16140_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_16141_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_16142_, _16141_, _16140_);
  and (_16143_, _16141_, _16140_);
  nor (_16144_, _16143_, _16142_);
  not (_16145_, _16144_);
  and (_16146_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_16147_, _16146_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_16148_, _16146_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_16149_, _16148_, _16147_);
  or (_16150_, _16149_, _16141_);
  and (_16151_, _16150_, _16145_);
  nor (_16152_, _16142_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_16153_, _16142_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_16154_, _16153_, _16152_);
  or (_16155_, _16147_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_36912_[3], _16155_, _38997_);
  and (_16156_, _36912_[3], _16154_);
  and (_36911_, _16156_, _16151_);
  not (_16157_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_16158_, _15699_, _16157_);
  and (_16159_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_16160_, _16158_);
  and (_16161_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_16162_, _16161_, _16159_);
  and (_36913_[31], _16162_, _38997_);
  and (_16163_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_16164_, _16158_, _34334_);
  or (_16165_, _16164_, _16163_);
  and (_36914_[31], _16165_, _38997_);
  and (_16166_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_16167_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16168_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _16167_);
  and (_16169_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_16170_, _16169_, _16166_);
  and (_36915_[7], _16170_, _38997_);
  and (_16171_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  or (_16172_, _16171_, _16168_);
  and (_36916_, _16172_, _38997_);
  or (_16173_, _16167_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_36917_, _16173_, _38997_);
  not (_16174_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_16175_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_16176_, _16175_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_16177_, _16167_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_16178_, _16177_, _38997_);
  and (_36918_[15], _16178_, _16176_);
  or (_16179_, _16167_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_36919_, _16179_, _38997_);
  nor (_16180_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_16181_, _16180_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16182_, _16181_, _38997_);
  and (_16183_, _36910_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_36920_, _16183_, _16182_);
  and (_16184_, _16157_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_16185_, _16184_, _16181_);
  and (_36921_, _16185_, _38997_);
  nand (_16186_, _16181_, _14189_);
  or (_16187_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_16188_, _16187_, _38997_);
  and (_36922_[15], _16188_, _16186_);
  and (_16189_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_16190_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_16191_, _15585_, _16190_);
  or (_16192_, _16191_, _16189_);
  and (_36889_[0], _16192_, _38997_);
  and (_16193_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_16194_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_16195_, _15585_, _16194_);
  or (_16196_, _16195_, _16193_);
  and (_36889_[1], _16196_, _38997_);
  and (_16197_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_16198_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_16199_, _15585_, _16198_);
  or (_16200_, _16199_, _16197_);
  and (_36889_[2], _16200_, _38997_);
  and (_16201_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_16202_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_16203_, _15585_, _16202_);
  or (_16204_, _16203_, _16201_);
  and (_36889_[3], _16204_, _38997_);
  and (_16205_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_16206_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_16207_, _15585_, _16206_);
  or (_16208_, _16207_, _16205_);
  and (_36889_[4], _16208_, _38997_);
  and (_16209_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_16210_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_16211_, _15585_, _16210_);
  or (_16212_, _16211_, _16209_);
  and (_36889_[5], _16212_, _38997_);
  and (_16213_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_16214_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_16215_, _15585_, _16214_);
  or (_16216_, _16215_, _16213_);
  and (_36889_[6], _16216_, _38997_);
  and (_16217_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_16218_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_16219_, _15585_, _16218_);
  or (_16220_, _16219_, _16217_);
  and (_36889_[7], _16220_, _38997_);
  and (_16221_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_16222_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_16223_, _15585_, _16222_);
  or (_16224_, _16223_, _16221_);
  and (_36889_[8], _16224_, _38997_);
  and (_16225_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_16226_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_16227_, _15585_, _16226_);
  or (_16228_, _16227_, _16225_);
  and (_36889_[9], _16228_, _38997_);
  and (_16229_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_16230_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_16231_, _15585_, _16230_);
  or (_16232_, _16231_, _16229_);
  and (_36889_[10], _16232_, _38997_);
  and (_16233_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_16234_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_16235_, _15585_, _16234_);
  or (_16236_, _16235_, _16233_);
  and (_36889_[11], _16236_, _38997_);
  and (_16237_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_16238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_16239_, _15585_, _16238_);
  or (_16240_, _16239_, _16237_);
  and (_36889_[12], _16240_, _38997_);
  and (_16241_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_16242_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_16243_, _15585_, _16242_);
  or (_16244_, _16243_, _16241_);
  and (_36889_[13], _16244_, _38997_);
  and (_16245_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_16246_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_16247_, _15585_, _16246_);
  or (_16248_, _16247_, _16245_);
  and (_36889_[14], _16248_, _38997_);
  or (_16249_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_16250_, _15585_, _16190_);
  and (_16251_, _16250_, _38997_);
  and (_36890_[0], _16251_, _16249_);
  or (_16252_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand (_16253_, _15585_, _16194_);
  and (_16254_, _16253_, _38997_);
  and (_36890_[1], _16254_, _16252_);
  or (_16255_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand (_16256_, _15585_, _16198_);
  and (_16257_, _16256_, _38997_);
  and (_36890_[2], _16257_, _16255_);
  or (_16258_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand (_16259_, _15585_, _16202_);
  and (_16260_, _16259_, _38997_);
  and (_36890_[3], _16260_, _16258_);
  or (_16261_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nand (_16262_, _15585_, _16206_);
  and (_16263_, _16262_, _38997_);
  and (_36890_[4], _16263_, _16261_);
  or (_16264_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand (_16265_, _15585_, _16210_);
  and (_16266_, _16265_, _38997_);
  and (_36890_[5], _16266_, _16264_);
  or (_16267_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand (_16268_, _15585_, _16214_);
  and (_16269_, _16268_, _38997_);
  and (_36890_[6], _16269_, _16267_);
  or (_16270_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nand (_16271_, _15585_, _16218_);
  and (_16272_, _16271_, _38997_);
  and (_36890_[7], _16272_, _16270_);
  or (_16273_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nand (_16274_, _15585_, _16222_);
  and (_16275_, _16274_, _38997_);
  and (_36890_[8], _16275_, _16273_);
  or (_16276_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nand (_16277_, _15585_, _16226_);
  and (_16278_, _16277_, _38997_);
  and (_36890_[9], _16278_, _16276_);
  or (_16279_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand (_16280_, _15585_, _16230_);
  and (_16281_, _16280_, _38997_);
  and (_36890_[10], _16281_, _16279_);
  or (_16282_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand (_16283_, _15585_, _16234_);
  and (_16284_, _16283_, _38997_);
  and (_36890_[11], _16284_, _16282_);
  or (_16285_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nand (_16286_, _15585_, _16238_);
  and (_16287_, _16286_, _38997_);
  and (_36890_[12], _16287_, _16285_);
  or (_16288_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nand (_16289_, _15585_, _16242_);
  and (_16290_, _16289_, _38997_);
  and (_36890_[13], _16290_, _16288_);
  or (_16291_, _15585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand (_16292_, _15585_, _16246_);
  and (_16293_, _16292_, _38997_);
  and (_36890_[14], _16293_, _16291_);
  and (_36892_[0], _33226_, _38997_);
  and (_36892_[1], _33250_, _38997_);
  and (_36892_[2], _33177_, _38997_);
  nor (_36892_[3], _34283_, rst);
  nor (_16294_, _16158_, _15469_);
  and (_16295_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_16296_, _16295_, _16294_);
  and (_36913_[0], _16296_, _38997_);
  and (_16297_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_16298_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_16299_, _16298_, _16158_);
  or (_16300_, _16299_, _16297_);
  and (_36913_[1], _16300_, _38997_);
  nor (_16301_, _16158_, _15501_);
  and (_16302_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_16303_, _16302_, _16301_);
  and (_36913_[2], _16303_, _38997_);
  nor (_16304_, _16158_, _15522_);
  and (_16305_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_16306_, _16305_, _16158_);
  or (_16307_, _16306_, _16304_);
  and (_36913_[3], _16307_, _38997_);
  nor (_16308_, _16158_, _15540_);
  and (_16309_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_16310_, _16309_, _16308_);
  and (_36913_[4], _16310_, _38997_);
  nor (_16311_, _16158_, _15555_);
  and (_16312_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_16313_, _16312_, _16311_);
  and (_36913_[5], _16313_, _38997_);
  nor (_16314_, _16158_, _15576_);
  and (_16315_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_16316_, _16315_, _16158_);
  or (_16317_, _16316_, _16314_);
  and (_36913_[6], _16317_, _38997_);
  nor (_16318_, _16158_, _15451_);
  and (_16319_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_16320_, _16319_, _16318_);
  and (_36913_[7], _16320_, _38997_);
  and (_16321_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_16322_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_16323_, _16322_, _16321_);
  and (_36913_[8], _16323_, _38997_);
  and (_16324_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_16325_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_16326_, _16325_, _16324_);
  and (_36913_[9], _16326_, _38997_);
  and (_16327_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_16328_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_16329_, _16328_, _16327_);
  and (_36913_[10], _16329_, _38997_);
  and (_16330_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_16331_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_16332_, _16331_, _16330_);
  and (_36913_[11], _16332_, _38997_);
  and (_16333_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_16334_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_16335_, _16334_, _16333_);
  and (_36913_[12], _16335_, _38997_);
  and (_16336_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_16337_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_16338_, _16337_, _16336_);
  and (_36913_[13], _16338_, _38997_);
  and (_16339_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_16340_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_16341_, _16340_, _16339_);
  and (_36913_[14], _16341_, _38997_);
  and (_16342_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_16343_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_16344_, _16343_, _16342_);
  and (_36913_[15], _16344_, _38997_);
  and (_16345_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_16346_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_16347_, _16346_, _16345_);
  and (_36913_[16], _16347_, _38997_);
  and (_16348_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_16349_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_16350_, _16349_, _16348_);
  and (_36913_[17], _16350_, _38997_);
  and (_16351_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_16352_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_16353_, _16352_, _16351_);
  and (_36913_[18], _16353_, _38997_);
  and (_16354_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_16355_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_16356_, _16355_, _16354_);
  and (_36913_[19], _16356_, _38997_);
  and (_16357_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_16358_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_16359_, _16358_, _16357_);
  and (_36913_[20], _16359_, _38997_);
  and (_16360_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_16361_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_16362_, _16361_, _16360_);
  and (_36913_[21], _16362_, _38997_);
  and (_16363_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_16364_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_16365_, _16364_, _16363_);
  and (_36913_[22], _16365_, _38997_);
  and (_16366_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_16367_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_16368_, _16367_, _16366_);
  and (_36913_[23], _16368_, _38997_);
  and (_16369_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_16370_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_16371_, _16370_, _16369_);
  and (_36913_[24], _16371_, _38997_);
  and (_16372_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_16373_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_16374_, _16373_, _16372_);
  and (_36913_[25], _16374_, _38997_);
  and (_16375_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_16376_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_16377_, _16376_, _16375_);
  and (_36913_[26], _16377_, _38997_);
  and (_16378_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_16379_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_16380_, _16379_, _16378_);
  and (_36913_[27], _16380_, _38997_);
  and (_16381_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_16382_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_16383_, _16382_, _16381_);
  and (_36913_[28], _16383_, _38997_);
  and (_16384_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_16385_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_16386_, _16385_, _16384_);
  and (_36913_[29], _16386_, _38997_);
  and (_16387_, _16158_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_16388_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_16389_, _16388_, _16387_);
  and (_36913_[30], _16389_, _38997_);
  nor (_36893_[0], _34441_, rst);
  nor (_36893_[1], _34548_, rst);
  nor (_36893_[2], _34741_, rst);
  nor (_36893_[3], _34391_, rst);
  nor (_36893_[4], _34517_, rst);
  nor (_36893_[5], _34634_, rst);
  nor (_36893_[6], _34669_, rst);
  and (_36898_[0], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _38997_);
  and (_36898_[1], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _38997_);
  and (_36898_[2], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _38997_);
  and (_36898_[3], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _38997_);
  and (_36898_[4], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _38997_);
  and (_36898_[5], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _38997_);
  and (_36898_[6], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _38997_);
  not (_16390_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_16391_, _15696_, _16390_);
  and (_16392_, _15021_, _33458_);
  and (_16393_, _15689_, _16392_);
  nor (_16394_, _15680_, _15842_);
  and (_16395_, _16394_, _15679_);
  nor (_16396_, _16395_, _16393_);
  and (_16397_, _16396_, _15632_);
  and (_16398_, _15621_, _34706_);
  and (_16399_, _16398_, _33658_);
  nor (_16400_, _16399_, _15685_);
  and (_16401_, _16400_, _16397_);
  or (_16402_, _15848_, _15826_);
  and (_16403_, _16402_, _14223_);
  nor (_16404_, _15827_, _15844_);
  and (_16405_, _16404_, _15772_);
  and (_16406_, _15828_, _15846_);
  and (_16407_, _16406_, _15864_);
  and (_16408_, _16407_, _15770_);
  or (_16409_, _16408_, _16405_);
  nor (_16410_, _15824_, _15839_);
  nor (_16411_, _16406_, _16410_);
  nor (_16412_, _15774_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_16413_, _16412_, _15775_);
  and (_16414_, _16413_, _16411_);
  or (_16415_, _16414_, _16409_);
  or (_16416_, _16415_, _16403_);
  and (_16417_, _16416_, _16401_);
  or (_16418_, _16417_, _16391_);
  and (_36899_[0], _16418_, _38997_);
  nand (_16419_, _16402_, _14289_);
  nand (_16420_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nand (_16421_, _16404_, _15765_);
  nand (_16422_, _16407_, _15763_);
  and (_16423_, _16422_, _16421_);
  and (_16424_, _16423_, _16420_);
  or (_16425_, _15777_, _15775_);
  nand (_16426_, _16425_, _16411_);
  or (_16427_, _16426_, _15778_);
  and (_16428_, _16427_, _16424_);
  and (_16429_, _16428_, _16419_);
  nand (_16430_, _16429_, _16401_);
  or (_16431_, _16401_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_16432_, _16431_, _38997_);
  and (_36899_[1], _16432_, _16430_);
  and (_16433_, _16402_, _14724_);
  and (_16434_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_16435_, _16404_, _15759_);
  and (_16436_, _16407_, _15757_);
  or (_16437_, _16436_, _16435_);
  or (_16438_, _16437_, _16434_);
  or (_16439_, _16438_, _16433_);
  not (_16440_, _15783_);
  or (_16441_, _15782_, _15779_);
  and (_16442_, _16441_, _16440_);
  nand (_16443_, _16442_, _16411_);
  nand (_16444_, _16443_, _16401_);
  or (_16445_, _16444_, _16439_);
  not (_16446_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_16447_, _15699_, _16446_);
  and (_16448_, _15699_, _16446_);
  nor (_16449_, _16448_, _16447_);
  or (_16450_, _16449_, _16401_);
  and (_16451_, _16450_, _38997_);
  and (_36899_[2], _16451_, _16445_);
  and (_16452_, _16402_, _14740_);
  not (_16453_, _15530_);
  and (_16454_, _16404_, _16453_);
  not (_16455_, _34417_);
  and (_16456_, _16407_, _16455_);
  or (_16457_, _16456_, _16454_);
  or (_16458_, _15755_, _15756_);
  not (_16459_, _16458_);
  nand (_16460_, _16459_, _15784_);
  or (_16461_, _16459_, _15784_);
  and (_16462_, _16461_, _16411_);
  and (_16463_, _16462_, _16460_);
  or (_16464_, _16463_, _16457_);
  or (_16465_, _16464_, _16452_);
  nand (_16466_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand (_16467_, _16466_, _16401_);
  or (_16468_, _16467_, _16465_);
  and (_16469_, _16447_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_16470_, _16447_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_16471_, _16470_, _16469_);
  or (_16472_, _16471_, _16401_);
  and (_16473_, _16472_, _38997_);
  and (_36899_[3], _16473_, _16468_);
  and (_16474_, _15702_, _15700_);
  nor (_16475_, _16469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_16476_, _16475_, _16474_);
  or (_16477_, _16476_, _15695_);
  and (_16478_, _16477_, _38997_);
  and (_16479_, _16402_, _14494_);
  or (_16480_, _15788_, _15786_);
  and (_16481_, _15830_, _15789_);
  and (_16482_, _16481_, _16480_);
  not (_16483_, _15548_);
  and (_16484_, _15836_, _16483_);
  not (_16485_, _34495_);
  and (_16486_, _15865_, _16485_);
  and (_16487_, _33469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_16488_, _16487_, _16486_);
  or (_16489_, _16488_, _16484_);
  nor (_16490_, _16489_, _16482_);
  nand (_16491_, _16490_, _15695_);
  or (_16492_, _16491_, _16479_);
  and (_36899_[4], _16492_, _16478_);
  nor (_16493_, _16474_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_16494_, _16493_, _15704_);
  or (_16495_, _16494_, _15695_);
  and (_16496_, _16495_, _38997_);
  and (_16497_, _16402_, _14767_);
  or (_16498_, _15746_, _15747_);
  and (_16499_, _16498_, _15790_);
  nor (_16500_, _16498_, _15790_);
  or (_16501_, _16500_, _16499_);
  and (_16502_, _16501_, _15830_);
  not (_16503_, _15566_);
  and (_16504_, _15836_, _16503_);
  not (_16505_, _34603_);
  and (_16506_, _15865_, _16505_);
  and (_16507_, _33469_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_16508_, _16507_, _16506_);
  or (_16509_, _16508_, _16504_);
  nor (_16510_, _16509_, _16502_);
  nand (_16511_, _16510_, _15695_);
  or (_16512_, _16511_, _16497_);
  and (_36899_[5], _16512_, _16496_);
  nor (_16513_, _15704_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_16514_, _16513_, _15705_);
  or (_16515_, _16514_, _15695_);
  and (_16516_, _16515_, _38997_);
  and (_16517_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_16518_, _16402_, _14632_);
  not (_16519_, _15584_);
  and (_16520_, _16404_, _16519_);
  and (_16521_, _16407_, _34686_);
  or (_16522_, _16521_, _16520_);
  or (_16523_, _15792_, _15742_);
  and (_16524_, _16411_, _15793_);
  and (_16525_, _16524_, _16523_);
  or (_16526_, _16525_, _16522_);
  or (_16527_, _16526_, _16518_);
  nor (_16528_, _16527_, _16517_);
  nand (_16529_, _16528_, _16401_);
  and (_36899_[6], _16529_, _16516_);
  nor (_16530_, _15705_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_16531_, _16530_, _15706_);
  or (_16532_, _16531_, _15695_);
  and (_16533_, _16532_, _38997_);
  or (_16534_, _15733_, _15734_);
  and (_16535_, _16534_, _15794_);
  nor (_16536_, _16534_, _15794_);
  or (_16537_, _16536_, _16535_);
  and (_16538_, _16537_, _16411_);
  and (_16539_, _16402_, _14683_);
  and (_16540_, _15842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_16541_, _15459_);
  and (_16542_, _16404_, _16541_);
  and (_16543_, _16407_, _15835_);
  or (_16544_, _16543_, _16542_);
  or (_16545_, _16544_, _16540_);
  or (_16546_, _16545_, _16539_);
  nor (_16547_, _16546_, _16538_);
  nand (_16548_, _16547_, _16401_);
  and (_36899_[7], _16548_, _16533_);
  nor (_16549_, _15706_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_16550_, _16549_, _15707_);
  or (_16551_, _16550_, _15695_);
  and (_16552_, _16551_, _38997_);
  and (_16553_, _15796_, _14110_);
  nor (_16554_, _15796_, _14110_);
  nor (_16555_, _16554_, _16553_);
  nor (_16556_, _16555_, _15732_);
  and (_16557_, _16555_, _15732_);
  or (_16558_, _16557_, _16556_);
  and (_16559_, _16558_, _15830_);
  and (_16560_, _14223_, _33469_);
  and (_16561_, _15826_, _14250_);
  nand (_16562_, _15836_, _15770_);
  and (_16563_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_16564_, _15865_, _14930_);
  nor (_16565_, _16564_, _16563_);
  and (_16566_, _16565_, _16562_);
  nand (_16567_, _16566_, _15695_);
  or (_16568_, _16567_, _16561_);
  or (_16569_, _16568_, _16560_);
  or (_16570_, _16569_, _16559_);
  and (_36899_[8], _16570_, _16552_);
  nor (_16571_, _15707_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_16572_, _16571_, _15708_);
  or (_16573_, _16572_, _15695_);
  and (_16574_, _16573_, _38997_);
  and (_16575_, _15796_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_16576_, _16575_, _15804_);
  nor (_16577_, _15805_, _15804_);
  nor (_16578_, _16577_, _16576_);
  nand (_16579_, _16578_, _14116_);
  or (_16580_, _16578_, _14116_);
  and (_16581_, _16580_, _15830_);
  and (_16582_, _16581_, _16579_);
  and (_16583_, _14289_, _33469_);
  nor (_16584_, _15833_, _14323_);
  and (_16585_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_16586_, _15836_, _15763_);
  or (_16587_, _16586_, _16585_);
  and (_16588_, _15865_, _33344_);
  or (_16589_, _16588_, _16587_);
  nor (_16590_, _16589_, _16584_);
  nand (_16591_, _16590_, _15695_);
  or (_16592_, _16591_, _16583_);
  or (_16593_, _16592_, _16582_);
  and (_36899_[9], _16593_, _16574_);
  nor (_16594_, _15708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_16595_, _16594_, _15709_);
  or (_16596_, _16595_, _15695_);
  and (_16597_, _16596_, _38997_);
  and (_16598_, _16577_, _14116_);
  and (_16599_, _16576_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_16600_, _16599_, _16598_);
  nand (_16601_, _16600_, _14121_);
  or (_16602_, _16600_, _14121_);
  and (_16603_, _16602_, _15830_);
  and (_16604_, _16603_, _16601_);
  nor (_16605_, _14356_, _33470_);
  nor (_16606_, _15833_, _14387_);
  and (_16607_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_16608_, _15836_, _15757_);
  and (_16609_, _15865_, _14931_);
  or (_16610_, _16609_, _16608_);
  or (_16611_, _16610_, _16607_);
  nor (_16612_, _16611_, _16606_);
  nand (_16613_, _16612_, _15695_);
  or (_16614_, _16613_, _16605_);
  or (_16615_, _16614_, _16604_);
  and (_36899_[10], _16615_, _16597_);
  nor (_16616_, _15709_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_16617_, _15709_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_16618_, _16617_, _16616_);
  or (_16619_, _16618_, _15695_);
  and (_16620_, _16619_, _38997_);
  and (_16621_, _15799_, _15804_);
  nor (_16622_, _15807_, _15804_);
  nor (_16623_, _16622_, _16621_);
  nor (_16624_, _16623_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_16625_, _16623_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_16626_, _16625_, _16624_);
  and (_16627_, _16626_, _15830_);
  nor (_16628_, _14423_, _33470_);
  nor (_16629_, _15833_, _14456_);
  and (_16630_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_16631_, _15836_, _16455_);
  or (_16632_, _16631_, _16630_);
  nor (_16633_, _15856_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_16634_, _16633_, _15857_);
  and (_16635_, _16634_, _15865_);
  or (_16636_, _16635_, _16632_);
  nor (_16637_, _16636_, _16629_);
  nand (_16638_, _16637_, _15695_);
  or (_16639_, _16638_, _16628_);
  or (_16640_, _16639_, _16627_);
  and (_36899_[11], _16640_, _16620_);
  nor (_16641_, _16617_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_16642_, _16641_, _15711_);
  or (_16643_, _16642_, _15695_);
  and (_16644_, _16643_, _38997_);
  nor (_16645_, _15808_, _15804_);
  and (_16646_, _15800_, _15804_);
  or (_16647_, _16646_, _16645_);
  nand (_16648_, _16647_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_16649_, _16647_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_16650_, _16649_, _15830_);
  and (_16651_, _16650_, _16648_);
  and (_16652_, _14494_, _33469_);
  nor (_16653_, _15833_, _14529_);
  and (_16654_, _15836_, _16485_);
  and (_16655_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_16656_, _15857_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_16657_, _16656_, _15858_);
  and (_16658_, _16657_, _15865_);
  or (_16659_, _16658_, _16655_);
  or (_16660_, _16659_, _16654_);
  nor (_16661_, _16660_, _16653_);
  nand (_16662_, _16661_, _15695_);
  or (_16663_, _16662_, _16652_);
  or (_16664_, _16663_, _16651_);
  and (_36899_[12], _16664_, _16644_);
  not (_16665_, _16401_);
  or (_16666_, _15809_, _15804_);
  nand (_16667_, _16646_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_16668_, _16667_, _16666_);
  nor (_16669_, _16668_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_16670_, _16668_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_16671_, _16670_, _16669_);
  and (_16672_, _16671_, _15830_);
  nor (_16673_, _14570_, _33470_);
  nor (_16674_, _15833_, _14602_);
  and (_16675_, _15836_, _16505_);
  and (_16676_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_16677_, _15858_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_16678_, _16677_, _15859_);
  and (_16679_, _16678_, _15865_);
  or (_16680_, _16679_, _16676_);
  or (_16681_, _16680_, _16675_);
  or (_16682_, _16681_, _16674_);
  or (_16683_, _16682_, _16673_);
  or (_16684_, _16683_, _16672_);
  or (_16685_, _16684_, _16665_);
  nor (_16686_, _15711_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_16687_, _16686_, _15712_);
  or (_16688_, _16687_, _16401_);
  and (_16689_, _16688_, _38997_);
  and (_36899_[13], _16689_, _16685_);
  and (_16690_, _14632_, _33469_);
  and (_16691_, _15826_, _14659_);
  and (_16692_, _15848_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_16693_, _15836_, _34686_);
  or (_16694_, _16693_, _16692_);
  or (_16695_, _15859_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_16696_, _16695_, _15860_);
  and (_16697_, _16696_, _15865_);
  or (_16698_, _16697_, _16694_);
  or (_16699_, _16698_, _16691_);
  or (_16700_, _16699_, _16690_);
  and (_16701_, _15811_, _15803_);
  nor (_16702_, _16701_, _14137_);
  and (_16703_, _16701_, _14137_);
  or (_16704_, _16703_, _16702_);
  and (_16705_, _16704_, _16411_);
  or (_16706_, _16705_, _16700_);
  or (_16707_, _16706_, _16665_);
  nor (_16708_, _15712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_16709_, _16708_, _15713_);
  or (_16710_, _16709_, _16401_);
  and (_16711_, _16710_, _38997_);
  and (_36899_[14], _16711_, _16707_);
  and (_16712_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_16713_, _16059_, _16057_);
  nor (_16714_, _16713_, _16060_);
  or (_16715_, _16714_, _15877_);
  or (_16716_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_16717_, _16716_, _16091_);
  and (_16718_, _16717_, _16715_);
  or (_36900_[0], _16718_, _16712_);
  and (_16719_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_16720_, _16062_, _16060_);
  and (_16721_, _16720_, _16063_);
  or (_16722_, _16721_, _15877_);
  or (_16723_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_16724_, _16723_, _16091_);
  and (_16725_, _16724_, _16722_);
  or (_36900_[1], _16725_, _16719_);
  and (_16726_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_16727_, _16067_, _16065_);
  nor (_16728_, _16727_, _16068_);
  or (_16729_, _16728_, _15877_);
  or (_16730_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_16731_, _16730_, _16091_);
  and (_16732_, _16731_, _16729_);
  or (_36900_[2], _16732_, _16726_);
  and (_16733_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_16734_, _16068_, _15952_);
  nor (_16735_, _16734_, _16069_);
  or (_16736_, _16735_, _15877_);
  or (_16737_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_16738_, _16737_, _16091_);
  and (_16739_, _16738_, _16736_);
  or (_36900_[3], _16739_, _16733_);
  nor (_16740_, _16072_, _16069_);
  nor (_16741_, _16740_, _16073_);
  or (_16742_, _16741_, _15877_);
  or (_16743_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_16744_, _16743_, _16091_);
  and (_16745_, _16744_, _16742_);
  and (_16746_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_36900_[4], _16746_, _16745_);
  nor (_16747_, _16073_, _15947_);
  nor (_16748_, _16747_, _16074_);
  or (_16749_, _16748_, _15877_);
  or (_16750_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_16751_, _16750_, _16091_);
  and (_16752_, _16751_, _16749_);
  and (_16753_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_36900_[5], _16753_, _16752_);
  nor (_16754_, _16074_, _15943_);
  nor (_16755_, _16754_, _16075_);
  or (_16756_, _16755_, _15877_);
  or (_16757_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_16758_, _16757_, _16091_);
  and (_16759_, _16758_, _16756_);
  and (_16760_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_36900_[6], _16760_, _16759_);
  and (_16761_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_16762_, _16075_, _15939_);
  nor (_16763_, _16762_, _16076_);
  or (_16764_, _16763_, _15877_);
  or (_16765_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_16766_, _16765_, _16091_);
  and (_16767_, _16766_, _16764_);
  or (_36900_[7], _16767_, _16761_);
  or (_16768_, _16078_, _16076_);
  nor (_16769_, _16079_, _15877_);
  and (_16770_, _16769_, _16768_);
  nor (_16771_, _15876_, _14110_);
  or (_16772_, _16771_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_16773_, _16772_, _16770_);
  or (_16774_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _33132_);
  and (_16775_, _16774_, _38997_);
  and (_36900_[8], _16775_, _16773_);
  nor (_16776_, _16079_, _15934_);
  nor (_16777_, _16776_, _16080_);
  or (_16778_, _16777_, _15877_);
  or (_16779_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_16780_, _16779_, _16091_);
  and (_16781_, _16780_, _16778_);
  and (_16782_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_36900_[9], _16782_, _16781_);
  nor (_16783_, _16080_, _15931_);
  nor (_16784_, _16783_, _16081_);
  or (_16785_, _16784_, _15877_);
  or (_16786_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_16787_, _16786_, _16091_);
  and (_16788_, _16787_, _16785_);
  and (_16789_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_36900_[10], _16789_, _16788_);
  and (_16790_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_16791_, _16081_, _15927_);
  nor (_16792_, _16791_, _16082_);
  or (_16793_, _16792_, _15877_);
  or (_16794_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_16795_, _16794_, _16091_);
  and (_16796_, _16795_, _16793_);
  or (_36900_[11], _16796_, _16790_);
  nor (_16797_, _16082_, _15923_);
  nor (_16798_, _16797_, _16083_);
  or (_16799_, _16798_, _15877_);
  or (_16800_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_16801_, _16800_, _16091_);
  and (_16802_, _16801_, _16799_);
  and (_16803_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_36900_[12], _16803_, _16802_);
  nor (_16804_, _16083_, _15920_);
  nor (_16805_, _16804_, _16084_);
  or (_16806_, _16805_, _15877_);
  or (_16807_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_16808_, _16807_, _16091_);
  and (_16809_, _16808_, _16806_);
  and (_16810_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_36900_[13], _16810_, _16809_);
  nor (_16811_, _16084_, _15917_);
  nor (_16812_, _16811_, _16085_);
  or (_16813_, _16812_, _15877_);
  or (_16814_, _15876_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_16815_, _16814_, _16091_);
  and (_16816_, _16815_, _16813_);
  and (_16817_, _15873_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_36900_[14], _16817_, _16816_);
  and (_16818_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_16819_, _16818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_36904_[0], _16819_, _38997_);
  and (_16820_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_16821_, _16820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_36904_[1], _16821_, _38997_);
  and (_16822_, _16102_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_16823_, _16822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_36904_[2], _16823_, _38997_);
  and (_16824_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_16825_, _16824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_36904_[3], _16825_, _38997_);
  and (_16826_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_16827_, _16826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_36904_[4], _16827_, _38997_);
  and (_16828_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_16829_, _16828_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_36904_[5], _16829_, _38997_);
  and (_16830_, _16103_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_16831_, _16830_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_36904_[6], _16831_, _38997_);
  nor (_16832_, _16056_, _34325_);
  nand (_16833_, _16832_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_16834_, _16832_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_16835_, _16834_, _16091_);
  and (_36905_[0], _16835_, _16833_);
  or (_16836_, _16115_, _16113_);
  and (_16837_, _16836_, _16116_);
  or (_16838_, _16837_, _34325_);
  or (_16839_, _33135_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_16840_, _16839_, _16091_);
  and (_36905_[1], _16840_, _16838_);
  and (_16841_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_16842_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_16843_, _16842_, _36910_);
  or (_36909_[0], _16843_, _16841_);
  and (_16844_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_16845_, _16298_, _36910_);
  or (_36909_[1], _16845_, _16844_);
  and (_16846_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_16847_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_16848_, _16847_, _36910_);
  or (_36909_[2], _16848_, _16846_);
  and (_16849_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_16850_, _16305_, _36910_);
  or (_36909_[3], _16850_, _16849_);
  and (_16851_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_16852_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_16853_, _16852_, _36910_);
  or (_36909_[4], _16853_, _16851_);
  and (_16854_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_16855_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_16856_, _16855_, _36910_);
  or (_36909_[5], _16856_, _16854_);
  and (_16857_, _16136_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_16858_, _16315_, _36910_);
  or (_36909_[6], _16858_, _16857_);
  and (_36912_[0], _16144_, _38997_);
  nor (_36912_[1], _16154_, rst);
  and (_36912_[2], _16150_, _38997_);
  or (_16859_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand (_16860_, _16158_, _15469_);
  and (_16861_, _16860_, _38997_);
  and (_36914_[0], _16861_, _16859_);
  and (_16862_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_16863_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_16864_, _16863_, _16862_);
  and (_36914_[1], _16864_, _38997_);
  or (_16865_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_16866_, _16158_, _15501_);
  and (_16867_, _16866_, _38997_);
  and (_36914_[2], _16867_, _16865_);
  or (_16868_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_16869_, _16158_, _15522_);
  and (_16870_, _16869_, _38997_);
  and (_36914_[3], _16870_, _16868_);
  or (_16871_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand (_16872_, _16158_, _15540_);
  and (_16873_, _16872_, _38997_);
  and (_36914_[4], _16873_, _16871_);
  or (_16874_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_16875_, _16158_, _15555_);
  and (_16876_, _16875_, _38997_);
  and (_36914_[5], _16876_, _16874_);
  or (_16877_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_16878_, _16158_, _15576_);
  and (_16879_, _16878_, _38997_);
  and (_36914_[6], _16879_, _16877_);
  or (_16880_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_16881_, _16158_, _15451_);
  and (_16882_, _16881_, _38997_);
  and (_36914_[7], _16882_, _16880_);
  and (_16883_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_16884_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_16885_, _16884_, _16883_);
  and (_36914_[8], _16885_, _38997_);
  and (_16886_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_16887_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_16888_, _16887_, _16886_);
  and (_36914_[9], _16888_, _38997_);
  and (_16889_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_16890_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_16891_, _16890_, _16889_);
  and (_36914_[10], _16891_, _38997_);
  and (_16892_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_16893_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_16894_, _16893_, _16892_);
  and (_36914_[11], _16894_, _38997_);
  and (_16895_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_16896_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_16897_, _16896_, _16895_);
  and (_36914_[12], _16897_, _38997_);
  and (_16898_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_16899_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_16900_, _16899_, _16898_);
  and (_36914_[13], _16900_, _38997_);
  and (_16901_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_16902_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_16903_, _16902_, _16901_);
  and (_36914_[14], _16903_, _38997_);
  and (_16904_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_16905_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_16906_, _16905_, _16904_);
  and (_36914_[15], _16906_, _38997_);
  and (_16907_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_16908_, _16158_, _33206_);
  or (_16909_, _16908_, _16907_);
  and (_36914_[16], _16909_, _38997_);
  and (_16910_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_16911_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_16912_, _16911_, _16910_);
  and (_36914_[17], _16912_, _38997_);
  and (_16913_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_16914_, _16158_, _33142_);
  or (_16915_, _16914_, _16913_);
  and (_36914_[18], _16915_, _38997_);
  and (_16916_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_16917_, _16158_, _33184_);
  or (_16918_, _16917_, _16916_);
  and (_36914_[19], _16918_, _38997_);
  and (_16919_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_16920_, _16158_, _33256_);
  or (_16921_, _16920_, _16919_);
  and (_36914_[20], _16921_, _38997_);
  and (_16922_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_16923_, _16158_, _33285_);
  or (_16924_, _16923_, _16922_);
  and (_36914_[21], _16924_, _38997_);
  and (_16925_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_16926_, _16158_, _33331_);
  or (_16927_, _16926_, _16925_);
  and (_36914_[22], _16927_, _38997_);
  and (_16928_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_16929_, _16158_, _33303_);
  or (_16930_, _16929_, _16928_);
  and (_36914_[23], _16930_, _38997_);
  and (_16931_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nor (_16932_, _16158_, _34445_);
  or (_16933_, _16932_, _16931_);
  and (_36914_[24], _16933_, _38997_);
  and (_16934_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_16935_, _16160_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_16936_, _16935_, _16934_);
  and (_36914_[25], _16936_, _38997_);
  and (_16937_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nor (_16938_, _16158_, _34747_);
  or (_16939_, _16938_, _16937_);
  and (_36914_[26], _16939_, _38997_);
  and (_16940_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nor (_16941_, _16158_, _34405_);
  or (_16942_, _16941_, _16940_);
  and (_36914_[27], _16942_, _38997_);
  and (_16943_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_16944_, _16158_, _34483_);
  or (_16945_, _16944_, _16943_);
  and (_36914_[28], _16945_, _38997_);
  and (_16946_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_16947_, _16158_, _34591_);
  or (_16948_, _16947_, _16946_);
  and (_36914_[29], _16948_, _38997_);
  and (_16949_, _16158_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_16950_, _16158_, _34673_);
  or (_16951_, _16950_, _16949_);
  and (_36914_[30], _16951_, _38997_);
  and (_16952_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16953_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_16954_, _16953_, _16952_);
  and (_36915_[0], _16954_, _38997_);
  and (_16955_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16956_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_16957_, _16956_, _16955_);
  and (_36915_[1], _16957_, _38997_);
  and (_16958_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16959_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_16960_, _16959_, _16958_);
  and (_36915_[2], _16960_, _38997_);
  and (_16961_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16962_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_16963_, _16962_, _16961_);
  and (_36915_[3], _16963_, _38997_);
  and (_16964_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16965_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_16966_, _16965_, _16964_);
  and (_36915_[4], _16966_, _38997_);
  and (_16967_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16968_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_16969_, _16968_, _16967_);
  and (_36915_[5], _16969_, _38997_);
  and (_16970_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_16971_, _16168_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_16972_, _16971_, _16970_);
  and (_36915_[6], _16972_, _38997_);
  and (_16973_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_16974_, _34441_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_16975_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_16976_, _16975_, _16167_);
  and (_16977_, _16976_, _16974_);
  or (_16978_, _16977_, _16973_);
  and (_36918_[0], _16978_, _38997_);
  and (_16979_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_16980_, _34548_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_16981_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_16982_, _16981_, _16167_);
  and (_16983_, _16982_, _16980_);
  or (_16984_, _16983_, _16979_);
  and (_36918_[1], _16984_, _38997_);
  and (_16985_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_16986_, _34741_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_16987_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_16988_, _16987_, _16167_);
  and (_16989_, _16988_, _16986_);
  or (_16990_, _16989_, _16985_);
  and (_36918_[2], _16990_, _38997_);
  and (_16991_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_16992_, _34391_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_16993_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_16994_, _16993_, _16167_);
  and (_16995_, _16994_, _16992_);
  or (_16996_, _16995_, _16991_);
  and (_36918_[3], _16996_, _38997_);
  and (_16997_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_16998_, _34517_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_16999_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_17000_, _16999_, _16167_);
  and (_17001_, _17000_, _16998_);
  or (_17002_, _17001_, _16997_);
  and (_36918_[4], _17002_, _38997_);
  and (_17003_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_17004_, _34634_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_17005_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_17006_, _17005_, _16167_);
  and (_17007_, _17006_, _17004_);
  or (_17008_, _17007_, _17003_);
  and (_36918_[5], _17008_, _38997_);
  and (_17009_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_17010_, _34669_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_17011_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_17012_, _17011_, _16167_);
  and (_17013_, _17012_, _17010_);
  or (_17014_, _17013_, _17009_);
  and (_36918_[6], _17014_, _38997_);
  and (_17015_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17016_, _34320_, _16174_);
  or (_17017_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_17018_, _17017_, _16167_);
  and (_17019_, _17018_, _17016_);
  or (_17020_, _17019_, _17015_);
  and (_36918_[7], _17020_, _38997_);
  and (_17021_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_17022_, _17021_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17023_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _16167_);
  and (_17024_, _17023_, _38997_);
  and (_36918_[8], _17024_, _17022_);
  and (_17025_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_17026_, _17025_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17027_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _16167_);
  and (_17028_, _17027_, _38997_);
  and (_36918_[9], _17028_, _17026_);
  and (_17029_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_17030_, _17029_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17031_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _16167_);
  and (_17032_, _17031_, _38997_);
  and (_36918_[10], _17032_, _17030_);
  and (_17033_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_17034_, _17033_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17035_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _16167_);
  and (_17036_, _17035_, _38997_);
  and (_36918_[11], _17036_, _17034_);
  and (_17037_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_17038_, _17037_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17039_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _16167_);
  and (_17040_, _17039_, _38997_);
  and (_36918_[12], _17040_, _17038_);
  and (_17041_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_17042_, _17041_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17043_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _16167_);
  and (_17044_, _17043_, _38997_);
  and (_36918_[13], _17044_, _17042_);
  and (_17045_, _16174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_17046_, _17045_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_17047_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _16167_);
  and (_17048_, _17047_, _38997_);
  and (_36918_[14], _17048_, _17046_);
  not (_17049_, _16181_);
  or (_17050_, _17049_, _14223_);
  or (_17051_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_17052_, _17051_, _38997_);
  and (_36922_[0], _17052_, _17050_);
  or (_17053_, _17049_, _14289_);
  or (_17054_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_17055_, _17054_, _38997_);
  and (_36922_[1], _17055_, _17053_);
  nand (_17056_, _16181_, _14356_);
  or (_17057_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_17058_, _17057_, _38997_);
  and (_36922_[2], _17058_, _17056_);
  nand (_17059_, _16181_, _14423_);
  or (_17060_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_17061_, _17060_, _38997_);
  and (_36922_[3], _17061_, _17059_);
  or (_17062_, _17049_, _14494_);
  or (_17063_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_17064_, _17063_, _38997_);
  and (_36922_[4], _17064_, _17062_);
  nand (_17065_, _16181_, _14570_);
  or (_17066_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_17067_, _17066_, _38997_);
  and (_36922_[5], _17067_, _17065_);
  or (_17068_, _17049_, _14632_);
  or (_17069_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_17070_, _17069_, _38997_);
  and (_36922_[6], _17070_, _17068_);
  nand (_17071_, _16181_, _14098_);
  or (_17072_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_17073_, _17072_, _38997_);
  and (_36922_[7], _17073_, _17071_);
  or (_17074_, _17049_, _14250_);
  or (_17075_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_17076_, _17075_, _38997_);
  and (_36922_[8], _17076_, _17074_);
  nand (_17077_, _16181_, _14323_);
  or (_17078_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_17079_, _17078_, _38997_);
  and (_36922_[9], _17079_, _17077_);
  nand (_17080_, _16181_, _14387_);
  or (_17081_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_17082_, _17081_, _38997_);
  and (_36922_[10], _17082_, _17080_);
  nand (_17083_, _16181_, _14456_);
  or (_17084_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_17085_, _17084_, _38997_);
  and (_36922_[11], _17085_, _17083_);
  nand (_17086_, _16181_, _14529_);
  or (_17087_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_17088_, _17087_, _38997_);
  and (_36922_[12], _17088_, _17086_);
  nand (_17089_, _16181_, _14602_);
  or (_17090_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_17091_, _17090_, _38997_);
  and (_36922_[13], _17091_, _17089_);
  or (_17092_, _17049_, _14659_);
  or (_17093_, _16181_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_17094_, _17093_, _38997_);
  and (_36922_[14], _17094_, _17092_);
  nor (_36880_, _34369_, rst);
  and (_17095_, _34258_, _34247_);
  nand (_17096_, _17095_, _34221_);
  or (_17097_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_17098_, _17097_, _38997_);
  and (_36881_[7], _17098_, _17096_);
  not (_17099_, _34260_);
  nor (_17100_, _17099_, _34221_);
  and (_17101_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_17102_, _17101_, _34248_);
  or (_17103_, _17102_, _17100_);
  or (_17104_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_17105_, _17104_, _38997_);
  and (_36882_[7], _17105_, _17103_);
  and (_17106_, _34263_, _34247_);
  not (_17107_, _17106_);
  nor (_17108_, _17107_, _34221_);
  and (_17109_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or (_17110_, _17109_, _17108_);
  and (_36883_[7], _17110_, _38997_);
  and (_17111_, _34255_, _34247_);
  not (_17112_, _17111_);
  nor (_17113_, _17112_, _34221_);
  and (_17114_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_17115_, _17114_, _17113_);
  and (_36884_[7], _17115_, _38997_);
  and (_17116_, _34268_, _34247_);
  not (_17117_, _17116_);
  nor (_17118_, _17117_, _34221_);
  and (_17119_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_17120_, _17119_, _17118_);
  and (_36885_[7], _17120_, _38997_);
  and (_17121_, _34269_, _34247_);
  and (_17122_, _17121_, _34318_);
  and (_17123_, _34270_, _34266_);
  nand (_17124_, _34261_, _34247_);
  or (_17125_, _17124_, _17123_);
  or (_17126_, _34255_, _34263_);
  or (_17127_, _34268_, _17126_);
  and (_17128_, _17127_, _34247_);
  or (_17129_, _17128_, _17125_);
  and (_17130_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or (_17131_, _17130_, _17122_);
  and (_36886_[7], _17131_, _38997_);
  and (_17132_, _34271_, _34247_);
  not (_17133_, _17132_);
  nor (_17134_, _17133_, _34221_);
  and (_17135_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or (_17136_, _17135_, _17134_);
  and (_36887_[7], _17136_, _38997_);
  not (_17137_, _34266_);
  or (_17138_, _34279_, _17137_);
  and (_17139_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_17140_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_17141_, _17140_, _34273_);
  nor (_17142_, _34278_, _34221_);
  or (_17143_, _17142_, _17141_);
  or (_17144_, _17143_, _17139_);
  and (_36888_[7], _17144_, _38997_);
  nand (_17145_, _17095_, _34148_);
  or (_17146_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_17147_, _17146_, _38997_);
  and (_36881_[0], _17147_, _17145_);
  not (_17148_, _17095_);
  or (_17149_, _17148_, _34122_);
  or (_17150_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_17151_, _17150_, _38997_);
  and (_36881_[1], _17151_, _17149_);
  or (_17152_, _17148_, _34089_);
  or (_17153_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_17154_, _17153_, _38997_);
  and (_36881_[2], _17154_, _17152_);
  nand (_17155_, _17095_, _34052_);
  or (_17156_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_17157_, _17156_, _38997_);
  and (_36881_[3], _17157_, _17155_);
  nand (_17158_, _17095_, _34017_);
  or (_17159_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_17160_, _17159_, _38997_);
  and (_36881_[4], _17160_, _17158_);
  or (_17161_, _17148_, _33978_);
  or (_17162_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_17163_, _17162_, _38997_);
  and (_36881_[5], _17163_, _17161_);
  or (_17164_, _17148_, _33942_);
  or (_17165_, _17095_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_17166_, _17165_, _38997_);
  and (_36881_[6], _17166_, _17164_);
  and (_17167_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_17168_, _34260_, _34149_);
  or (_17169_, _17168_, _34248_);
  or (_17170_, _17169_, _17167_);
  or (_17171_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_17172_, _17171_, _38997_);
  and (_36882_[0], _17172_, _17170_);
  and (_17173_, _34260_, _34122_);
  and (_17174_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_17175_, _17174_, _34248_);
  or (_17176_, _17175_, _17173_);
  or (_17177_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_17178_, _17177_, _38997_);
  and (_36882_[1], _17178_, _17176_);
  and (_17179_, _34260_, _34089_);
  and (_17180_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_17181_, _17180_, _34248_);
  or (_17182_, _17181_, _17179_);
  or (_17183_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_17184_, _17183_, _38997_);
  and (_36882_[2], _17184_, _17182_);
  nor (_17185_, _17099_, _34052_);
  and (_17186_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_17187_, _17186_, _34248_);
  or (_17188_, _17187_, _17185_);
  or (_17189_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_17190_, _17189_, _38997_);
  and (_36882_[3], _17190_, _17188_);
  nor (_17191_, _17099_, _34017_);
  and (_17192_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_17193_, _17192_, _34248_);
  or (_17194_, _17193_, _17191_);
  or (_17195_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_17196_, _17195_, _38997_);
  and (_36882_[4], _17196_, _17194_);
  and (_17197_, _34260_, _33978_);
  and (_17198_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_17199_, _17198_, _34248_);
  or (_17200_, _17199_, _17197_);
  or (_17201_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_17202_, _17201_, _38997_);
  and (_36882_[5], _17202_, _17200_);
  and (_17203_, _34260_, _33942_);
  and (_17204_, _17099_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_17205_, _17204_, _34248_);
  or (_17206_, _17205_, _17203_);
  or (_17207_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_17208_, _17207_, _38997_);
  and (_36882_[6], _17208_, _17206_);
  or (_17209_, _34265_, _34248_);
  and (_17210_, _17209_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand (_17211_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_17212_, _17211_, _34261_);
  and (_17213_, _17106_, _34149_);
  or (_17214_, _17213_, _17212_);
  or (_17215_, _17214_, _17210_);
  and (_36883_[0], _17215_, _38997_);
  and (_17216_, _17106_, _34122_);
  and (_17217_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_17218_, _17217_, _17216_);
  and (_36883_[1], _17218_, _38997_);
  and (_17219_, _17106_, _34089_);
  and (_17220_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_17221_, _17220_, _17219_);
  and (_36883_[2], _17221_, _38997_);
  nor (_17222_, _17107_, _34052_);
  and (_17223_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_17224_, _17223_, _17222_);
  and (_36883_[3], _17224_, _38997_);
  and (_17225_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_17226_, _17107_, _34017_);
  or (_17227_, _17226_, _17225_);
  and (_36883_[4], _17227_, _38997_);
  and (_17228_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_17229_, _17106_, _33978_);
  or (_17230_, _17229_, _17228_);
  and (_36883_[5], _17230_, _38997_);
  and (_17231_, _17106_, _33942_);
  and (_17232_, _17107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_17233_, _17232_, _17231_);
  and (_36883_[6], _17233_, _38997_);
  and (_17234_, _17111_, _34149_);
  and (_17235_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_17236_, _17235_, _17234_);
  and (_36884_[0], _17236_, _38997_);
  and (_17237_, _17111_, _34122_);
  and (_17238_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_17239_, _17238_, _17237_);
  and (_36884_[1], _17239_, _38997_);
  and (_17240_, _17111_, _34089_);
  and (_17241_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_17242_, _17241_, _17240_);
  and (_36884_[2], _17242_, _38997_);
  and (_17243_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_17244_, _17112_, _34052_);
  or (_17245_, _17244_, _17243_);
  and (_36884_[3], _17245_, _38997_);
  nor (_17246_, _17112_, _34017_);
  and (_17247_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_17248_, _17247_, _17246_);
  and (_36884_[4], _17248_, _38997_);
  and (_17249_, _17111_, _33978_);
  and (_17250_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_17251_, _17250_, _17249_);
  and (_36884_[5], _17251_, _38997_);
  and (_17252_, _17111_, _33942_);
  and (_17253_, _17112_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or (_17254_, _17253_, _17252_);
  and (_36884_[6], _17254_, _38997_);
  and (_17255_, _17116_, _34149_);
  and (_17256_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or (_17257_, _17256_, _17255_);
  and (_36885_[0], _17257_, _38997_);
  and (_17258_, _17116_, _34122_);
  and (_17259_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or (_17260_, _17259_, _17258_);
  and (_36885_[1], _17260_, _38997_);
  and (_17261_, _17116_, _34089_);
  and (_17262_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_17263_, _17262_, _17261_);
  and (_36885_[2], _17263_, _38997_);
  nor (_17264_, _17117_, _34052_);
  and (_17265_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_17266_, _17265_, _17264_);
  and (_36885_[3], _17266_, _38997_);
  nor (_17267_, _17117_, _34017_);
  and (_17268_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_17269_, _17268_, _17267_);
  and (_36885_[4], _17269_, _38997_);
  and (_17270_, _34268_, _33978_);
  and (_17271_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_17272_, _17271_, _17270_);
  or (_17273_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_17274_, _17273_, _38997_);
  and (_36885_[5], _17274_, _17272_);
  and (_17275_, _17117_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_17276_, _17116_, _33942_);
  or (_17277_, _17276_, _17275_);
  and (_36885_[6], _17277_, _38997_);
  and (_17278_, _17121_, _34149_);
  and (_17279_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or (_17280_, _17279_, _17278_);
  and (_36886_[0], _17280_, _38997_);
  or (_17281_, _17127_, _17125_);
  and (_17282_, _17281_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_17283_, _17121_, _34122_);
  or (_17284_, _17283_, _17282_);
  and (_36886_[1], _17284_, _38997_);
  and (_17285_, _17121_, _34089_);
  and (_17286_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or (_17287_, _17286_, _17285_);
  and (_36886_[2], _17287_, _38997_);
  and (_17288_, _17121_, _34389_);
  and (_17289_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_17290_, _17289_, _17288_);
  and (_36886_[3], _17290_, _38997_);
  and (_17291_, _17121_, _34515_);
  and (_17292_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or (_17293_, _17292_, _17291_);
  and (_36886_[4], _17293_, _38997_);
  and (_17294_, _17121_, _33978_);
  and (_17295_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or (_17296_, _17295_, _17294_);
  and (_36886_[5], _17296_, _38997_);
  and (_17297_, _17121_, _33942_);
  and (_17298_, _17129_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_17299_, _17298_, _17297_);
  and (_36886_[6], _17299_, _38997_);
  and (_17300_, _17132_, _34149_);
  and (_17301_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or (_17302_, _17301_, _17300_);
  and (_36887_[0], _17302_, _38997_);
  not (_17303_, _34265_);
  or (_17304_, _34275_, _17303_);
  and (_17305_, _17304_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand (_17306_, _34270_, _34256_);
  and (_17307_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_17308_, _17307_, _17306_);
  and (_17309_, _17132_, _34122_);
  or (_17310_, _17309_, _17308_);
  or (_17311_, _17310_, _17305_);
  and (_36887_[1], _17311_, _38997_);
  and (_17312_, _17132_, _34089_);
  and (_17313_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_17314_, _17313_, _17312_);
  and (_36887_[2], _17314_, _38997_);
  nor (_17315_, _17133_, _34052_);
  and (_17316_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_17317_, _17316_, _17315_);
  and (_36887_[3], _17317_, _38997_);
  nor (_17318_, _17133_, _34017_);
  and (_17319_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or (_17320_, _17319_, _17318_);
  and (_36887_[4], _17320_, _38997_);
  and (_17321_, _17132_, _33978_);
  and (_17322_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_17323_, _17322_, _17321_);
  and (_36887_[5], _17323_, _38997_);
  and (_17324_, _17133_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_17325_, _17132_, _33942_);
  or (_17326_, _17325_, _17324_);
  and (_36887_[6], _17326_, _38997_);
  and (_17327_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_17328_, _34267_, _34254_);
  and (_17329_, _17328_, _34149_);
  not (_17330_, _34273_);
  and (_17331_, _17330_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_17332_, _17331_, _17329_);
  and (_17333_, _17332_, _34247_);
  or (_17334_, _17333_, _17327_);
  and (_36888_[0], _17334_, _38997_);
  and (_17335_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_17336_, _17328_, _34122_);
  and (_17337_, _17330_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or (_17338_, _17337_, _17336_);
  and (_17339_, _17338_, _34247_);
  or (_17340_, _17339_, _17335_);
  and (_36888_[1], _17340_, _38997_);
  and (_17341_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nand (_17342_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_17343_, _17342_, _34273_);
  and (_17344_, _34277_, _34089_);
  or (_17345_, _17344_, _17343_);
  or (_17346_, _17345_, _17341_);
  and (_36888_[2], _17346_, _38997_);
  and (_17347_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nand (_17348_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_17349_, _17348_, _34273_);
  nor (_17350_, _34278_, _34052_);
  or (_17351_, _17350_, _17349_);
  or (_17352_, _17351_, _17347_);
  and (_36888_[3], _17352_, _38997_);
  and (_17353_, _17138_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nand (_17354_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_17355_, _17354_, _34273_);
  nor (_17356_, _34278_, _34017_);
  or (_17357_, _17356_, _17355_);
  or (_17358_, _17357_, _17353_);
  and (_36888_[4], _17358_, _38997_);
  and (_17359_, _34279_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_17360_, _34277_, _33978_);
  nand (_17361_, _34247_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_17362_, _17361_, _34274_);
  or (_17363_, _17362_, _17360_);
  or (_17364_, _17363_, _17359_);
  and (_36888_[5], _17364_, _38997_);
  and (_17365_, _34277_, _33942_);
  and (_17366_, _34278_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_17367_, _17366_, _17365_);
  and (_36888_[6], _17367_, _38997_);
  not (_17368_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_17369_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_17370_, _17369_, _17368_);
  and (_17371_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _38997_);
  and (_38985_, _17371_, _17370_);
  nor (_17372_, _17370_, rst);
  nand (_17373_, _17369_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_17374_, _17369_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_17375_, _17374_, _17373_);
  and (_38986_[3], _17375_, _17372_);
  not (_17376_, _34691_);
  and (_17377_, _34637_, _17376_);
  and (_17378_, _34421_, _34346_);
  and (_17379_, _17378_, _34699_);
  and (_17380_, _17379_, _17377_);
  not (_17381_, _34770_);
  nand (_17382_, _14846_, _14832_);
  or (_17383_, _14846_, _14832_);
  nand (_17384_, _17383_, _17382_);
  or (_17385_, _14869_, _14858_);
  nand (_17386_, _14869_, _14858_);
  nand (_17387_, _17386_, _17385_);
  nand (_17388_, _17387_, _17384_);
  or (_17389_, _17387_, _17384_);
  nand (_17390_, _17389_, _17388_);
  or (_17391_, _14894_, _14882_);
  nand (_17392_, _14894_, _14882_);
  nand (_17393_, _17392_, _17391_);
  or (_17394_, _14904_, _14815_);
  nand (_17395_, _14904_, _14815_);
  and (_17396_, _17395_, _17394_);
  nand (_17397_, _17396_, _17393_);
  or (_17398_, _17396_, _17393_);
  nand (_17399_, _17398_, _17397_);
  nand (_17400_, _17399_, _17390_);
  or (_17401_, _17399_, _17390_);
  and (_17402_, _17401_, _17400_);
  or (_17403_, _17402_, _17381_);
  and (_17404_, _34579_, _34471_);
  or (_17405_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_17406_, _17405_, _17404_);
  and (_17407_, _17406_, _17403_);
  not (_17408_, _34579_);
  nor (_17409_, _17408_, _34471_);
  and (_17410_, _17409_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_17411_, _17408_, _34471_);
  and (_17412_, _17411_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_17413_, _17412_, _17410_);
  and (_17414_, _17413_, _17381_);
  nor (_17415_, _34579_, _34471_);
  nor (_17416_, _34770_, _13513_);
  and (_17417_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_17418_, _17417_, _17416_);
  and (_17419_, _17418_, _17415_);
  and (_17420_, _17409_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_17421_, _17411_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_17422_, _17421_, _17420_);
  and (_17423_, _17422_, _34770_);
  or (_17424_, _17423_, _17419_);
  or (_17425_, _17424_, _17414_);
  or (_17426_, _17425_, _17407_);
  and (_17427_, _17426_, _17380_);
  not (_17428_, _34421_);
  nor (_17429_, _34637_, _17376_);
  nor (_17430_, _34770_, _12205_);
  and (_17431_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_17432_, _17431_, _17430_);
  and (_17433_, _17432_, _17409_);
  and (_17434_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_17435_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_17436_, _17435_, _17434_);
  and (_17437_, _17436_, _17411_);
  nor (_17438_, _34770_, _12203_);
  and (_17439_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_17440_, _17439_, _17438_);
  and (_17441_, _17440_, _17404_);
  or (_17442_, _17441_, _17437_);
  and (_17443_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_17444_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_17445_, _17444_, _17443_);
  and (_17446_, _17445_, _17415_);
  or (_17447_, _17446_, _17442_);
  or (_17448_, _17447_, _17433_);
  and (_17449_, _34699_, _34346_);
  and (_17450_, _17449_, _17448_);
  and (_17451_, _34529_, _34346_);
  and (_17452_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_17453_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_17454_, _17453_, _17452_);
  and (_17455_, _17454_, _17415_);
  and (_17456_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_17457_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_17458_, _17457_, _17456_);
  and (_17459_, _17458_, _17411_);
  nor (_17460_, _34770_, _12174_);
  and (_17461_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_17462_, _17461_, _17460_);
  and (_17463_, _17462_, _17404_);
  or (_17464_, _17463_, _17459_);
  nor (_17465_, _34770_, _12178_);
  and (_17466_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_17467_, _17466_, _17465_);
  and (_17468_, _17467_, _17409_);
  or (_17469_, _17468_, _17464_);
  or (_17470_, _17469_, _17455_);
  and (_17471_, _17470_, _17451_);
  or (_17472_, _17471_, _17450_);
  and (_17473_, _17472_, _17429_);
  and (_17474_, _34637_, _34691_);
  nor (_17475_, _34770_, _11307_);
  and (_17476_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_17477_, _17476_, _17475_);
  and (_17478_, _17477_, _17409_);
  nor (_17479_, _34770_, _10903_);
  and (_17480_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_17481_, _17480_, _17479_);
  and (_17482_, _17481_, _17411_);
  nor (_17483_, _34770_, _10920_);
  and (_17484_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_17485_, _17484_, _17483_);
  and (_17486_, _17485_, _17404_);
  or (_17487_, _17486_, _17482_);
  nor (_17488_, _34770_, _11281_);
  and (_17489_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_17490_, _17489_, _17488_);
  and (_17491_, _17490_, _17415_);
  or (_17492_, _17491_, _17487_);
  or (_17493_, _17492_, _17478_);
  and (_17494_, _17493_, _17449_);
  nor (_17495_, _34770_, _11404_);
  and (_17496_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_17497_, _17496_, _17495_);
  and (_17498_, _17497_, _17411_);
  nor (_17499_, _34770_, _11494_);
  and (_17500_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_17501_, _17500_, _17499_);
  and (_17502_, _17501_, _17404_);
  or (_17503_, _17502_, _17498_);
  and (_17504_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_17505_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_17506_, _17505_, _17504_);
  and (_17507_, _17506_, _17415_);
  and (_17508_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_17509_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_17510_, _17509_, _17508_);
  and (_17511_, _17510_, _17409_);
  or (_17512_, _17511_, _17507_);
  or (_17513_, _17512_, _17503_);
  and (_17514_, _17513_, _17451_);
  or (_17515_, _17514_, _17494_);
  and (_17516_, _17515_, _17474_);
  or (_17517_, _17516_, _17473_);
  and (_17518_, _17517_, _17428_);
  and (_17519_, _17451_, _34421_);
  not (_17520_, _34355_);
  not (_17521_, _33433_);
  and (_17522_, _33201_, _33381_);
  nor (_17523_, _17522_, _33396_);
  and (_17524_, _17523_, _17521_);
  and (_17525_, _17524_, _17520_);
  and (_17526_, _17525_, _15407_);
  nor (_17527_, _33348_, _33323_);
  and (_17528_, _33515_, _17527_);
  or (_17529_, _15124_, _33430_);
  or (_17530_, _17529_, _17528_);
  nor (_17531_, _17530_, _15061_);
  and (_17532_, _17531_, _15400_);
  and (_17533_, _17532_, _17526_);
  and (_17534_, _17533_, _33428_);
  nor (_17535_, _17534_, _33477_);
  or (_17536_, _17535_, p0_in[4]);
  not (_17537_, _17535_);
  or (_17538_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_17539_, _17538_, _17536_);
  and (_17540_, _17539_, _17381_);
  or (_17541_, _17535_, p0_in[0]);
  or (_17542_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_17543_, _17542_, _17541_);
  and (_17544_, _17543_, _34770_);
  or (_17545_, _17544_, _17540_);
  and (_17546_, _17545_, _17404_);
  or (_17547_, _17535_, p0_in[7]);
  or (_17548_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_17549_, _17548_, _17547_);
  and (_17550_, _17549_, _17381_);
  or (_17551_, _17535_, p0_in[3]);
  or (_17552_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_17553_, _17552_, _17551_);
  and (_17554_, _17553_, _34770_);
  or (_17555_, _17554_, _17550_);
  and (_17556_, _17555_, _17415_);
  or (_17557_, _17556_, _17546_);
  or (_17558_, _17535_, p0_in[5]);
  or (_17559_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_17560_, _17559_, _17558_);
  and (_17561_, _17560_, _17381_);
  or (_17562_, _17535_, p0_in[1]);
  or (_17563_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_17564_, _17563_, _17562_);
  and (_17565_, _17564_, _34770_);
  or (_17566_, _17565_, _17561_);
  and (_17567_, _17566_, _17409_);
  nor (_17568_, _17535_, p0_in[6]);
  and (_17569_, _17535_, _13246_);
  nor (_17570_, _17569_, _17568_);
  and (_17571_, _17570_, _17381_);
  or (_17572_, _17535_, p0_in[2]);
  nand (_17573_, _17535_, _13190_);
  and (_17574_, _17573_, _17572_);
  and (_17575_, _17574_, _34770_);
  or (_17576_, _17575_, _17571_);
  and (_17577_, _17576_, _17411_);
  or (_17578_, _17577_, _17567_);
  or (_17579_, _17578_, _17557_);
  and (_17580_, _17579_, _17519_);
  or (_17581_, _17535_, p1_in[4]);
  or (_17582_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_17583_, _17582_, _17581_);
  and (_17584_, _17583_, _17381_);
  or (_17585_, _17535_, p1_in[0]);
  or (_17586_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_17587_, _17586_, _17585_);
  and (_17588_, _17587_, _34770_);
  or (_17589_, _17588_, _17584_);
  and (_17590_, _17589_, _17404_);
  or (_17591_, _17535_, p1_in[7]);
  or (_17592_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_17593_, _17592_, _17591_);
  and (_17594_, _17593_, _17381_);
  or (_17595_, _17535_, p1_in[3]);
  or (_17596_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_17597_, _17596_, _17595_);
  and (_17598_, _17597_, _34770_);
  or (_17599_, _17598_, _17594_);
  and (_17600_, _17599_, _17415_);
  or (_17601_, _17600_, _17590_);
  or (_17602_, _17535_, p1_in[5]);
  or (_17603_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_17604_, _17603_, _17602_);
  and (_17605_, _17604_, _17381_);
  or (_17606_, _17535_, p1_in[1]);
  or (_17607_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_17608_, _17607_, _17606_);
  and (_17609_, _17608_, _34770_);
  or (_17610_, _17609_, _17605_);
  and (_17611_, _17610_, _17409_);
  nor (_17612_, _17535_, p1_in[6]);
  and (_17613_, _17535_, _13330_);
  nor (_17614_, _17613_, _17612_);
  and (_17615_, _17614_, _17381_);
  or (_17616_, _17535_, p1_in[2]);
  or (_17617_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_17618_, _17617_, _17616_);
  and (_17619_, _17618_, _34770_);
  or (_17620_, _17619_, _17615_);
  and (_17621_, _17620_, _17411_);
  or (_17622_, _17621_, _17611_);
  or (_17623_, _17622_, _17601_);
  and (_17624_, _17623_, _17379_);
  or (_17625_, _17624_, _17580_);
  and (_17626_, _17625_, _17474_);
  nor (_17627_, _34637_, _34691_);
  nor (_17628_, _34770_, _14686_);
  and (_17629_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_17630_, _17629_, _17628_);
  and (_17631_, _17630_, _17415_);
  nor (_17632_, _34770_, _14782_);
  and (_17633_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_17634_, _17633_, _17632_);
  and (_17635_, _17634_, _17411_);
  nor (_17636_, _34770_, _14755_);
  and (_17637_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_17638_, _17637_, _17636_);
  and (_17639_, _17638_, _17404_);
  or (_17640_, _17639_, _17635_);
  nor (_17641_, _34770_, _14769_);
  and (_17642_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_17643_, _17642_, _17641_);
  and (_17644_, _17643_, _17409_);
  or (_17645_, _17644_, _17640_);
  or (_17646_, _17645_, _17631_);
  and (_17647_, _17646_, _17627_);
  or (_17648_, _17535_, p3_in[7]);
  or (_17649_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_17650_, _17649_, _17648_);
  and (_17651_, _17650_, _17381_);
  or (_17652_, _17535_, p3_in[3]);
  or (_17653_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_17654_, _17653_, _17652_);
  and (_17655_, _17654_, _34770_);
  or (_17656_, _17655_, _17651_);
  and (_17657_, _17656_, _17415_);
  nor (_17658_, _17535_, p3_in[6]);
  and (_17659_, _17535_, _13500_);
  nor (_17660_, _17659_, _17658_);
  and (_17661_, _17660_, _17381_);
  or (_17662_, _17535_, p3_in[2]);
  or (_17663_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_17664_, _17663_, _17662_);
  and (_17665_, _17664_, _34770_);
  or (_17666_, _17665_, _17661_);
  and (_17667_, _17666_, _17411_);
  or (_17668_, _17667_, _17657_);
  or (_17669_, _17535_, p3_in[4]);
  or (_17670_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_17671_, _17670_, _17669_);
  and (_17672_, _17671_, _17381_);
  or (_17673_, _17535_, p3_in[0]);
  or (_17674_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_17675_, _17674_, _17673_);
  and (_17676_, _17675_, _34770_);
  or (_17677_, _17676_, _17672_);
  and (_17678_, _17677_, _17404_);
  or (_17679_, _17535_, p3_in[5]);
  or (_17680_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_17681_, _17680_, _17679_);
  and (_17682_, _17681_, _17381_);
  or (_17683_, _17535_, p3_in[1]);
  or (_17684_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_17685_, _17684_, _17683_);
  and (_17686_, _17685_, _34770_);
  or (_17687_, _17686_, _17682_);
  and (_17688_, _17687_, _17409_);
  or (_17689_, _17688_, _17678_);
  or (_17690_, _17689_, _17668_);
  and (_17691_, _17690_, _17429_);
  or (_17692_, _17691_, _17647_);
  and (_17693_, _17692_, _17379_);
  and (_17694_, _15621_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_17695_, _17451_, _17377_);
  and (_17696_, _17695_, _17428_);
  nand (_17697_, _34691_, _34346_);
  or (_17698_, _17697_, _34421_);
  nand (_17699_, _17698_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nand (_17700_, _34529_, _34637_);
  or (_17701_, _17700_, _34691_);
  and (_17702_, _17701_, _17378_);
  or (_17703_, _17702_, _17699_);
  nor (_17704_, _17703_, _17696_);
  and (_17705_, _17627_, _17519_);
  nor (_17706_, _34770_, _33984_);
  and (_17707_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_17708_, _17707_, _17706_);
  and (_17709_, _17708_, _17404_);
  nor (_17710_, _34770_, _34193_);
  and (_17711_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_17712_, _17711_, _17710_);
  and (_17713_, _17712_, _17415_);
  or (_17714_, _17713_, _17709_);
  nor (_17715_, _34770_, _33773_);
  and (_17716_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_17717_, _17716_, _17715_);
  and (_17718_, _17717_, _17411_);
  nor (_17719_, _34770_, _33948_);
  and (_17720_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_17721_, _17720_, _17719_);
  and (_17722_, _17721_, _17409_);
  or (_17723_, _17722_, _17718_);
  or (_17724_, _17723_, _17714_);
  and (_17725_, _17724_, _17705_);
  or (_17726_, _17725_, _17704_);
  nor (_17727_, _34770_, _13097_);
  and (_17728_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_17729_, _17728_, _17727_);
  and (_17730_, _17729_, _17411_);
  nor (_17731_, _34770_, _11000_);
  and (_17732_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_17733_, _17732_, _17731_);
  and (_17734_, _17733_, _17404_);
  or (_17735_, _17734_, _17730_);
  and (_17736_, _17381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_17737_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_17738_, _17737_, _17736_);
  and (_17739_, _17738_, _17415_);
  nor (_17740_, _34770_, _10900_);
  and (_17741_, _34770_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_17742_, _17741_, _17740_);
  and (_17743_, _17742_, _17409_);
  or (_17744_, _17743_, _17739_);
  or (_17745_, _17744_, _17735_);
  and (_17746_, _17745_, _17696_);
  and (_17747_, _17519_, _17429_);
  or (_17748_, _17535_, p2_in[7]);
  or (_17749_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_17750_, _17749_, _17748_);
  and (_17751_, _17750_, _17381_);
  or (_17752_, _17535_, p2_in[3]);
  or (_17753_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_17754_, _17753_, _17752_);
  and (_17755_, _17754_, _34770_);
  or (_17756_, _17755_, _17751_);
  and (_17757_, _17756_, _17415_);
  or (_17758_, _17535_, p2_in[5]);
  or (_17759_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_17760_, _17759_, _17758_);
  and (_17761_, _17760_, _17381_);
  or (_17762_, _17535_, p2_in[1]);
  or (_17763_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_17764_, _17763_, _17762_);
  and (_17765_, _17764_, _34770_);
  or (_17766_, _17765_, _17761_);
  and (_17767_, _17766_, _17409_);
  or (_17768_, _17767_, _17757_);
  or (_17769_, _17535_, p2_in[4]);
  or (_17770_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_17771_, _17770_, _17769_);
  and (_17772_, _17771_, _17381_);
  or (_17773_, _17535_, p2_in[0]);
  or (_17774_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_17775_, _17774_, _17773_);
  and (_17776_, _17775_, _34770_);
  or (_17777_, _17776_, _17772_);
  and (_17778_, _17777_, _17404_);
  nor (_17779_, _17535_, p2_in[6]);
  and (_17780_, _17535_, _13415_);
  nor (_17781_, _17780_, _17779_);
  and (_17782_, _17781_, _17381_);
  or (_17783_, _17535_, p2_in[2]);
  or (_17784_, _17537_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_17785_, _17784_, _17783_);
  and (_17786_, _17785_, _34770_);
  or (_17787_, _17786_, _17782_);
  and (_17788_, _17787_, _17411_);
  or (_17789_, _17788_, _17778_);
  or (_17790_, _17789_, _17768_);
  and (_17791_, _17790_, _17747_);
  or (_17792_, _17791_, _17746_);
  or (_17793_, _17792_, _17726_);
  or (_17794_, _17793_, _17694_);
  or (_17795_, _17794_, _17693_);
  or (_17796_, _17795_, _17626_);
  or (_17797_, _17796_, _17518_);
  or (_17798_, _17797_, _17427_);
  and (_17799_, _17705_, _14795_);
  nor (_17800_, _17799_, _15630_);
  nand (_17801_, _17694_, _35722_);
  and (_17802_, _17801_, _17800_);
  and (_17803_, _17802_, _17798_);
  nor (_17804_, _34770_, _34221_);
  and (_17805_, _34770_, _34389_);
  or (_17806_, _17805_, _17804_);
  and (_17807_, _17806_, _17415_);
  and (_17808_, _17381_, _33942_);
  and (_17809_, _34770_, _34089_);
  or (_17810_, _17809_, _17808_);
  and (_17811_, _17810_, _17411_);
  nor (_17812_, _34770_, _34017_);
  and (_17813_, _34770_, _34149_);
  or (_17814_, _17813_, _17812_);
  and (_17815_, _17814_, _17404_);
  or (_17816_, _17815_, _17811_);
  and (_17817_, _17381_, _33978_);
  and (_17818_, _34770_, _34122_);
  or (_17819_, _17818_, _17817_);
  and (_17820_, _17819_, _17409_);
  or (_17821_, _17820_, _17816_);
  nor (_17822_, _17821_, _17807_);
  nor (_17823_, _17822_, _17800_);
  or (_17824_, _17823_, _17803_);
  and (_38987_, _17824_, _38997_);
  and (_17825_, _34770_, _34421_);
  and (_17826_, _17474_, _17451_);
  and (_17827_, _17826_, _17415_);
  and (_17828_, _17827_, _17825_);
  and (_17829_, _17828_, _14101_);
  and (_17830_, _34699_, _34637_);
  nor (_17831_, _34691_, _35178_);
  and (_17832_, _17825_, _17404_);
  and (_17833_, _17832_, _17831_);
  and (_17834_, _17833_, _17830_);
  and (_17835_, _17834_, _13518_);
  nor (_17836_, _17835_, _17829_);
  nor (_17837_, _17836_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_17838_, _17837_);
  not (_17839_, _11084_);
  and (_17840_, _17415_, _17381_);
  nor (_17841_, _17840_, _17839_);
  and (_17842_, _17841_, _15608_);
  nor (_17843_, _34699_, _34637_);
  and (_17844_, _17843_, _17833_);
  and (_17845_, _17844_, _14819_);
  nor (_17846_, _17845_, _17842_);
  and (_17847_, _17846_, _15624_);
  and (_17848_, _17847_, _17838_);
  and (_17849_, _17825_, _17411_);
  and (_17850_, _17849_, _17826_);
  and (_17851_, _17850_, _14101_);
  or (_17852_, _17851_, rst);
  nor (_38988_, _17852_, _17848_);
  and (_17853_, _34770_, _17428_);
  and (_17854_, _17853_, _17404_);
  and (_17855_, _17854_, _17826_);
  and (_17856_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_17857_, _17853_, _17415_);
  and (_17858_, _17857_, _17695_);
  and (_17859_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_17860_, _17859_, _17856_);
  and (_17861_, _17840_, _34421_);
  and (_17862_, _17449_, _17429_);
  and (_17863_, _17862_, _17861_);
  and (_17864_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_17865_, _17451_, _17429_);
  and (_17866_, _17865_, _17854_);
  and (_17867_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_17868_, _17867_, _17864_);
  or (_17869_, _17868_, _17860_);
  and (_17870_, _17854_, _17695_);
  and (_17871_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_17872_, _34770_, _34421_);
  and (_17873_, _17872_, _17404_);
  and (_17874_, _17873_, _17695_);
  and (_17875_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_17876_, _17875_, _17871_);
  and (_17877_, _17872_, _17409_);
  and (_17878_, _17877_, _17695_);
  and (_17879_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_17880_, _17853_, _17411_);
  and (_17881_, _17880_, _17695_);
  and (_17882_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_17883_, _17882_, _17879_);
  or (_17884_, _17883_, _17876_);
  or (_17885_, _17884_, _17869_);
  and (_17886_, _17857_, _17826_);
  and (_17887_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_17888_, _17853_, _17409_);
  and (_17889_, _17888_, _17826_);
  and (_17890_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_17891_, _17890_, _17887_);
  and (_17892_, _17877_, _17826_);
  and (_17893_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_17894_, _17880_, _17826_);
  and (_17895_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_17896_, _17895_, _17893_);
  or (_17897_, _17896_, _17891_);
  and (_17898_, _17474_, _17449_);
  and (_17899_, _17898_, _17854_);
  and (_17900_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_17901_, _17888_, _17898_);
  and (_17902_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_17903_, _17902_, _17900_);
  and (_17904_, _17873_, _17826_);
  and (_17905_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_17906_, _17861_, _17826_);
  and (_17907_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_17908_, _17907_, _17905_);
  or (_17909_, _17908_, _17903_);
  or (_17910_, _17909_, _17897_);
  or (_17911_, _17910_, _17885_);
  and (_17912_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_17913_, _17825_, _17415_);
  and (_17914_, _17913_, _17826_);
  and (_17915_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_17916_, _17915_, _17912_);
  and (_17917_, _17627_, _17449_);
  and (_17918_, _17917_, _17832_);
  and (_17919_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_17920_, _17825_, _17409_);
  and (_17921_, _17920_, _17826_);
  and (_17922_, _17921_, _34223_);
  or (_17923_, _17922_, _17919_);
  or (_17924_, _17923_, _17916_);
  and (_17925_, _17865_, _17832_);
  and (_17926_, _17925_, _17750_);
  and (_17927_, _17862_, _17832_);
  and (_17928_, _17927_, _17650_);
  or (_17929_, _17928_, _17926_);
  and (_17930_, _17832_, _17826_);
  and (_17931_, _17930_, _17549_);
  and (_17932_, _17898_, _17832_);
  and (_17933_, _17932_, _17593_);
  or (_17934_, _17933_, _17931_);
  or (_17935_, _17934_, _17929_);
  or (_17936_, _17935_, _17924_);
  and (_17937_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_17938_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_17939_, _17938_, _17937_);
  or (_17940_, _17939_, _17936_);
  or (_17941_, _17940_, _17911_);
  and (_17942_, _17941_, _17848_);
  nor (_17943_, _17881_, _17878_);
  nand (_17944_, _17696_, _17404_);
  and (_17945_, _17944_, _17943_);
  nor (_17946_, _17858_, _17855_);
  nor (_17947_, _17866_, _17863_);
  and (_17948_, _17947_, _17946_);
  and (_17949_, _17948_, _17945_);
  nor (_17950_, _17889_, _17886_);
  nor (_17951_, _17894_, _17892_);
  and (_17952_, _17951_, _17950_);
  nor (_17953_, _17906_, _17904_);
  nor (_17954_, _17901_, _17899_);
  and (_17955_, _17954_, _17953_);
  and (_17956_, _17955_, _17952_);
  and (_17957_, _17956_, _17949_);
  not (_17958_, _17832_);
  or (_17959_, _17958_, _17697_);
  nor (_17960_, _17914_, _17850_);
  nor (_17961_, _17921_, _17918_);
  and (_17962_, _17961_, _17960_);
  and (_17963_, _17962_, _17959_);
  nor (_17964_, _17844_, _17834_);
  and (_17965_, _17964_, _17963_);
  nand (_17966_, _17965_, _17957_);
  nand (_17967_, _17966_, _17848_);
  and (_17968_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_17969_, _17968_, _17942_);
  or (_17970_, _17969_, _17851_);
  nand (_17971_, _17851_, _14098_);
  and (_17972_, _17971_, _38997_);
  and (_38989_[7], _17972_, _17970_);
  nor (_38986_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_17973_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_17974_, _17369_, rst);
  and (_38986_[1], _17974_, _17973_);
  nor (_17975_, _17369_, _17368_);
  or (_17976_, _17975_, _17370_);
  and (_17977_, _17373_, _38997_);
  and (_38986_[2], _17977_, _17976_);
  and (_17978_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_17979_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_17980_, _17979_, _17978_);
  and (_17981_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_17982_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_17983_, _17982_, _17981_);
  or (_17984_, _17983_, _17980_);
  and (_17985_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_17986_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_17987_, _17986_, _17985_);
  and (_17988_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_17989_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_17990_, _17989_, _17988_);
  or (_17991_, _17990_, _17987_);
  or (_17992_, _17991_, _17984_);
  and (_17993_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_17994_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_17995_, _17994_, _17993_);
  and (_17996_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_17997_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_17998_, _17997_, _17996_);
  or (_17999_, _17998_, _17995_);
  and (_18000_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_18001_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_18002_, _18001_, _18000_);
  and (_18003_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_18004_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_18005_, _18004_, _18003_);
  or (_18006_, _18005_, _18002_);
  or (_18007_, _18006_, _17999_);
  or (_18008_, _18007_, _17992_);
  and (_18009_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_18010_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_18011_, _18010_, _18009_);
  and (_18012_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_18013_, _17921_);
  nor (_18014_, _18013_, _34466_);
  or (_18015_, _18014_, _18012_);
  or (_18016_, _18015_, _18011_);
  and (_18017_, _17927_, _17675_);
  and (_18018_, _17925_, _17775_);
  or (_18019_, _18018_, _18017_);
  and (_18020_, _17930_, _17543_);
  and (_18021_, _17932_, _17587_);
  or (_18022_, _18021_, _18020_);
  or (_18023_, _18022_, _18019_);
  or (_18024_, _18023_, _18016_);
  and (_18025_, _17834_, _17402_);
  and (_18026_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_18027_, _18026_, _18025_);
  or (_18028_, _18027_, _18024_);
  or (_18029_, _18028_, _18008_);
  and (_18030_, _18029_, _17848_);
  and (_18031_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_18032_, _18031_, _17851_);
  or (_18033_, _18032_, _18030_);
  nand (_18034_, _17851_, _14224_);
  and (_18035_, _18034_, _38997_);
  and (_38989_[0], _18035_, _18033_);
  and (_18036_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  not (_18037_, _17851_);
  and (_18038_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_18039_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_18040_, _18039_, _18038_);
  and (_18041_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_18042_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_18043_, _18042_, _18041_);
  or (_18044_, _18043_, _18040_);
  and (_18045_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_18046_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_18047_, _18046_, _18045_);
  and (_18048_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_18049_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_18050_, _18049_, _18048_);
  or (_18051_, _18050_, _18047_);
  or (_18052_, _18051_, _18044_);
  and (_18053_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_18054_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_18055_, _18054_, _18053_);
  and (_18056_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_18057_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_18058_, _18057_, _18056_);
  or (_18059_, _18058_, _18055_);
  and (_18060_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_18061_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_18062_, _18061_, _18060_);
  and (_18063_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_18064_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_18065_, _18064_, _18063_);
  or (_18066_, _18065_, _18062_);
  or (_18067_, _18066_, _18059_);
  or (_18068_, _18067_, _18052_);
  and (_18069_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_18070_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_18071_, _18070_, _18069_);
  and (_18072_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18073_, _17921_, _34558_);
  or (_18074_, _18073_, _18072_);
  or (_18075_, _18074_, _18071_);
  and (_18076_, _17932_, _17608_);
  and (_18077_, _17930_, _17564_);
  or (_18078_, _18077_, _18076_);
  and (_18079_, _17927_, _17685_);
  and (_18080_, _17925_, _17764_);
  or (_18081_, _18080_, _18079_);
  or (_18082_, _18081_, _18078_);
  or (_18083_, _18082_, _18075_);
  and (_18084_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_18085_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_18086_, _18085_, _18084_);
  or (_18087_, _18086_, _18083_);
  or (_18088_, _18087_, _18068_);
  nand (_18089_, _18088_, _17848_);
  nand (_18090_, _18089_, _18037_);
  or (_18091_, _18090_, _18036_);
  nand (_18092_, _17851_, _14290_);
  and (_18093_, _18092_, _38997_);
  and (_38989_[1], _18093_, _18091_);
  and (_18094_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_18095_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_18096_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_18097_, _18096_, _18095_);
  and (_18098_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_18099_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_18100_, _18099_, _18098_);
  or (_18101_, _18100_, _18097_);
  and (_18102_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_18103_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_18104_, _18103_, _18102_);
  and (_18105_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_18106_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_18107_, _18106_, _18105_);
  or (_18108_, _18107_, _18104_);
  or (_18109_, _18108_, _18101_);
  and (_18110_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_18111_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  or (_18112_, _18111_, _18110_);
  and (_18113_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_18114_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_18115_, _18114_, _18113_);
  or (_18116_, _18115_, _18112_);
  and (_18117_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_18118_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_18119_, _18118_, _18117_);
  and (_18120_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_18121_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_18122_, _18121_, _18120_);
  or (_18123_, _18122_, _18119_);
  or (_18124_, _18123_, _18116_);
  or (_18125_, _18124_, _18109_);
  and (_18126_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_18127_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_18128_, _18127_, _18126_);
  and (_18129_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_18130_, _17921_, _34767_);
  or (_18131_, _18130_, _18129_);
  or (_18132_, _18131_, _18128_);
  and (_18133_, _17925_, _17785_);
  and (_18134_, _17927_, _17664_);
  or (_18135_, _18134_, _18133_);
  and (_18136_, _17930_, _17574_);
  and (_18137_, _17932_, _17618_);
  or (_18138_, _18137_, _18136_);
  or (_18139_, _18138_, _18135_);
  or (_18140_, _18139_, _18132_);
  and (_18141_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_18142_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_18143_, _18142_, _18141_);
  or (_18144_, _18143_, _18140_);
  or (_18145_, _18144_, _18125_);
  and (_18146_, _18145_, _17848_);
  or (_18147_, _18146_, _17851_);
  or (_18148_, _18147_, _18094_);
  nand (_18149_, _17851_, _14356_);
  and (_18150_, _18149_, _38997_);
  and (_38989_[2], _18150_, _18148_);
  and (_18151_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_18152_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_18153_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_18154_, _18153_, _18152_);
  and (_18155_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_18156_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_18157_, _18156_, _18155_);
  or (_18158_, _18157_, _18154_);
  and (_18159_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_18160_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_18161_, _18160_, _18159_);
  and (_18162_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_18163_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_18164_, _18163_, _18162_);
  or (_18165_, _18164_, _18161_);
  or (_18166_, _18165_, _18158_);
  and (_18167_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_18168_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_18169_, _18168_, _18167_);
  and (_18170_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_18171_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_18172_, _18171_, _18170_);
  or (_18173_, _18172_, _18169_);
  and (_18174_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_18175_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_18176_, _18175_, _18174_);
  and (_18177_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_18178_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_18179_, _18178_, _18177_);
  or (_18180_, _18179_, _18176_);
  or (_18181_, _18180_, _18173_);
  or (_18182_, _18181_, _18166_);
  and (_18183_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_18184_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_18185_, _18184_, _18183_);
  and (_18186_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_18187_, _17921_, _34401_);
  or (_18188_, _18187_, _18186_);
  or (_18189_, _18188_, _18185_);
  and (_18190_, _17925_, _17754_);
  and (_18191_, _17927_, _17654_);
  or (_18192_, _18191_, _18190_);
  and (_18193_, _17930_, _17553_);
  and (_18194_, _17932_, _17597_);
  or (_18195_, _18194_, _18193_);
  or (_18196_, _18195_, _18192_);
  or (_18197_, _18196_, _18189_);
  and (_18198_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_18199_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_18200_, _18199_, _18198_);
  or (_18201_, _18200_, _18197_);
  or (_18202_, _18201_, _18182_);
  nand (_18203_, _18202_, _17848_);
  nand (_18204_, _18203_, _18037_);
  or (_18205_, _18204_, _18151_);
  nand (_18206_, _17851_, _14423_);
  and (_18207_, _18206_, _38997_);
  and (_38989_[3], _18207_, _18205_);
  and (_18208_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_18209_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_18210_, _18209_, _18208_);
  and (_18211_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_18212_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_18213_, _18212_, _18211_);
  or (_18214_, _18213_, _18210_);
  and (_18215_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_18216_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_18217_, _18216_, _18215_);
  and (_18218_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_18219_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_18220_, _18219_, _18218_);
  or (_18221_, _18220_, _18217_);
  or (_18222_, _18221_, _18214_);
  and (_18223_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_18224_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_18225_, _18224_, _18223_);
  and (_18226_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_18227_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or (_18228_, _18227_, _18226_);
  or (_18229_, _18228_, _18225_);
  and (_18230_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_18231_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_18232_, _18231_, _18230_);
  and (_18233_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_18234_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_18235_, _18234_, _18233_);
  or (_18236_, _18235_, _18232_);
  or (_18237_, _18236_, _18229_);
  or (_18238_, _18237_, _18222_);
  and (_18239_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_18240_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_18241_, _18240_, _18239_);
  and (_18242_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_18243_, _17921_, _34525_);
  or (_18244_, _18243_, _18242_);
  or (_18245_, _18244_, _18241_);
  and (_18246_, _17930_, _17539_);
  and (_18247_, _17932_, _17583_);
  or (_18248_, _18247_, _18246_);
  and (_18249_, _17927_, _17671_);
  and (_18250_, _17925_, _17771_);
  or (_18251_, _18250_, _18249_);
  or (_18252_, _18251_, _18248_);
  or (_18253_, _18252_, _18245_);
  and (_18254_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_18255_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_18256_, _18255_, _18254_);
  or (_18257_, _18256_, _18253_);
  or (_18258_, _18257_, _18238_);
  and (_18259_, _18258_, _17848_);
  and (_18260_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or (_18261_, _18260_, _18259_);
  or (_18262_, _18261_, _17851_);
  nand (_18263_, _17851_, _14495_);
  and (_18264_, _18263_, _38997_);
  and (_38989_[4], _18264_, _18262_);
  and (_18265_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_18266_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_18267_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_18268_, _18267_, _18266_);
  and (_18269_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_18270_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_18271_, _18270_, _18269_);
  or (_18272_, _18271_, _18268_);
  and (_18273_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_18274_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_18275_, _18274_, _18273_);
  and (_18276_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_18277_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_18278_, _18277_, _18276_);
  or (_18279_, _18278_, _18275_);
  or (_18280_, _18279_, _18272_);
  and (_18281_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_18282_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_18283_, _18282_, _18281_);
  and (_18284_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_18285_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_18286_, _18285_, _18284_);
  or (_18287_, _18286_, _18283_);
  and (_18288_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_18289_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_18290_, _18289_, _18288_);
  and (_18291_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_18292_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_18293_, _18292_, _18291_);
  or (_18294_, _18293_, _18290_);
  or (_18295_, _18294_, _18287_);
  or (_18296_, _18295_, _18280_);
  and (_18297_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_18298_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_18299_, _18298_, _18297_);
  and (_18300_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_18301_, _18013_, _34615_);
  or (_18302_, _18301_, _18300_);
  or (_18303_, _18302_, _18299_);
  and (_18304_, _17932_, _17604_);
  and (_18305_, _17930_, _17560_);
  or (_18306_, _18305_, _18304_);
  and (_18307_, _17927_, _17681_);
  and (_18308_, _17925_, _17760_);
  or (_18309_, _18308_, _18307_);
  or (_18310_, _18309_, _18306_);
  or (_18311_, _18310_, _18303_);
  and (_18312_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_18313_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_18314_, _18313_, _18312_);
  or (_18315_, _18314_, _18311_);
  or (_18316_, _18315_, _18296_);
  nand (_18317_, _18316_, _17848_);
  nand (_18318_, _18317_, _18037_);
  or (_18319_, _18318_, _18265_);
  nand (_18320_, _17851_, _14570_);
  and (_18321_, _18320_, _38997_);
  and (_38989_[5], _18321_, _18319_);
  and (_18322_, _17967_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_18323_, _17855_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nand (_18324_, _17858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_18325_, _18324_, _18323_);
  nand (_18326_, _17863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand (_18327_, _17866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_18328_, _18327_, _18326_);
  and (_18329_, _18328_, _18325_);
  nand (_18330_, _17870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_18331_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_18332_, _18331_, _18330_);
  nand (_18333_, _17878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand (_18334_, _17881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_18335_, _18334_, _18333_);
  and (_18336_, _18335_, _18332_);
  and (_18337_, _18336_, _18329_);
  nand (_18338_, _17886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_18339_, _17889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_18340_, _18339_, _18338_);
  nand (_18341_, _17892_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_18342_, _17894_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_18343_, _18342_, _18341_);
  and (_18344_, _18343_, _18340_);
  nand (_18345_, _17899_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand (_18346_, _17901_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_18347_, _18346_, _18345_);
  nand (_18348_, _17906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand (_18349_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_18350_, _18349_, _18348_);
  and (_18351_, _18350_, _18347_);
  and (_18352_, _18351_, _18344_);
  and (_18353_, _18352_, _18337_);
  nand (_18354_, _17850_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand (_18355_, _17914_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_18356_, _18355_, _18354_);
  nand (_18357_, _17918_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_18358_, _18013_, _34649_);
  and (_18359_, _18358_, _18357_);
  and (_18360_, _18359_, _18356_);
  nand (_18361_, _17927_, _17660_);
  nand (_18362_, _17925_, _17781_);
  and (_18363_, _18362_, _18361_);
  nand (_18364_, _17932_, _17614_);
  nand (_18365_, _17930_, _17570_);
  and (_18366_, _18365_, _18364_);
  and (_18367_, _18366_, _18363_);
  and (_18368_, _18367_, _18360_);
  nand (_18369_, _17844_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_18370_, _17834_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_18371_, _18370_, _18369_);
  and (_18372_, _18371_, _18368_);
  nand (_18373_, _18372_, _18353_);
  nand (_18374_, _18373_, _17848_);
  nand (_18375_, _18374_, _18037_);
  or (_18376_, _18375_, _18322_);
  or (_18377_, _18037_, _14632_);
  and (_18378_, _18377_, _38997_);
  and (_38989_[6], _18378_, _18376_);
  and (_36924_, _34788_, _38997_);
  and (_36925_[7], _35813_, _38997_);
  nor (_36927_[2], _34770_, rst);
  and (_36925_[0], _35732_, _38997_);
  and (_36925_[1], _35748_, _38997_);
  and (_36925_[2], _35757_, _38997_);
  and (_36925_[3], _35767_, _38997_);
  and (_36925_[4], _35778_, _38997_);
  and (_36925_[5], _35791_, _38997_);
  and (_36925_[6], _35802_, _38997_);
  nor (_36927_[0], _34471_, rst);
  nor (_36927_[1], _34579_, rst);
  nor (_18379_, _16449_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_18380_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18381_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _18380_);
  nor (_18382_, _18381_, _18379_);
  nor (_18383_, _16471_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18384_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _18380_);
  nor (_18385_, _18384_, _18383_);
  nor (_18386_, _18385_, _18382_);
  and (_18387_, _18386_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_18388_, _18385_, _18382_);
  and (_18389_, _18388_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_18390_, _18389_, _18387_);
  not (_18391_, _18382_);
  and (_18392_, _18385_, _18391_);
  and (_18393_, _18392_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18394_, _18385_, _18391_);
  and (_18395_, _18394_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_18396_, _18395_, _18393_);
  and (_18397_, _18396_, _18390_);
  nor (_18398_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18399_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _18380_);
  nor (_18400_, _18399_, _18398_);
  nor (_18401_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_18402_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _18380_);
  nor (_18403_, _18402_, _18401_);
  and (_18404_, _18403_, _18400_);
  not (_18405_, _18404_);
  nor (_18406_, _18405_, _18397_);
  and (_18407_, _18394_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_18408_, _18386_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_18409_, _18408_, _18407_);
  and (_18410_, _18392_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_18411_, _18388_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_18412_, _18411_, _18410_);
  and (_18413_, _18412_, _18409_);
  nor (_18414_, _18403_, _18400_);
  not (_18415_, _18414_);
  nor (_18416_, _18415_, _18413_);
  nor (_18417_, _18416_, _18406_);
  and (_18418_, _18392_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_18419_, _18386_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_18420_, _18419_, _18418_);
  and (_18421_, _18394_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_18422_, _18388_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_18423_, _18422_, _18421_);
  and (_18424_, _18423_, _18420_);
  not (_18425_, _18403_);
  and (_18426_, _18425_, _18400_);
  not (_18427_, _18426_);
  nor (_18428_, _18427_, _18424_);
  and (_18429_, _18388_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_18430_, _18386_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_18431_, _18430_, _18429_);
  and (_18432_, _18392_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_18433_, _18394_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_18434_, _18433_, _18432_);
  and (_18435_, _18434_, _18431_);
  not (_18436_, _18400_);
  and (_18437_, _18403_, _18436_);
  not (_18438_, _18437_);
  nor (_18439_, _18438_, _18435_);
  nor (_18440_, _18439_, _18428_);
  and (_18441_, _18440_, _18417_);
  and (_18442_, _18441_, word_in[7]);
  not (_18443_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_18444_, _18400_, _18443_);
  or (_18445_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_18446_, _18445_, _18444_);
  nor (_18447_, _18403_, _18382_);
  and (_18448_, _18447_, _18446_);
  or (_18449_, _18448_, _18385_);
  and (_18450_, _18403_, _18382_);
  not (_18451_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_18452_, _18400_, _18451_);
  or (_18453_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_18454_, _18453_, _18452_);
  and (_18455_, _18454_, _18450_);
  and (_18456_, _18425_, _18382_);
  not (_18457_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_18458_, _18400_, _18457_);
  or (_18459_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_18460_, _18459_, _18458_);
  and (_18461_, _18460_, _18456_);
  not (_18462_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_18463_, _18400_, _18462_);
  or (_18464_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_18465_, _18464_, _18463_);
  nor (_18466_, _18425_, _18382_);
  and (_18467_, _18466_, _18465_);
  or (_18468_, _18467_, _18461_);
  or (_18469_, _18468_, _18455_);
  or (_18470_, _18469_, _18449_);
  not (_18471_, _18385_);
  not (_18472_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_18473_, _18400_, _18472_);
  or (_18474_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_18475_, _18474_, _18473_);
  and (_18476_, _18475_, _18447_);
  or (_18477_, _18476_, _18471_);
  not (_18478_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_18479_, _18400_, _18478_);
  or (_18480_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_18481_, _18480_, _18479_);
  and (_18482_, _18481_, _18456_);
  not (_18483_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_18484_, _18400_, _18483_);
  or (_18485_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_18486_, _18485_, _18484_);
  and (_18487_, _18486_, _18450_);
  or (_18488_, _18487_, _18482_);
  not (_18489_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_18490_, _18400_, _18489_);
  or (_18491_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_18492_, _18491_, _18490_);
  and (_18493_, _18492_, _18466_);
  or (_18494_, _18493_, _18488_);
  or (_18495_, _18494_, _18477_);
  nand (_18496_, _18495_, _18470_);
  nor (_18497_, _18496_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _18497_, _18442_);
  nor (_18498_, _18404_, _18382_);
  and (_18499_, _18404_, _18382_);
  nor (_18500_, _18499_, _18498_);
  not (_18501_, _18500_);
  nor (_18502_, _18499_, _18471_);
  and (_18503_, _18404_, _18394_);
  nor (_18504_, _18503_, _18502_);
  and (_18505_, _18504_, _18501_);
  and (_18506_, _18505_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_18507_, _18506_);
  not (_18508_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand (_18509_, _18504_, _18508_);
  nor (_18510_, _18504_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_18511_, _18510_, _18501_);
  and (_18512_, _18511_, _18509_);
  nor (_18513_, _18504_, _18500_);
  and (_18514_, _18513_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18515_, _18514_, _18512_);
  and (_18516_, _18515_, _18507_);
  nor (_18517_, _18516_, _18415_);
  and (_18518_, _18505_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_18519_, _18518_);
  not (_18520_, _18504_);
  or (_18521_, _18520_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_18522_, _18504_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_18523_, _18522_, _18501_);
  and (_18524_, _18523_, _18521_);
  and (_18525_, _18513_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18526_, _18525_, _18524_);
  and (_18527_, _18526_, _18519_);
  nor (_18528_, _18527_, _18438_);
  nor (_18529_, _18528_, _18517_);
  and (_18530_, _18505_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_18531_, _18530_);
  not (_18532_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand (_18533_, _18504_, _18532_);
  nor (_18534_, _18504_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_18535_, _18534_, _18501_);
  and (_18536_, _18535_, _18533_);
  and (_18537_, _18513_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_18538_, _18537_, _18536_);
  and (_18539_, _18538_, _18531_);
  nor (_18540_, _18539_, _18405_);
  and (_18541_, _18505_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_18542_, _18541_);
  not (_18543_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand (_18544_, _18504_, _18543_);
  nor (_18545_, _18504_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_18546_, _18545_, _18501_);
  and (_18547_, _18546_, _18544_);
  and (_18548_, _18513_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18549_, _18548_, _18547_);
  and (_18550_, _18549_, _18542_);
  nor (_18551_, _18550_, _18427_);
  nor (_18552_, _18551_, _18540_);
  and (_18553_, _18552_, _18529_);
  and (_18554_, _18553_, word_in[15]);
  or (_18555_, _18414_, _18404_);
  not (_18556_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_18557_, _18400_, _18556_);
  or (_18558_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_18559_, _18558_, _18557_);
  and (_18560_, _18559_, _18555_);
  not (_18561_, _18555_);
  and (_18562_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor (_18563_, _18400_, _18462_);
  or (_18564_, _18563_, _18562_);
  and (_18565_, _18564_, _18561_);
  nor (_18566_, _18565_, _18560_);
  nor (_18567_, _18566_, _18500_);
  and (_18568_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_18569_, _18400_, _18457_);
  or (_18570_, _18569_, _18568_);
  and (_18571_, _18570_, _18555_);
  not (_18572_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_18573_, _18400_, _18572_);
  or (_18574_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_18575_, _18574_, _18573_);
  and (_18576_, _18575_, _18561_);
  or (_18577_, _18576_, _18571_);
  and (_18578_, _18577_, _18500_);
  nor (_18579_, _18578_, _18567_);
  nand (_18580_, _18579_, _18504_);
  not (_18581_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_18582_, _18400_, _18581_);
  or (_18583_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_18584_, _18583_, _18582_);
  and (_18585_, _18584_, _18555_);
  not (_18586_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_18587_, _18400_, _18586_);
  or (_18588_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_18589_, _18588_, _18587_);
  and (_18590_, _18589_, _18561_);
  nor (_18591_, _18590_, _18585_);
  nor (_18592_, _18591_, _18500_);
  not (_18593_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_18594_, _18400_, _18593_);
  or (_18595_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_18596_, _18595_, _18594_);
  and (_18597_, _18596_, _18555_);
  not (_18598_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_18599_, _18400_, _18598_);
  or (_18600_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_18601_, _18600_, _18599_);
  and (_18602_, _18601_, _18561_);
  or (_18603_, _18602_, _18597_);
  and (_18604_, _18603_, _18500_);
  or (_18605_, _18604_, _18592_);
  or (_18606_, _18605_, _18504_);
  nand (_18607_, _18606_, _18580_);
  nor (_18608_, _18607_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _18608_, _18554_);
  not (_18609_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_18610_, _18450_, _18471_);
  not (_18611_, _18610_);
  or (_18612_, _18450_, _18471_);
  and (_18613_, _18612_, _18611_);
  and (_18614_, _18613_, _18609_);
  nor (_18615_, _18450_, _18447_);
  not (_18616_, _18615_);
  and (_18617_, _18616_, _18613_);
  and (_18618_, _18616_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18619_, _18618_, _18617_);
  nor (_18620_, _18619_, _18614_);
  and (_18621_, _18613_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_18622_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_18623_, _18613_, _18622_);
  nor (_18624_, _18623_, _18621_);
  nor (_18625_, _18624_, _18391_);
  nor (_18626_, _18625_, _18620_);
  nor (_18627_, _18626_, _18403_);
  and (_18628_, _18613_, _18508_);
  not (_18629_, _18466_);
  not (_18630_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_18631_, _18385_, _18630_);
  nor (_18632_, _18631_, _18629_);
  not (_18633_, _18632_);
  nor (_18634_, _18633_, _18628_);
  not (_18635_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_18636_, _18613_, _18635_);
  and (_18637_, _18450_, _18385_);
  and (_18638_, _18450_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18639_, _18638_, _18637_);
  nor (_18640_, _18639_, _18636_);
  or (_18641_, _18640_, _18436_);
  or (_18642_, _18641_, _18634_);
  nor (_18643_, _18642_, _18627_);
  not (_18644_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_18645_, _18613_, _18644_);
  not (_18646_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18647_, _18615_, _18646_);
  nor (_18648_, _18647_, _18617_);
  nor (_18649_, _18648_, _18645_);
  and (_18650_, _18613_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_18651_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_18652_, _18613_, _18651_);
  nor (_18653_, _18652_, _18650_);
  nor (_18654_, _18653_, _18391_);
  nor (_18655_, _18654_, _18649_);
  nor (_18656_, _18655_, _18403_);
  not (_18657_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_18658_, _18613_, _18657_);
  and (_18659_, _18450_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_18660_, _18659_, _18637_);
  nor (_18661_, _18660_, _18658_);
  and (_18662_, _18613_, _18532_);
  not (_18663_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18664_, _18385_, _18663_);
  nor (_18665_, _18664_, _18629_);
  not (_18666_, _18665_);
  nor (_18667_, _18666_, _18662_);
  or (_18668_, _18667_, _18400_);
  or (_18669_, _18668_, _18661_);
  nor (_18670_, _18669_, _18656_);
  nor (_18671_, _18670_, _18643_);
  not (_18672_, _18671_);
  and (_18673_, _18672_, word_in[23]);
  and (_18674_, _18466_, _18460_);
  and (_18675_, _18465_, _18447_);
  or (_18676_, _18675_, _18674_);
  and (_18677_, _18456_, _18454_);
  and (_18678_, _18450_, _18446_);
  or (_18679_, _18678_, _18677_);
  nor (_18680_, _18679_, _18676_);
  nand (_18681_, _18680_, _18613_);
  and (_18682_, _18481_, _18466_);
  and (_18683_, _18492_, _18447_);
  or (_18684_, _18683_, _18682_);
  and (_18685_, _18486_, _18456_);
  and (_18686_, _18475_, _18450_);
  or (_18687_, _18686_, _18685_);
  or (_18688_, _18687_, _18684_);
  or (_18689_, _18688_, _18613_);
  and (_18690_, _18689_, _18681_);
  and (_18691_, _18690_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _18691_, _18673_);
  and (_18692_, _18415_, _18382_);
  and (_18693_, _18692_, _18385_);
  nor (_18694_, _18692_, _18385_);
  nor (_18695_, _18694_, _18693_);
  nor (_18696_, _18695_, \oc8051_symbolic_cxrom1.regvalid [5]);
  not (_18697_, _18696_);
  nor (_18698_, _18415_, _18382_);
  nor (_18699_, _18692_, _18698_);
  not (_18700_, _18699_);
  nor (_18701_, _18700_, _18631_);
  and (_18702_, _18701_, _18697_);
  nor (_18703_, _18695_, _18635_);
  and (_18704_, _18695_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18705_, _18704_, _18703_);
  nor (_18706_, _18705_, _18699_);
  nor (_18707_, _18706_, _18702_);
  nor (_18708_, _18707_, _18438_);
  nor (_18709_, _18695_, _18657_);
  and (_18710_, _18695_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_18711_, _18710_, _18709_);
  nor (_18712_, _18711_, _18699_);
  nor (_18713_, _18695_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_18714_, _18713_);
  nor (_18715_, _18700_, _18664_);
  and (_18716_, _18715_, _18714_);
  nor (_18717_, _18716_, _18712_);
  nor (_18718_, _18717_, _18427_);
  nor (_18719_, _18718_, _18708_);
  nor (_18720_, _18695_, _18609_);
  and (_18721_, _18695_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_18722_, _18721_, _18720_);
  nor (_18723_, _18722_, _18699_);
  nand (_18724_, _18695_, _18622_);
  nor (_18725_, _18695_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_18726_, _18725_, _18700_);
  and (_18727_, _18726_, _18724_);
  nor (_18728_, _18727_, _18723_);
  nor (_18729_, _18728_, _18415_);
  nor (_18730_, _18695_, _18644_);
  and (_18731_, _18695_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18732_, _18731_, _18730_);
  nor (_18733_, _18732_, _18699_);
  nand (_18734_, _18695_, _18651_);
  nor (_18735_, _18695_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_18736_, _18735_, _18700_);
  and (_18737_, _18736_, _18734_);
  nor (_18738_, _18737_, _18733_);
  nor (_18739_, _18738_, _18405_);
  nor (_18740_, _18739_, _18729_);
  and (_18741_, _18740_, _18719_);
  and (_18742_, _18601_, _18555_);
  and (_18743_, _18596_, _18561_);
  or (_18744_, _18743_, _18742_);
  and (_18745_, _18744_, _18699_);
  and (_18746_, _18589_, _18555_);
  and (_18747_, _18584_, _18561_);
  nor (_18748_, _18747_, _18746_);
  nor (_18749_, _18748_, _18699_);
  or (_18750_, _18749_, _18745_);
  and (_18751_, _18750_, _18695_);
  not (_18752_, _18695_);
  and (_18753_, _18575_, _18555_);
  and (_18754_, _18570_, _18561_);
  or (_18755_, _18754_, _18753_);
  and (_18756_, _18755_, _18699_);
  and (_18757_, _18564_, _18555_);
  and (_18758_, _18559_, _18561_);
  nor (_18759_, _18758_, _18757_);
  nor (_18760_, _18759_, _18699_);
  or (_18761_, _18760_, _18756_);
  and (_18762_, _18761_, _18752_);
  nor (_18763_, _18762_, _18751_);
  nor (_18764_, _18763_, _18741_);
  and (_18765_, _18741_, word_in[31]);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _18765_, _18764_);
  or (_18766_, _18388_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_36729_[15], _18766_, _38997_);
  and (_18767_, _18741_, _38997_);
  and (_18768_, _18767_, word_in[31]);
  and (_18769_, _18414_, _18388_);
  and (_18770_, _18767_, _18769_);
  and (_18771_, _18770_, _18768_);
  not (_18772_, _18770_);
  and (_18773_, _18643_, _38997_);
  and (_18774_, _18773_, _18425_);
  not (_18775_, _18613_);
  nor (_18776_, _18671_, rst);
  and (_18777_, _18776_, _18775_);
  and (_18778_, _18777_, _18615_);
  and (_18779_, _18778_, _18774_);
  and (_18780_, _18553_, _38997_);
  and (_18781_, _18780_, _18500_);
  and (_18782_, _18781_, _18520_);
  and (_18783_, _18782_, _18437_);
  and (_18784_, _18499_, _18385_);
  and (_18785_, _18441_, _38997_);
  and (_18786_, _18785_, _18784_);
  and (_18787_, _18786_, word_in[7]);
  nor (_18788_, _18786_, _18483_);
  nor (_18789_, _18788_, _18787_);
  nor (_18790_, _18789_, _18783_);
  and (_18791_, _18780_, word_in[15]);
  and (_18792_, _18791_, _18783_);
  nor (_18793_, _18792_, _18790_);
  nor (_18794_, _18793_, _18779_);
  and (_18795_, _18776_, word_in[23]);
  and (_18796_, _18795_, _18779_);
  or (_18797_, _18796_, _18794_);
  and (_18798_, _18797_, _18772_);
  or (_36785_, _18798_, _18771_);
  and (_18799_, _18414_, _18386_);
  or (_18800_, _18693_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_18801_, _18800_, _18799_);
  and (_36858_, _18801_, _38997_);
  and (_18802_, _18425_, _18386_);
  or (_18803_, _18784_, _18802_);
  and (_18804_, _18437_, _18388_);
  or (_18805_, _18804_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_18806_, _18805_, _18803_);
  and (_36729_[1], _18806_, _38997_);
  and (_18807_, _18437_, _18386_);
  or (_18808_, _18807_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_18809_, _18808_, _18803_);
  and (_36729_[2], _18809_, _38997_);
  or (_18810_, _18386_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_36729_[3], _18810_, _38997_);
  and (_18811_, _18414_, _18394_);
  nand (_18812_, _18694_, _18405_);
  and (_18813_, _18812_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_18814_, _18813_, _18811_);
  nor (_18815_, _18814_, _18386_);
  and (_18816_, _18404_, _18386_);
  and (_18817_, _18426_, _18386_);
  and (_18818_, _18799_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_18819_, _18818_, _18817_);
  or (_18820_, _18819_, _18816_);
  or (_18821_, _18820_, _18807_);
  or (_18822_, _18821_, _18815_);
  and (_36729_[4], _18822_, _38997_);
  nor (_18823_, _18784_, _18386_);
  and (_18824_, _18426_, _18394_);
  or (_18825_, _18824_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_18826_, _18694_, _18784_);
  and (_18827_, _18826_, _18825_);
  nor (_18828_, _18385_, _18508_);
  and (_18829_, _18466_, _18828_);
  or (_18830_, _18829_, _18811_);
  or (_18831_, _18830_, _18827_);
  and (_18832_, _18831_, _18823_);
  and (_18833_, _18817_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_18834_, _18833_, _18807_);
  and (_18835_, _18698_, _18828_);
  and (_18836_, _18825_, _18784_);
  or (_18837_, _18836_, _18835_);
  or (_18838_, _18837_, _18834_);
  or (_18839_, _18838_, _18816_);
  or (_18840_, _18839_, _18832_);
  and (_36729_[5], _18840_, _38997_);
  not (_18841_, _18824_);
  nor (_18842_, _18816_, _18811_);
  nand (_18843_, _18842_, _18841_);
  and (_18844_, _18405_, _18386_);
  and (_18845_, _18844_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_18846_, _18450_, _18385_);
  and (_18847_, _18437_, _18394_);
  or (_18848_, _18400_, _18385_);
  nor (_18849_, _18386_, _18543_);
  and (_18850_, _18849_, _18848_);
  or (_18851_, _18850_, _18847_);
  and (_18852_, _18851_, _18846_);
  or (_18853_, _18852_, _18845_);
  or (_18854_, _18853_, _18843_);
  and (_36729_[6], _18854_, _38997_);
  or (_18855_, _18502_, _18610_);
  and (_18856_, _18425_, _18395_);
  nand (_18857_, _18438_, _18394_);
  and (_18858_, _18857_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_18859_, _18858_, _18856_);
  and (_18860_, _18859_, _18502_);
  or (_18861_, _18856_, _18610_);
  or (_18862_, _18861_, _18860_);
  and (_18863_, _18862_, _18855_);
  and (_18864_, _18859_, _18784_);
  and (_18865_, _18807_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_18866_, _18816_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_18867_, _18802_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_18868_, _18867_, _18811_);
  or (_18869_, _18868_, _18866_);
  or (_18870_, _18869_, _18865_);
  or (_18871_, _18870_, _18864_);
  or (_18872_, _18871_, _18824_);
  or (_18873_, _18872_, _18863_);
  and (_36729_[7], _18873_, _38997_);
  and (_18874_, _18561_, _18386_);
  not (_18875_, _18698_);
  nand (_18876_, _18842_, _18875_);
  or (_18877_, _18876_, _18874_);
  and (_18878_, _18877_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_18879_, _18400_, _18394_);
  or (_18880_, _18698_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_18881_, _18880_, _18385_);
  or (_18882_, _18881_, _18879_);
  or (_18883_, _18882_, _18847_);
  or (_18884_, _18883_, _18878_);
  and (_36729_[8], _18884_, _38997_);
  not (_18885_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_18886_, _18846_, _18885_);
  and (_18887_, _18846_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_18888_, _18426_, _18392_);
  or (_18889_, _18888_, _18698_);
  or (_18890_, _18889_, _18887_);
  and (_18891_, _18890_, _18385_);
  or (_18892_, _18891_, _18610_);
  or (_18893_, _18892_, _18886_);
  and (_36729_[9], _18893_, _38997_);
  and (_18894_, _18615_, _18385_);
  or (_18895_, _18894_, _18804_);
  or (_18896_, _18895_, _18784_);
  nand (_18897_, _18561_, _18394_);
  nand (_18898_, _18842_, _18897_);
  and (_18899_, _18898_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_18900_, _18437_, _18392_);
  and (_18901_, _18799_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_18902_, _18874_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_18903_, _18902_, _18901_);
  or (_18904_, _18903_, _18900_);
  and (_18905_, _18698_, _18385_);
  or (_18906_, _18905_, _18503_);
  and (_18907_, _18906_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_18908_, _18498_, _18471_);
  or (_18909_, _18908_, _18888_);
  and (_18910_, _18909_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_18911_, _18910_, _18907_);
  or (_18912_, _18911_, _18904_);
  or (_18913_, _18912_, _18899_);
  and (_18914_, _18913_, _18896_);
  nor (_18915_, _18824_, _18807_);
  and (_18916_, _18915_, _18842_);
  nor (_18917_, _18916_, _18646_);
  and (_18918_, _18847_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_18919_, _18802_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_18920_, _18919_, _18503_);
  or (_18921_, _18920_, _18918_);
  or (_18922_, _18921_, _18917_);
  or (_18923_, _18922_, _18888_);
  or (_18924_, _18923_, _18905_);
  or (_18925_, _18924_, _18914_);
  and (_36729_[10], _18925_, _38997_);
  and (_18926_, _18404_, _18392_);
  or (_18927_, _18926_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_18928_, _18500_, _18385_);
  and (_18929_, _18928_, _18927_);
  or (_18930_, _18811_, _18824_);
  and (_18931_, _18930_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_18932_, _18847_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_18933_, _18932_, _18931_);
  and (_18934_, _18816_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_18935_, _18934_, _18933_);
  and (_18936_, _18905_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_18937_, _18874_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_18938_, _18937_, _18936_);
  and (_18939_, _18888_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_18940_, _18503_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_18941_, _18940_, _18900_);
  or (_18942_, _18941_, _18939_);
  or (_18943_, _18942_, _18938_);
  or (_18944_, _18943_, _18935_);
  or (_18945_, _18944_, _18929_);
  and (_18946_, _18945_, _18895_);
  or (_18947_, _18937_, _18940_);
  or (_18948_, _18947_, _18935_);
  and (_18949_, _18799_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_18950_, _18784_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_18951_, _18950_, _18949_);
  or (_18952_, _18951_, _18905_);
  or (_18953_, _18952_, _18948_);
  or (_18954_, _18953_, _18888_);
  or (_18955_, _18954_, _18946_);
  and (_36729_[11], _18955_, _38997_);
  and (_18956_, _18693_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18957_, _18415_, _18394_);
  and (_18958_, _18957_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18959_, _18816_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18960_, _18811_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18961_, _18698_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_18962_, _18961_, _18888_);
  or (_18963_, _18962_, _18960_);
  or (_18964_, _18963_, _18959_);
  and (_18965_, _18874_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_18966_, _18426_, _18388_);
  not (_18967_, _18966_);
  and (_18968_, _18894_, _18967_);
  or (_18969_, _18968_, _18965_);
  or (_18970_, _18969_, _18964_);
  or (_18971_, _18970_, _18958_);
  or (_18972_, _18971_, _18956_);
  and (_36729_[12], _18972_, _38997_);
  or (_18973_, _18894_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_36729_[13], _18973_, _38997_);
  or (_18974_, _18928_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_36729_[14], _18974_, _38997_);
  and (_18975_, _18767_, _18699_);
  and (_18976_, _18767_, _18695_);
  nor (_18977_, _18976_, _18975_);
  and (_18978_, _18977_, _18426_);
  and (_18979_, _18978_, _18767_);
  and (_18980_, _18776_, _18425_);
  nor (_18981_, _18980_, _18773_);
  and (_18982_, _18981_, _18776_);
  and (_18983_, _18982_, _18617_);
  and (_18984_, _18780_, _18784_);
  not (_18985_, _18984_);
  or (_18986_, _18985_, word_in[8]);
  not (_18987_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_18988_, _18785_, _18799_);
  nor (_18989_, _18988_, _18987_);
  and (_18990_, _18988_, word_in[0]);
  or (_18991_, _18990_, _18989_);
  or (_18992_, _18991_, _18984_);
  and (_18993_, _18992_, _18986_);
  or (_18994_, _18993_, _18983_);
  not (_18995_, _18983_);
  or (_18996_, _18995_, word_in[16]);
  and (_18997_, _18996_, _18994_);
  or (_18998_, _18997_, _18979_);
  not (_18999_, _18979_);
  or (_19000_, _18999_, word_in[24]);
  and (_36730_, _19000_, _18998_);
  and (_19001_, _18780_, word_in[9]);
  and (_19002_, _19001_, _18984_);
  not (_19003_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_19004_, _18988_, _19003_);
  and (_19005_, _18988_, word_in[1]);
  nor (_19006_, _19005_, _19004_);
  nor (_19007_, _19006_, _18984_);
  or (_19008_, _19007_, _19002_);
  or (_19009_, _19008_, _18983_);
  or (_19010_, _18995_, word_in[17]);
  and (_19011_, _19010_, _19009_);
  or (_19012_, _19011_, _18979_);
  or (_19013_, _18999_, word_in[25]);
  and (_36731_, _19013_, _19012_);
  or (_19014_, _18985_, word_in[10]);
  and (_19015_, _18988_, word_in[2]);
  not (_19016_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_19017_, _18988_, _19016_);
  or (_19018_, _19017_, _19015_);
  or (_19019_, _19018_, _18984_);
  and (_19020_, _19019_, _19014_);
  or (_19021_, _19020_, _18983_);
  or (_19022_, _18995_, word_in[18]);
  and (_19023_, _19022_, _19021_);
  or (_19024_, _19023_, _18979_);
  or (_19025_, _18999_, word_in[26]);
  and (_36732_, _19025_, _19024_);
  or (_19026_, _18985_, word_in[11]);
  not (_19027_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_19028_, _18988_, _19027_);
  and (_19029_, _18988_, word_in[3]);
  or (_19030_, _19029_, _19028_);
  or (_19031_, _19030_, _18984_);
  and (_19032_, _19031_, _19026_);
  or (_19033_, _19032_, _18983_);
  or (_19034_, _18995_, word_in[19]);
  and (_19035_, _19034_, _19033_);
  or (_19036_, _19035_, _18979_);
  or (_19037_, _18999_, word_in[27]);
  and (_36733_, _19037_, _19036_);
  and (_19038_, _18767_, word_in[28]);
  and (_19039_, _19038_, _18978_);
  or (_19040_, _18995_, word_in[20]);
  or (_19041_, _18985_, word_in[12]);
  not (_19042_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_19043_, _18988_, _19042_);
  and (_19044_, _18988_, word_in[4]);
  or (_19045_, _19044_, _19043_);
  or (_19046_, _19045_, _18984_);
  and (_19047_, _19046_, _19041_);
  or (_19048_, _19047_, _18983_);
  and (_19049_, _19048_, _18999_);
  and (_19050_, _19049_, _19040_);
  or (_36734_, _19050_, _19039_);
  or (_19051_, _18995_, word_in[21]);
  or (_19052_, _18985_, word_in[13]);
  and (_19053_, _18988_, word_in[5]);
  not (_19054_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_19055_, _18988_, _19054_);
  or (_19056_, _19055_, _19053_);
  or (_19057_, _19056_, _18984_);
  and (_19058_, _19057_, _19052_);
  or (_19059_, _19058_, _18983_);
  and (_19060_, _19059_, _18999_);
  and (_19061_, _19060_, _19051_);
  and (_19062_, _18979_, word_in[29]);
  or (_36735_, _19062_, _19061_);
  or (_19063_, _18985_, word_in[14]);
  and (_19064_, _18988_, word_in[6]);
  not (_19065_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_19066_, _18988_, _19065_);
  or (_19067_, _19066_, _19064_);
  or (_19068_, _19067_, _18984_);
  and (_19069_, _19068_, _19063_);
  or (_19070_, _19069_, _18983_);
  or (_19071_, _18995_, word_in[22]);
  and (_19072_, _19071_, _19070_);
  or (_19073_, _19072_, _18979_);
  or (_19074_, _18999_, word_in[30]);
  and (_36736_, _19074_, _19073_);
  or (_19075_, _18985_, word_in[15]);
  and (_19076_, _18988_, word_in[7]);
  nor (_19077_, _18988_, _18556_);
  or (_19078_, _19077_, _19076_);
  or (_19079_, _19078_, _18984_);
  and (_19080_, _19079_, _19075_);
  or (_19081_, _19080_, _18983_);
  or (_19082_, _18995_, word_in[23]);
  and (_19083_, _19082_, _19081_);
  or (_19084_, _19083_, _18979_);
  or (_19085_, _18999_, word_in[31]);
  and (_36737_, _19085_, _19084_);
  and (_19086_, _18767_, _18437_);
  and (_19087_, _19086_, _18977_);
  not (_19088_, _18617_);
  and (_19089_, _18776_, _19088_);
  and (_19090_, _18773_, _18403_);
  not (_19091_, _19090_);
  nor (_19092_, _19091_, _19089_);
  and (_19093_, _18780_, _18799_);
  nand (_19094_, _18785_, _18817_);
  and (_19095_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_19096_, _18785_, word_in[0]);
  and (_19097_, _19096_, _18817_);
  or (_19098_, _19097_, _19095_);
  or (_19099_, _19098_, _19093_);
  not (_19100_, _19093_);
  or (_19101_, _19100_, word_in[8]);
  and (_19102_, _19101_, _19099_);
  or (_19103_, _19102_, _19092_);
  and (_19104_, _18776_, word_in[16]);
  not (_19105_, _19092_);
  or (_19106_, _19105_, _19104_);
  and (_19107_, _19106_, _19103_);
  or (_19108_, _19107_, _19087_);
  not (_19109_, _19087_);
  or (_19110_, _19109_, word_in[24]);
  and (_36786_, _19110_, _19108_);
  and (_19111_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_19112_, _18785_, word_in[1]);
  and (_19113_, _19112_, _18817_);
  nor (_19114_, _19113_, _19111_);
  nor (_19115_, _19114_, _19093_);
  and (_19116_, _19093_, word_in[9]);
  nor (_19117_, _19116_, _19115_);
  nor (_19118_, _19117_, _19092_);
  and (_19119_, _18776_, word_in[17]);
  and (_19120_, _19092_, _19119_);
  or (_19121_, _19120_, _19087_);
  or (_19122_, _19121_, _19118_);
  or (_19123_, _19109_, word_in[25]);
  and (_36787_, _19123_, _19122_);
  and (_19124_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_19125_, _18785_, word_in[2]);
  and (_19126_, _19125_, _18817_);
  nor (_19127_, _19126_, _19124_);
  nor (_19128_, _19127_, _19093_);
  and (_19129_, _19093_, word_in[10]);
  nor (_19130_, _19129_, _19128_);
  nor (_19131_, _19130_, _19092_);
  and (_19132_, _18776_, word_in[18]);
  and (_19133_, _19092_, _19132_);
  or (_19134_, _19133_, _19087_);
  or (_19135_, _19134_, _19131_);
  or (_19136_, _19109_, word_in[26]);
  and (_36788_, _19136_, _19135_);
  and (_19137_, _18785_, word_in[3]);
  and (_19138_, _19137_, _18817_);
  and (_19139_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_19140_, _19139_, _19138_);
  nor (_19141_, _19140_, _19093_);
  and (_19142_, _19093_, word_in[11]);
  nor (_19143_, _19142_, _19141_);
  nor (_19144_, _19143_, _19092_);
  and (_19145_, _18776_, word_in[19]);
  and (_19146_, _19092_, _19145_);
  or (_19147_, _19146_, _19087_);
  or (_19148_, _19147_, _19144_);
  or (_19149_, _19109_, word_in[27]);
  and (_36789_, _19149_, _19148_);
  and (_19150_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_19151_, _18785_, word_in[4]);
  and (_19152_, _19151_, _18817_);
  or (_19153_, _19152_, _19150_);
  or (_19154_, _19153_, _19093_);
  or (_19155_, _19100_, word_in[12]);
  and (_19156_, _19155_, _19154_);
  or (_19157_, _19156_, _19092_);
  and (_19158_, _18776_, word_in[20]);
  or (_19159_, _19105_, _19158_);
  and (_19160_, _19159_, _19157_);
  or (_19161_, _19160_, _19087_);
  or (_19162_, _19109_, word_in[28]);
  and (_36790_, _19162_, _19161_);
  and (_19163_, _18785_, word_in[5]);
  and (_19164_, _19163_, _18817_);
  and (_19165_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_19166_, _19165_, _19164_);
  nor (_19167_, _19166_, _19093_);
  and (_19168_, _19093_, word_in[13]);
  nor (_19169_, _19168_, _19167_);
  nor (_19170_, _19169_, _19092_);
  and (_19171_, _18776_, word_in[21]);
  and (_19172_, _19092_, _19171_);
  or (_19173_, _19172_, _19087_);
  or (_19174_, _19173_, _19170_);
  or (_19175_, _19109_, word_in[29]);
  and (_36791_, _19175_, _19174_);
  and (_19176_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_19177_, _18785_, word_in[6]);
  and (_19178_, _19177_, _18817_);
  nor (_19179_, _19178_, _19176_);
  nor (_19180_, _19179_, _19093_);
  and (_19181_, _19093_, word_in[14]);
  nor (_19182_, _19181_, _19180_);
  nor (_19183_, _19182_, _19092_);
  and (_19184_, _18776_, word_in[22]);
  and (_19185_, _19092_, _19184_);
  or (_19186_, _19185_, _19087_);
  or (_19187_, _19186_, _19183_);
  or (_19188_, _19109_, word_in[30]);
  and (_36792_, _19188_, _19187_);
  and (_19189_, _18785_, word_in[7]);
  and (_19190_, _19189_, _18817_);
  and (_19191_, _19094_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_19192_, _19191_, _19190_);
  nor (_19193_, _19192_, _19093_);
  and (_19194_, _19093_, word_in[15]);
  nor (_19195_, _19194_, _19193_);
  nor (_19196_, _19195_, _19092_);
  and (_19197_, _19092_, _18795_);
  or (_19198_, _19197_, _19087_);
  or (_19199_, _19198_, _19196_);
  or (_19200_, _19109_, word_in[31]);
  and (_36793_, _19200_, _19199_);
  and (_19201_, _18767_, _18404_);
  and (_19202_, _19201_, _18977_);
  not (_19203_, _19202_);
  not (_19204_, _18773_);
  and (_19205_, _18980_, _19204_);
  and (_19206_, _19205_, _18617_);
  and (_19207_, _18780_, _18817_);
  and (_19208_, _19096_, _18807_);
  nand (_19209_, _18785_, _18807_);
  and (_19210_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_19211_, _19210_, _19208_);
  nor (_19212_, _19211_, _19207_);
  and (_19213_, _19207_, word_in[8]);
  nor (_19214_, _19213_, _19212_);
  nor (_19215_, _19214_, _19206_);
  and (_19216_, _19206_, _19104_);
  or (_19217_, _19216_, _19215_);
  and (_19218_, _19217_, _19203_);
  and (_19219_, _19202_, word_in[24]);
  or (_36794_, _19219_, _19218_);
  and (_19220_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_19221_, _19112_, _18807_);
  nor (_19222_, _19221_, _19220_);
  nor (_19223_, _19222_, _19207_);
  and (_19224_, _19207_, word_in[9]);
  nor (_19225_, _19224_, _19223_);
  nor (_19226_, _19225_, _19206_);
  and (_19227_, _19206_, _19119_);
  or (_19228_, _19227_, _19226_);
  and (_19229_, _19228_, _19203_);
  and (_19230_, _19202_, word_in[25]);
  or (_36795_, _19230_, _19229_);
  and (_19231_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_19232_, _19125_, _18807_);
  nor (_19233_, _19232_, _19231_);
  nor (_19234_, _19233_, _19207_);
  and (_19235_, _19207_, word_in[10]);
  nor (_19236_, _19235_, _19234_);
  nor (_19237_, _19236_, _19206_);
  and (_19238_, _19206_, _19132_);
  or (_19239_, _19238_, _19237_);
  and (_19240_, _19239_, _19203_);
  and (_19241_, _19202_, word_in[26]);
  or (_36796_, _19241_, _19240_);
  and (_19242_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_19243_, _19137_, _18807_);
  nor (_19244_, _19243_, _19242_);
  nor (_19245_, _19244_, _19207_);
  and (_19246_, _19207_, word_in[11]);
  nor (_19247_, _19246_, _19245_);
  nor (_19248_, _19247_, _19206_);
  and (_19249_, _19206_, _19145_);
  or (_19250_, _19249_, _19248_);
  and (_19251_, _19250_, _19203_);
  and (_19252_, _19202_, word_in[27]);
  or (_36797_, _19252_, _19251_);
  and (_19253_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_19254_, _19151_, _18807_);
  or (_19255_, _19254_, _19253_);
  or (_19256_, _19255_, _19207_);
  not (_19257_, word_in[12]);
  nand (_19258_, _19207_, _19257_);
  nand (_19259_, _19258_, _19256_);
  nor (_19260_, _19259_, _19206_);
  and (_19261_, _19206_, _19158_);
  or (_19262_, _19261_, _19260_);
  or (_19263_, _19262_, _19202_);
  or (_19264_, _19203_, word_in[28]);
  and (_36798_, _19264_, _19263_);
  and (_19265_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_19266_, _19163_, _18807_);
  nor (_19267_, _19266_, _19265_);
  nor (_19268_, _19267_, _19207_);
  and (_19269_, _19207_, word_in[13]);
  nor (_19270_, _19269_, _19268_);
  nor (_19271_, _19270_, _19206_);
  and (_19272_, _19206_, _19171_);
  or (_19273_, _19272_, _19271_);
  and (_19274_, _19273_, _19203_);
  and (_19275_, _19202_, word_in[29]);
  or (_36799_, _19275_, _19274_);
  and (_19276_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_19277_, _19177_, _18807_);
  nor (_19278_, _19277_, _19276_);
  nor (_19279_, _19278_, _19207_);
  and (_19280_, _19207_, word_in[14]);
  nor (_19281_, _19280_, _19279_);
  nor (_19282_, _19281_, _19206_);
  and (_19283_, _19206_, _19184_);
  or (_19284_, _19283_, _19282_);
  and (_19285_, _19284_, _19203_);
  and (_19286_, _19202_, word_in[30]);
  or (_36800_, _19286_, _19285_);
  and (_19287_, _19209_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_19288_, _19189_, _18807_);
  nor (_19289_, _19288_, _19287_);
  nor (_19290_, _19289_, _19207_);
  and (_19291_, _19207_, word_in[15]);
  nor (_19292_, _19291_, _19290_);
  nor (_19293_, _19292_, _19206_);
  and (_19294_, _19206_, _18795_);
  or (_19295_, _19294_, _19293_);
  and (_19296_, _19295_, _19203_);
  and (_19297_, _19202_, word_in[31]);
  or (_36801_, _19297_, _19296_);
  and (_19298_, _18767_, _18799_);
  not (_19299_, _19298_);
  not (_19300_, _18774_);
  nor (_19301_, _19089_, _19300_);
  and (_19302_, _18780_, _18807_);
  nand (_19303_, _18785_, _18816_);
  and (_19304_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_19305_, _19096_, _18816_);
  nor (_19306_, _19305_, _19304_);
  nor (_19307_, _19306_, _19302_);
  and (_19308_, _19302_, word_in[8]);
  nor (_19309_, _19308_, _19307_);
  nor (_19310_, _19309_, _19301_);
  and (_19311_, _19301_, _19104_);
  or (_19312_, _19311_, _19310_);
  and (_19313_, _19312_, _19299_);
  and (_19314_, _19298_, word_in[24]);
  or (_36802_, _19314_, _19313_);
  and (_19315_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_19316_, _19112_, _18816_);
  nor (_19317_, _19316_, _19315_);
  nor (_19318_, _19317_, _19302_);
  and (_19319_, _19302_, word_in[9]);
  nor (_19320_, _19319_, _19318_);
  nor (_19321_, _19320_, _19301_);
  and (_19322_, _19301_, _19119_);
  or (_19323_, _19322_, _19321_);
  and (_19324_, _19323_, _19299_);
  and (_19325_, _19298_, word_in[25]);
  or (_36803_, _19325_, _19324_);
  and (_19326_, _19125_, _18816_);
  and (_19327_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_19328_, _19327_, _19326_);
  nor (_19329_, _19328_, _19302_);
  and (_19330_, _19302_, word_in[10]);
  nor (_19331_, _19330_, _19329_);
  nor (_19332_, _19331_, _19301_);
  and (_19333_, _19301_, _19132_);
  or (_19334_, _19333_, _19332_);
  and (_19335_, _19334_, _19299_);
  and (_19336_, _19298_, word_in[26]);
  or (_36804_, _19336_, _19335_);
  and (_19337_, _19137_, _18816_);
  and (_19338_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_19339_, _19338_, _19337_);
  nor (_19340_, _19339_, _19302_);
  and (_19341_, _19302_, word_in[11]);
  nor (_19342_, _19341_, _19340_);
  nor (_19343_, _19342_, _19301_);
  and (_19344_, _19301_, _19145_);
  or (_19345_, _19344_, _19343_);
  and (_19346_, _19345_, _19299_);
  and (_19347_, _19298_, word_in[27]);
  or (_36805_, _19347_, _19346_);
  and (_19348_, _19298_, _19038_);
  and (_19349_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_19350_, _19151_, _18816_);
  or (_19351_, _19350_, _19349_);
  or (_19352_, _19351_, _19302_);
  nand (_19353_, _19302_, _19257_);
  and (_19354_, _19353_, _19352_);
  or (_19355_, _19354_, _19301_);
  not (_19356_, _19301_);
  or (_19357_, _19356_, _19158_);
  and (_19358_, _19357_, _19299_);
  and (_19359_, _19358_, _19355_);
  or (_36806_, _19359_, _19348_);
  and (_19360_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_19361_, _19163_, _18816_);
  nor (_19362_, _19361_, _19360_);
  nor (_19363_, _19362_, _19302_);
  and (_19364_, _19302_, word_in[13]);
  nor (_19365_, _19364_, _19363_);
  nor (_19366_, _19365_, _19301_);
  and (_19367_, _19301_, _19171_);
  or (_19368_, _19367_, _19366_);
  and (_19369_, _19368_, _19299_);
  and (_19370_, _19298_, word_in[29]);
  or (_36807_, _19370_, _19369_);
  and (_19371_, _19177_, _18816_);
  and (_19372_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_19373_, _19372_, _19371_);
  nor (_19374_, _19373_, _19302_);
  and (_19375_, _19302_, word_in[14]);
  nor (_19376_, _19375_, _19374_);
  nor (_19377_, _19376_, _19301_);
  and (_19378_, _19301_, _19184_);
  or (_19379_, _19378_, _19377_);
  and (_19380_, _19379_, _19299_);
  and (_19381_, _19298_, word_in[30]);
  or (_36808_, _19381_, _19380_);
  and (_19382_, _19189_, _18816_);
  and (_19383_, _19303_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  or (_19384_, _19383_, _19382_);
  or (_19385_, _19384_, _19302_);
  not (_19386_, word_in[15]);
  nand (_19387_, _19302_, _19386_);
  and (_19388_, _19387_, _19385_);
  or (_19389_, _19388_, _19301_);
  or (_19390_, _19356_, _18795_);
  and (_19391_, _19390_, _19389_);
  or (_19392_, _19391_, _19298_);
  or (_19393_, _19299_, word_in[31]);
  and (_36809_, _19393_, _19392_);
  and (_19394_, _18975_, _18752_);
  and (_19395_, _19394_, _18426_);
  not (_19396_, _19395_);
  not (_19397_, _18916_);
  and (_19398_, _19397_, _18776_);
  and (_19399_, _19398_, _18981_);
  and (_19400_, _18781_, _18504_);
  and (_19401_, _19400_, _18404_);
  nand (_19402_, _18785_, _18811_);
  and (_19403_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_19404_, _19096_, _18811_);
  nor (_19405_, _19404_, _19403_);
  nor (_19406_, _19405_, _19401_);
  and (_19407_, _18780_, word_in[8]);
  and (_19408_, _19401_, _19407_);
  nor (_19409_, _19408_, _19406_);
  nor (_19410_, _19409_, _19399_);
  and (_19411_, _19399_, _19104_);
  or (_19412_, _19411_, _19410_);
  and (_19413_, _19412_, _19396_);
  and (_19414_, _18767_, word_in[24]);
  and (_19415_, _19395_, _19414_);
  or (_36810_, _19415_, _19413_);
  and (_19416_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_19417_, _19112_, _18811_);
  nor (_19418_, _19417_, _19416_);
  nor (_19419_, _19418_, _19401_);
  and (_19420_, _19401_, _19001_);
  nor (_19421_, _19420_, _19419_);
  nor (_19422_, _19421_, _19399_);
  and (_19423_, _19399_, _19119_);
  or (_19424_, _19423_, _19422_);
  and (_19425_, _19424_, _19396_);
  and (_19426_, _18767_, word_in[25]);
  and (_19427_, _19395_, _19426_);
  or (_36811_, _19427_, _19425_);
  and (_19428_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_19429_, _19125_, _18811_);
  nor (_19430_, _19429_, _19428_);
  nor (_19431_, _19430_, _19401_);
  and (_19432_, _18780_, word_in[10]);
  and (_19433_, _19401_, _19432_);
  nor (_19434_, _19433_, _19431_);
  nor (_19435_, _19434_, _19399_);
  and (_19436_, _19399_, _19132_);
  or (_19437_, _19436_, _19395_);
  or (_19438_, _19437_, _19435_);
  and (_19439_, _18767_, word_in[26]);
  or (_19440_, _19396_, _19439_);
  and (_36812_, _19440_, _19438_);
  and (_19441_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_19442_, _19137_, _18811_);
  nor (_19443_, _19442_, _19441_);
  nor (_19444_, _19443_, _19401_);
  and (_19445_, _18780_, word_in[11]);
  and (_19446_, _19401_, _19445_);
  nor (_19447_, _19446_, _19444_);
  nor (_19448_, _19447_, _19399_);
  and (_19449_, _19399_, _19145_);
  or (_19450_, _19449_, _19448_);
  and (_19451_, _19450_, _19396_);
  and (_19452_, _18767_, word_in[27]);
  and (_19453_, _19395_, _19452_);
  or (_36813_, _19453_, _19451_);
  and (_19454_, _18780_, word_in[12]);
  not (_19455_, _19401_);
  or (_19456_, _19455_, _19454_);
  and (_19457_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_19458_, _19151_, _18811_);
  or (_19459_, _19458_, _19457_);
  or (_19460_, _19459_, _19401_);
  and (_19461_, _19460_, _19456_);
  or (_19462_, _19461_, _19399_);
  not (_19463_, _19399_);
  or (_19464_, _19463_, _19158_);
  and (_19465_, _19464_, _19396_);
  and (_19466_, _19465_, _19462_);
  and (_19467_, _19395_, _19038_);
  or (_36814_, _19467_, _19466_);
  and (_19468_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_19469_, _19163_, _18811_);
  nor (_19470_, _19469_, _19468_);
  nor (_19471_, _19470_, _19401_);
  and (_19472_, _18780_, word_in[13]);
  and (_19473_, _19401_, _19472_);
  nor (_19474_, _19473_, _19471_);
  nor (_19475_, _19474_, _19399_);
  and (_19476_, _19399_, _19171_);
  or (_19477_, _19476_, _19475_);
  and (_19478_, _19477_, _19396_);
  and (_19479_, _18767_, word_in[29]);
  and (_19480_, _19395_, _19479_);
  or (_36815_, _19480_, _19478_);
  and (_19481_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_19482_, _19177_, _18811_);
  nor (_19483_, _19482_, _19481_);
  nor (_19484_, _19483_, _19401_);
  and (_19485_, _18780_, word_in[14]);
  and (_19486_, _19401_, _19485_);
  nor (_19487_, _19486_, _19484_);
  nor (_19488_, _19487_, _19399_);
  and (_19489_, _19399_, _19184_);
  or (_19490_, _19489_, _19488_);
  and (_19491_, _19490_, _19396_);
  and (_19492_, _18767_, word_in[30]);
  and (_19493_, _19395_, _19492_);
  or (_36816_, _19493_, _19491_);
  or (_19494_, _19455_, _18791_);
  and (_19495_, _19402_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_19496_, _19189_, _18811_);
  or (_19497_, _19496_, _19495_);
  or (_19498_, _19497_, _19401_);
  and (_19499_, _19498_, _19494_);
  or (_19500_, _19499_, _19399_);
  or (_19501_, _19463_, _18795_);
  and (_19502_, _19501_, _19396_);
  and (_19503_, _19502_, _19500_);
  and (_19504_, _19395_, _18768_);
  or (_36857_[7], _19504_, _19503_);
  and (_19505_, _19398_, _19090_);
  and (_19506_, _19400_, _18414_);
  and (_19507_, _19096_, _18824_);
  nand (_19508_, _18785_, _18824_);
  and (_19509_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or (_19510_, _19509_, _19507_);
  or (_19511_, _19510_, _19506_);
  not (_19512_, _19506_);
  or (_19513_, _19512_, _19407_);
  and (_19514_, _19513_, _19511_);
  or (_19515_, _19514_, _19505_);
  and (_19516_, _19394_, _18437_);
  not (_19517_, _19516_);
  not (_19518_, _19505_);
  or (_19519_, _19518_, _19104_);
  and (_19520_, _19519_, _19517_);
  and (_19521_, _19520_, _19515_);
  and (_19522_, _19516_, _19414_);
  or (_36817_, _19522_, _19521_);
  and (_19523_, _19112_, _18824_);
  and (_19524_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  or (_19525_, _19524_, _19523_);
  or (_19526_, _19525_, _19506_);
  or (_19527_, _19512_, _19001_);
  and (_19528_, _19527_, _19526_);
  or (_19529_, _19528_, _19505_);
  or (_19530_, _19518_, _19119_);
  and (_19531_, _19530_, _19517_);
  and (_19532_, _19531_, _19529_);
  and (_19533_, _19516_, _19426_);
  or (_36818_, _19533_, _19532_);
  and (_19534_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_19535_, _19125_, _18824_);
  nor (_19536_, _19535_, _19534_);
  nor (_19537_, _19536_, _19506_);
  and (_19538_, _19506_, _19432_);
  or (_19539_, _19538_, _19537_);
  and (_19540_, _19539_, _19518_);
  and (_19541_, _19505_, _19132_);
  or (_19542_, _19541_, _19516_);
  or (_19543_, _19542_, _19540_);
  or (_19544_, _19517_, _19439_);
  and (_36819_, _19544_, _19543_);
  and (_19545_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_19546_, _19137_, _18824_);
  nor (_19547_, _19546_, _19545_);
  nor (_19548_, _19547_, _19506_);
  and (_19549_, _19506_, _19445_);
  or (_19550_, _19549_, _19548_);
  and (_19551_, _19550_, _19518_);
  and (_19552_, _19505_, _19145_);
  or (_19553_, _19552_, _19516_);
  or (_19554_, _19553_, _19551_);
  or (_19555_, _19517_, _19452_);
  and (_36820_, _19555_, _19554_);
  and (_19556_, _19505_, _19158_);
  and (_19557_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_19558_, _19151_, _18824_);
  nor (_19559_, _19558_, _19557_);
  nor (_19560_, _19559_, _19506_);
  and (_19561_, _19506_, _19454_);
  or (_19562_, _19561_, _19560_);
  and (_19563_, _19562_, _19518_);
  or (_19564_, _19563_, _19556_);
  and (_19565_, _19564_, _19517_);
  and (_19566_, _19516_, _19038_);
  or (_36821_, _19566_, _19565_);
  and (_19567_, _19505_, _19171_);
  and (_19568_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_19569_, _19163_, _18824_);
  nor (_19570_, _19569_, _19568_);
  nor (_19571_, _19570_, _19506_);
  and (_19572_, _19506_, _19472_);
  or (_19573_, _19572_, _19571_);
  and (_19574_, _19573_, _19518_);
  or (_19575_, _19574_, _19567_);
  and (_19576_, _19575_, _19517_);
  and (_19577_, _19516_, _19479_);
  or (_36822_, _19577_, _19576_);
  and (_19578_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_19579_, _19177_, _18824_);
  nor (_19580_, _19579_, _19578_);
  nor (_19581_, _19580_, _19506_);
  and (_19582_, _19506_, _19485_);
  or (_19583_, _19582_, _19581_);
  and (_19584_, _19583_, _19518_);
  and (_19585_, _19505_, _19184_);
  or (_19586_, _19585_, _19516_);
  or (_19587_, _19586_, _19584_);
  or (_19588_, _19517_, _19492_);
  and (_36823_, _19588_, _19587_);
  and (_19589_, _19508_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_19590_, _19189_, _18824_);
  nor (_19591_, _19590_, _19589_);
  nor (_19592_, _19591_, _19506_);
  and (_19593_, _19506_, _18791_);
  or (_19594_, _19593_, _19592_);
  and (_19595_, _19594_, _19518_);
  and (_19596_, _19505_, _18795_);
  or (_19597_, _19596_, _19516_);
  or (_19598_, _19597_, _19595_);
  or (_19599_, _19517_, _18768_);
  and (_36824_, _19599_, _19598_);
  and (_19600_, _19205_, _19397_);
  and (_19601_, _19400_, _18426_);
  and (_19602_, _18785_, _18847_);
  and (_19603_, _19602_, word_in[0]);
  not (_19604_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_19605_, _19602_, _19604_);
  nor (_19606_, _19605_, _19603_);
  nor (_19607_, _19606_, _19601_);
  and (_19608_, _19601_, _19407_);
  or (_19609_, _19608_, _19607_);
  or (_19610_, _19609_, _19600_);
  and (_19611_, _19394_, _18404_);
  not (_19612_, _19611_);
  not (_19613_, _19600_);
  or (_19614_, _19613_, _19104_);
  and (_19615_, _19614_, _19612_);
  and (_19616_, _19615_, _19610_);
  and (_19617_, _19611_, _19414_);
  or (_36825_, _19617_, _19616_);
  not (_19618_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_19619_, _19602_, _19618_);
  and (_19620_, _19602_, _19112_);
  or (_19621_, _19620_, _19619_);
  or (_19622_, _19621_, _19601_);
  not (_19623_, _19601_);
  or (_19624_, _19623_, _19001_);
  and (_19625_, _19624_, _19622_);
  or (_19626_, _19625_, _19600_);
  or (_19627_, _19613_, _19119_);
  and (_19628_, _19627_, _19612_);
  and (_19629_, _19628_, _19626_);
  and (_19630_, _19611_, _19426_);
  or (_36826_, _19630_, _19629_);
  and (_19631_, _19602_, word_in[2]);
  not (_19632_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_19633_, _19602_, _19632_);
  nor (_19634_, _19633_, _19631_);
  nor (_19635_, _19634_, _19601_);
  and (_19636_, _19601_, _19432_);
  nor (_19637_, _19636_, _19635_);
  nor (_19638_, _19637_, _19600_);
  and (_19639_, _19600_, _19132_);
  or (_19640_, _19639_, _19611_);
  or (_19641_, _19640_, _19638_);
  or (_19642_, _19612_, _19439_);
  and (_36827_, _19642_, _19641_);
  and (_19643_, _19600_, _19145_);
  and (_19644_, _19602_, word_in[3]);
  not (_19645_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_19646_, _19602_, _19645_);
  nor (_19647_, _19646_, _19644_);
  nor (_19648_, _19647_, _19601_);
  and (_19649_, _19601_, _19445_);
  nor (_19650_, _19649_, _19648_);
  nor (_19651_, _19650_, _19600_);
  or (_19652_, _19651_, _19643_);
  and (_19653_, _19652_, _19612_);
  and (_19654_, _19611_, _19452_);
  or (_36828_, _19654_, _19653_);
  and (_19655_, _19600_, _19158_);
  and (_19656_, _19602_, word_in[4]);
  not (_19657_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_19658_, _19602_, _19657_);
  nor (_19659_, _19658_, _19656_);
  nor (_19660_, _19659_, _19601_);
  and (_19661_, _19601_, _19454_);
  nor (_19662_, _19661_, _19660_);
  nor (_19663_, _19662_, _19600_);
  or (_19664_, _19663_, _19655_);
  and (_19665_, _19664_, _19612_);
  and (_19666_, _19611_, _19038_);
  or (_36829_, _19666_, _19665_);
  not (_19667_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_19668_, _19602_, _19667_);
  and (_19669_, _19602_, _19163_);
  or (_19670_, _19669_, _19668_);
  or (_19671_, _19670_, _19601_);
  or (_19672_, _19623_, _19472_);
  and (_19673_, _19672_, _19671_);
  or (_19674_, _19673_, _19600_);
  or (_19675_, _19613_, _19171_);
  and (_19676_, _19675_, _19612_);
  and (_19677_, _19676_, _19674_);
  and (_19678_, _19611_, _19479_);
  or (_36830_, _19678_, _19677_);
  not (_19679_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_19680_, _19602_, _19679_);
  and (_19681_, _19602_, _19177_);
  or (_19682_, _19681_, _19680_);
  or (_19683_, _19682_, _19601_);
  or (_19684_, _19623_, _19485_);
  and (_19685_, _19684_, _19683_);
  or (_19686_, _19685_, _19600_);
  or (_19687_, _19613_, _19184_);
  and (_19688_, _19687_, _19612_);
  and (_19689_, _19688_, _19686_);
  and (_19690_, _19611_, _19492_);
  or (_36831_, _19690_, _19689_);
  and (_19691_, _19602_, word_in[7]);
  nor (_19692_, _19602_, _18572_);
  nor (_19693_, _19692_, _19691_);
  nor (_19694_, _19693_, _19601_);
  and (_19695_, _19601_, _18791_);
  nor (_19696_, _19695_, _19694_);
  nor (_19697_, _19696_, _19600_);
  and (_19698_, _19600_, _18795_);
  or (_19699_, _19698_, _19697_);
  and (_19700_, _19699_, _19612_);
  and (_19701_, _19611_, _18768_);
  or (_36832_, _19701_, _19700_);
  and (_19702_, _18767_, _18811_);
  and (_19703_, _19398_, _18774_);
  and (_19704_, _19400_, _18437_);
  not (_19705_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_19706_, _18785_, _18503_);
  nor (_19707_, _19706_, _19705_);
  and (_19708_, _19706_, _19096_);
  or (_19709_, _19708_, _19707_);
  or (_19710_, _19709_, _19704_);
  not (_19711_, _19704_);
  or (_19712_, _19711_, _19407_);
  and (_19713_, _19712_, _19710_);
  or (_19714_, _19713_, _19703_);
  not (_19715_, _19703_);
  or (_19716_, _19715_, word_in[16]);
  and (_19717_, _19716_, _19714_);
  or (_19718_, _19717_, _19702_);
  not (_19719_, _19702_);
  or (_19720_, _19719_, word_in[24]);
  and (_36833_, _19720_, _19718_);
  not (_19721_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_19722_, _19706_, _19721_);
  and (_19723_, _19706_, word_in[1]);
  nor (_19724_, _19723_, _19722_);
  nor (_19725_, _19724_, _19704_);
  and (_19726_, _19704_, _19001_);
  or (_19727_, _19726_, _19725_);
  and (_19728_, _19727_, _19715_);
  and (_19729_, _19703_, word_in[17]);
  or (_19730_, _19729_, _19728_);
  and (_19731_, _19730_, _19719_);
  and (_19732_, _19702_, word_in[25]);
  or (_36834_, _19732_, _19731_);
  and (_19733_, _19702_, word_in[26]);
  and (_19734_, _19706_, word_in[2]);
  not (_19735_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_19736_, _19706_, _19735_);
  nor (_19737_, _19736_, _19734_);
  nor (_19738_, _19737_, _19704_);
  and (_19739_, _19704_, _19432_);
  or (_19740_, _19739_, _19738_);
  and (_19741_, _19740_, _19715_);
  and (_19742_, _19703_, word_in[18]);
  or (_19743_, _19742_, _19741_);
  and (_19744_, _19743_, _19719_);
  or (_36835_, _19744_, _19733_);
  not (_19745_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_19746_, _19706_, _19745_);
  and (_19747_, _19706_, _19137_);
  or (_19748_, _19747_, _19746_);
  or (_19749_, _19748_, _19704_);
  or (_19750_, _19711_, _19445_);
  and (_19751_, _19750_, _19749_);
  or (_19752_, _19751_, _19703_);
  or (_19753_, _19715_, _19145_);
  and (_19754_, _19753_, _19719_);
  and (_19755_, _19754_, _19752_);
  and (_19756_, _19702_, word_in[27]);
  or (_36836_, _19756_, _19755_);
  and (_19757_, _19038_, _18811_);
  and (_19758_, _19706_, word_in[4]);
  not (_19759_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_19760_, _19706_, _19759_);
  nor (_19761_, _19760_, _19758_);
  nor (_19762_, _19761_, _19704_);
  and (_19763_, _19704_, _19454_);
  or (_19764_, _19763_, _19762_);
  or (_19765_, _19764_, _19703_);
  or (_19766_, _19715_, _19158_);
  and (_19767_, _19766_, _19719_);
  and (_19768_, _19767_, _19765_);
  or (_36837_, _19768_, _19757_);
  and (_19769_, _19706_, word_in[5]);
  not (_19770_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_19771_, _19706_, _19770_);
  nor (_19772_, _19771_, _19769_);
  nor (_19773_, _19772_, _19704_);
  and (_19774_, _19704_, _19472_);
  or (_19775_, _19774_, _19773_);
  and (_19776_, _19775_, _19715_);
  and (_19777_, _19703_, word_in[21]);
  or (_19778_, _19777_, _19776_);
  and (_19779_, _19778_, _19719_);
  and (_19780_, _19702_, word_in[29]);
  or (_36838_, _19780_, _19779_);
  and (_19781_, _19702_, word_in[30]);
  not (_19782_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_19783_, _19706_, _19782_);
  and (_19784_, _19706_, _19177_);
  or (_19785_, _19784_, _19783_);
  or (_19786_, _19785_, _19704_);
  or (_19787_, _19711_, _19485_);
  and (_19788_, _19787_, _19786_);
  or (_19789_, _19788_, _19703_);
  or (_19790_, _19715_, word_in[22]);
  and (_19791_, _19790_, _19719_);
  and (_19792_, _19791_, _19789_);
  or (_36839_, _19792_, _19781_);
  and (_19793_, _19702_, word_in[31]);
  and (_19794_, _19706_, word_in[7]);
  nor (_19795_, _19706_, _18451_);
  nor (_19796_, _19795_, _19794_);
  nor (_19797_, _19796_, _19704_);
  and (_19798_, _19704_, _18791_);
  or (_19799_, _19798_, _19797_);
  and (_19800_, _19799_, _19715_);
  and (_19801_, _19703_, word_in[23]);
  or (_19802_, _19801_, _19800_);
  and (_19803_, _19802_, _19719_);
  or (_36840_, _19803_, _19793_);
  and (_19804_, _18777_, _18616_);
  and (_19805_, _19804_, _18981_);
  and (_19806_, _18780_, _18503_);
  not (_19807_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_19808_, _18785_, _18905_);
  nor (_19809_, _19808_, _19807_);
  and (_19810_, _19808_, _19096_);
  or (_19811_, _19810_, _19809_);
  or (_19812_, _19811_, _19806_);
  not (_19813_, _19806_);
  or (_19814_, _19813_, word_in[8]);
  nand (_19815_, _19814_, _19812_);
  nor (_19816_, _19815_, _19805_);
  and (_19817_, _18976_, _18700_);
  and (_19818_, _19817_, _18426_);
  and (_19819_, _19805_, _19104_);
  or (_19820_, _19819_, _19818_);
  or (_19821_, _19820_, _19816_);
  not (_19822_, _19818_);
  or (_19823_, _19822_, _19414_);
  and (_36841_, _19823_, _19821_);
  and (_19824_, _19808_, word_in[1]);
  not (_19825_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_19826_, _19808_, _19825_);
  nor (_19827_, _19826_, _19824_);
  nor (_19828_, _19827_, _19806_);
  and (_19829_, _19806_, word_in[9]);
  nor (_19830_, _19829_, _19828_);
  nor (_19831_, _19830_, _19805_);
  and (_19832_, _19805_, _19119_);
  or (_19833_, _19832_, _19831_);
  and (_19834_, _19833_, _19822_);
  and (_19835_, _19818_, _19426_);
  or (_36842_, _19835_, _19834_);
  and (_19836_, _19808_, word_in[2]);
  not (_19837_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_19838_, _19808_, _19837_);
  nor (_19839_, _19838_, _19836_);
  nor (_19840_, _19839_, _19806_);
  and (_19841_, _19806_, word_in[10]);
  nor (_19842_, _19841_, _19840_);
  nor (_19843_, _19842_, _19805_);
  and (_19844_, _19805_, _19132_);
  or (_19845_, _19844_, _19843_);
  and (_19846_, _19845_, _19822_);
  and (_19847_, _19818_, _19439_);
  or (_36843_, _19847_, _19846_);
  and (_19848_, _19808_, word_in[3]);
  not (_19849_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_19850_, _19808_, _19849_);
  nor (_19851_, _19850_, _19848_);
  nor (_19852_, _19851_, _19806_);
  and (_19853_, _19806_, word_in[11]);
  nor (_19854_, _19853_, _19852_);
  nor (_19855_, _19854_, _19805_);
  and (_19856_, _19805_, _19145_);
  or (_19857_, _19856_, _19855_);
  and (_19858_, _19857_, _19822_);
  and (_19859_, _19818_, _19452_);
  or (_36844_, _19859_, _19858_);
  not (_19860_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_19861_, _19808_, _19860_);
  and (_19862_, _19808_, _19151_);
  or (_19863_, _19862_, _19861_);
  or (_19864_, _19863_, _19806_);
  nand (_19865_, _19806_, _19257_);
  nand (_19866_, _19865_, _19864_);
  nor (_19867_, _19866_, _19805_);
  and (_19868_, _19805_, _19158_);
  or (_19869_, _19868_, _19867_);
  or (_19870_, _19869_, _19818_);
  or (_19871_, _19822_, _19038_);
  and (_36845_, _19871_, _19870_);
  and (_19872_, _19808_, word_in[5]);
  not (_19873_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_19874_, _19808_, _19873_);
  nor (_19875_, _19874_, _19872_);
  nor (_19876_, _19875_, _19806_);
  and (_19877_, _19806_, word_in[13]);
  nor (_19878_, _19877_, _19876_);
  nor (_19879_, _19878_, _19805_);
  and (_19880_, _19805_, _19171_);
  or (_19881_, _19880_, _19879_);
  and (_19882_, _19881_, _19822_);
  and (_19883_, _19818_, _19479_);
  or (_36846_, _19883_, _19882_);
  and (_19884_, _19808_, word_in[6]);
  not (_19885_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_19886_, _19808_, _19885_);
  nor (_19887_, _19886_, _19884_);
  nor (_19888_, _19887_, _19806_);
  and (_19889_, _19806_, word_in[14]);
  nor (_19890_, _19889_, _19888_);
  nor (_19891_, _19890_, _19805_);
  and (_19892_, _19805_, _19184_);
  or (_19893_, _19892_, _19891_);
  and (_19894_, _19893_, _19822_);
  and (_19895_, _19818_, _19492_);
  or (_36847_, _19895_, _19894_);
  and (_19896_, _19808_, word_in[7]);
  nor (_19897_, _19808_, _18581_);
  nor (_19898_, _19897_, _19896_);
  nor (_19899_, _19898_, _19806_);
  and (_19900_, _19806_, word_in[15]);
  nor (_19901_, _19900_, _19899_);
  nor (_19902_, _19901_, _19805_);
  and (_19903_, _19805_, _18795_);
  or (_19904_, _19903_, _19902_);
  and (_19905_, _19904_, _19822_);
  and (_19906_, _19818_, _18768_);
  or (_36848_, _19906_, _19905_);
  and (_19907_, _19817_, _18437_);
  not (_19908_, _19907_);
  and (_19909_, _19804_, _19090_);
  and (_19910_, _18780_, _18513_);
  and (_19911_, _19910_, _18414_);
  and (_19912_, _19096_, _18888_);
  not (_19913_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_19914_, _18785_, _18888_);
  nor (_19915_, _19914_, _19913_);
  nor (_19916_, _19915_, _19912_);
  nor (_19917_, _19916_, _19911_);
  and (_19918_, _19911_, _19407_);
  nor (_19919_, _19918_, _19917_);
  nor (_19920_, _19919_, _19909_);
  and (_19921_, _19909_, _19104_);
  or (_19922_, _19921_, _19920_);
  and (_19923_, _19922_, _19908_);
  and (_19924_, _19907_, _19414_);
  or (_36849_, _19924_, _19923_);
  not (_19925_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_19926_, _19914_, _19925_);
  and (_19927_, _19112_, _18888_);
  nor (_19928_, _19927_, _19926_);
  nor (_19929_, _19928_, _19911_);
  and (_19930_, _19911_, _19001_);
  nor (_19931_, _19930_, _19929_);
  nor (_19932_, _19931_, _19909_);
  and (_19933_, _19909_, _19119_);
  or (_19934_, _19933_, _19932_);
  and (_19935_, _19934_, _19908_);
  and (_19936_, _19907_, _19426_);
  or (_36850_, _19936_, _19935_);
  not (_19937_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_19938_, _19914_, _19937_);
  and (_19939_, _19125_, _18888_);
  or (_19940_, _19939_, _19938_);
  or (_19941_, _19940_, _19911_);
  not (_19942_, _19911_);
  or (_19943_, _19942_, _19432_);
  and (_19944_, _19943_, _19941_);
  or (_19945_, _19944_, _19909_);
  not (_19946_, _19909_);
  or (_19947_, _19946_, _19132_);
  and (_19948_, _19947_, _19945_);
  or (_19949_, _19948_, _19907_);
  or (_19950_, _19908_, _19439_);
  and (_36851_, _19950_, _19949_);
  not (_19951_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_19952_, _19914_, _19951_);
  and (_19953_, _19137_, _18888_);
  nor (_19954_, _19953_, _19952_);
  nor (_19955_, _19954_, _19911_);
  and (_19956_, _19911_, _19445_);
  nor (_19957_, _19956_, _19955_);
  nor (_19958_, _19957_, _19909_);
  and (_19959_, _19909_, _19145_);
  or (_19960_, _19959_, _19907_);
  or (_19961_, _19960_, _19958_);
  or (_19962_, _19908_, _19452_);
  and (_36852_, _19962_, _19961_);
  not (_19963_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_19964_, _19914_, _19963_);
  and (_19965_, _19151_, _18888_);
  or (_19966_, _19965_, _19964_);
  or (_19967_, _19966_, _19911_);
  or (_19968_, _19942_, _19454_);
  and (_19969_, _19968_, _19967_);
  or (_19970_, _19969_, _19909_);
  or (_19971_, _19946_, _19158_);
  and (_19972_, _19971_, _19970_);
  or (_19973_, _19972_, _19907_);
  or (_19974_, _19908_, _19038_);
  and (_36853_, _19974_, _19973_);
  not (_19975_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_19976_, _19914_, _19975_);
  and (_19977_, _19163_, _18888_);
  or (_19978_, _19977_, _19976_);
  or (_19979_, _19978_, _19911_);
  or (_19980_, _19942_, _19472_);
  nand (_19981_, _19980_, _19979_);
  nor (_19982_, _19981_, _19909_);
  and (_19983_, _19909_, _19171_);
  or (_19984_, _19983_, _19907_);
  or (_19985_, _19984_, _19982_);
  or (_19986_, _19908_, _19479_);
  and (_36854_, _19986_, _19985_);
  and (_19987_, _19914_, word_in[6]);
  not (_19988_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_19989_, _19914_, _19988_);
  nor (_19990_, _19989_, _19987_);
  nor (_19991_, _19990_, _19911_);
  and (_19992_, _19911_, _19485_);
  nor (_19993_, _19992_, _19991_);
  nor (_19994_, _19993_, _19909_);
  and (_19995_, _19909_, _19184_);
  or (_19996_, _19995_, _19994_);
  and (_19997_, _19996_, _19908_);
  and (_19998_, _19907_, _19492_);
  or (_36855_, _19998_, _19997_);
  nor (_19999_, _19914_, _18472_);
  and (_20000_, _19914_, _19189_);
  or (_20001_, _20000_, _19999_);
  or (_20002_, _20001_, _19911_);
  or (_20003_, _19942_, _18791_);
  and (_20004_, _20003_, _20002_);
  or (_20005_, _20004_, _19909_);
  or (_20006_, _19946_, _18795_);
  and (_20007_, _20006_, _19908_);
  and (_20008_, _20007_, _20005_);
  and (_20009_, _19907_, _18768_);
  or (_36856_, _20009_, _20008_);
  and (_20010_, _18976_, _18499_);
  not (_20011_, _20010_);
  and (_20012_, _19804_, _19205_);
  and (_20013_, _19910_, _18426_);
  and (_20014_, _18785_, _18900_);
  and (_20015_, _20014_, _19096_);
  not (_20016_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_20017_, _20014_, _20016_);
  nor (_20018_, _20017_, _20015_);
  nor (_20019_, _20018_, _20013_);
  and (_20020_, _20013_, _19407_);
  nor (_20021_, _20020_, _20019_);
  nor (_20022_, _20021_, _20012_);
  and (_20023_, _20012_, _19104_);
  or (_20024_, _20023_, _20022_);
  and (_20025_, _20024_, _20011_);
  and (_20026_, _20010_, word_in[24]);
  or (_36738_, _20026_, _20025_);
  and (_20027_, _20014_, word_in[1]);
  not (_20028_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_20029_, _20014_, _20028_);
  nor (_20030_, _20029_, _20027_);
  nor (_20031_, _20030_, _20013_);
  and (_20032_, _20013_, _19001_);
  nor (_20033_, _20032_, _20031_);
  nor (_20034_, _20033_, _20012_);
  and (_20035_, _20012_, _19119_);
  or (_20036_, _20035_, _20010_);
  or (_20037_, _20036_, _20034_);
  or (_20038_, _20011_, _19426_);
  and (_36739_, _20038_, _20037_);
  and (_20039_, _20014_, word_in[2]);
  not (_20040_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_20041_, _20014_, _20040_);
  nor (_20042_, _20041_, _20039_);
  nor (_20043_, _20042_, _20013_);
  and (_20044_, _20013_, _19432_);
  nor (_20045_, _20044_, _20043_);
  nor (_20046_, _20045_, _20012_);
  and (_20047_, _20012_, _19132_);
  or (_20048_, _20047_, _20010_);
  or (_20049_, _20048_, _20046_);
  or (_20050_, _20011_, _19439_);
  and (_36740_, _20050_, _20049_);
  and (_20051_, _20014_, word_in[3]);
  not (_20052_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_20053_, _20014_, _20052_);
  nor (_20054_, _20053_, _20051_);
  nor (_20055_, _20054_, _20013_);
  and (_20056_, _20013_, _19445_);
  nor (_20057_, _20056_, _20055_);
  nor (_20058_, _20057_, _20012_);
  and (_20059_, _20012_, _19145_);
  or (_20060_, _20059_, _20058_);
  and (_20061_, _20060_, _20011_);
  and (_20062_, _20010_, word_in[27]);
  or (_36741_, _20062_, _20061_);
  and (_20063_, _20014_, word_in[4]);
  not (_20064_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_20065_, _20014_, _20064_);
  nor (_20066_, _20065_, _20063_);
  nor (_20067_, _20066_, _20013_);
  and (_20068_, _20013_, _19454_);
  nor (_20069_, _20068_, _20067_);
  nor (_20070_, _20069_, _20012_);
  and (_20071_, _20012_, _19158_);
  or (_20072_, _20071_, _20070_);
  and (_20073_, _20072_, _20011_);
  and (_20074_, _20010_, word_in[28]);
  or (_36742_, _20074_, _20073_);
  and (_20075_, _20014_, word_in[5]);
  not (_20076_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_20077_, _20014_, _20076_);
  nor (_20078_, _20077_, _20075_);
  nor (_20079_, _20078_, _20013_);
  and (_20080_, _20013_, _19472_);
  nor (_20081_, _20080_, _20079_);
  nor (_20082_, _20081_, _20012_);
  and (_20083_, _20012_, _19171_);
  or (_20084_, _20083_, _20082_);
  and (_20085_, _20084_, _20011_);
  and (_20086_, _20010_, word_in[29]);
  or (_36743_, _20086_, _20085_);
  not (_20087_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_20088_, _20014_, _20087_);
  and (_20089_, _20014_, word_in[6]);
  nor (_20090_, _20089_, _20088_);
  nor (_20091_, _20090_, _20013_);
  and (_20092_, _20013_, _19485_);
  nor (_20093_, _20092_, _20091_);
  nor (_20094_, _20093_, _20012_);
  and (_20095_, _20012_, _19184_);
  or (_20096_, _20095_, _20094_);
  and (_20097_, _20096_, _20011_);
  and (_20098_, _20010_, word_in[30]);
  or (_36744_, _20098_, _20097_);
  and (_20099_, _20014_, word_in[7]);
  nor (_20100_, _20014_, _18586_);
  nor (_20101_, _20100_, _20099_);
  nor (_20102_, _20101_, _20013_);
  and (_20103_, _20013_, _18791_);
  nor (_20104_, _20103_, _20102_);
  nor (_20105_, _20104_, _20012_);
  and (_20106_, _20012_, _18795_);
  or (_20107_, _20106_, _20010_);
  or (_20108_, _20107_, _20105_);
  or (_20109_, _20011_, _18768_);
  and (_36745_, _20109_, _20108_);
  and (_20110_, _18767_, _18905_);
  not (_20111_, _20110_);
  and (_20112_, _19804_, _18774_);
  and (_20113_, _19910_, _18437_);
  and (_20114_, _18785_, _18926_);
  and (_20115_, _20114_, word_in[0]);
  not (_20116_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_20117_, _20114_, _20116_);
  nor (_20118_, _20117_, _20115_);
  nor (_20119_, _20118_, _20113_);
  and (_20120_, _20113_, _19407_);
  nor (_20121_, _20120_, _20119_);
  nor (_20122_, _20121_, _20112_);
  and (_20123_, _20112_, _19104_);
  or (_20124_, _20123_, _20122_);
  and (_20125_, _20124_, _20111_);
  and (_20126_, _20110_, word_in[24]);
  or (_36746_, _20126_, _20125_);
  not (_20127_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_20128_, _20114_, _20127_);
  and (_20129_, _20114_, word_in[1]);
  or (_20130_, _20129_, _20128_);
  or (_20131_, _20130_, _20113_);
  not (_20132_, _20113_);
  or (_20133_, _20132_, _19001_);
  and (_20134_, _20133_, _20131_);
  or (_20135_, _20134_, _20112_);
  not (_20136_, _20112_);
  or (_20137_, _20136_, _19119_);
  and (_20138_, _20137_, _20111_);
  and (_20139_, _20138_, _20135_);
  and (_20140_, _20110_, word_in[25]);
  or (_36747_, _20140_, _20139_);
  and (_20141_, _20114_, word_in[2]);
  not (_20142_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_20143_, _20114_, _20142_);
  nor (_20144_, _20143_, _20141_);
  nor (_20145_, _20144_, _20113_);
  and (_20146_, _20113_, _19432_);
  nor (_20147_, _20146_, _20145_);
  nor (_20148_, _20147_, _20112_);
  and (_20149_, _20112_, _19132_);
  or (_20150_, _20149_, _20148_);
  and (_20151_, _20150_, _20111_);
  and (_20152_, _20110_, word_in[26]);
  or (_36748_, _20152_, _20151_);
  and (_20153_, _20114_, word_in[3]);
  not (_20154_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_20155_, _20114_, _20154_);
  nor (_20156_, _20155_, _20153_);
  nor (_20157_, _20156_, _20113_);
  and (_20158_, _20113_, _19445_);
  nor (_20159_, _20158_, _20157_);
  nor (_20160_, _20159_, _20112_);
  and (_20161_, _20112_, _19145_);
  or (_20162_, _20161_, _20160_);
  and (_20163_, _20162_, _20111_);
  and (_20164_, _20110_, word_in[27]);
  or (_36749_, _20164_, _20163_);
  not (_20165_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_20166_, _20114_, _20165_);
  and (_20167_, _20114_, word_in[4]);
  or (_20168_, _20167_, _20166_);
  or (_20169_, _20168_, _20113_);
  or (_20170_, _20132_, _19454_);
  and (_20171_, _20170_, _20169_);
  or (_20172_, _20171_, _20112_);
  or (_20173_, _20136_, _19158_);
  and (_20174_, _20173_, _20111_);
  and (_20175_, _20174_, _20172_);
  and (_20176_, _20110_, word_in[28]);
  or (_36750_, _20176_, _20175_);
  and (_20177_, _20114_, word_in[5]);
  not (_20178_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_20179_, _20114_, _20178_);
  nor (_20180_, _20179_, _20177_);
  nor (_20181_, _20180_, _20113_);
  and (_20182_, _20113_, _19472_);
  nor (_20183_, _20182_, _20181_);
  nor (_20184_, _20183_, _20112_);
  and (_20185_, _20112_, _19171_);
  or (_20186_, _20185_, _20184_);
  and (_20187_, _20186_, _20111_);
  and (_20188_, _20110_, word_in[29]);
  or (_36751_, _20188_, _20187_);
  and (_20189_, _20114_, word_in[6]);
  not (_20190_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_20191_, _20114_, _20190_);
  nor (_20192_, _20191_, _20189_);
  nor (_20193_, _20192_, _20113_);
  and (_20194_, _20113_, _19485_);
  nor (_20195_, _20194_, _20193_);
  nor (_20196_, _20195_, _20112_);
  and (_20197_, _20112_, _19184_);
  or (_20198_, _20197_, _20196_);
  and (_20199_, _20198_, _20111_);
  and (_20200_, _20110_, word_in[30]);
  or (_36752_, _20200_, _20199_);
  nor (_20201_, _20114_, _18489_);
  and (_20202_, _20114_, word_in[7]);
  or (_20203_, _20202_, _20201_);
  or (_20204_, _20203_, _20113_);
  or (_20205_, _20132_, _18791_);
  and (_20206_, _20205_, _20204_);
  or (_20207_, _20206_, _20112_);
  or (_20208_, _20136_, _18795_);
  and (_20209_, _20208_, _20111_);
  and (_20210_, _20209_, _20207_);
  and (_20211_, _20110_, word_in[31]);
  or (_36753_, _20211_, _20210_);
  and (_20212_, _18975_, _18695_);
  and (_20213_, _20212_, _18426_);
  and (_20214_, _18981_, _18778_);
  and (_20215_, _18780_, _18926_);
  and (_20216_, _18785_, _18769_);
  and (_20217_, _20216_, _19096_);
  not (_20218_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_20219_, _20216_, _20218_);
  or (_20220_, _20219_, _20217_);
  or (_20221_, _20220_, _20215_);
  not (_20222_, _20215_);
  or (_20223_, _20222_, word_in[8]);
  and (_20224_, _20223_, _20221_);
  or (_20225_, _20224_, _20214_);
  not (_20226_, _20214_);
  or (_20227_, _20226_, _19104_);
  and (_20228_, _20227_, _20225_);
  or (_20229_, _20228_, _20213_);
  not (_20230_, _20213_);
  or (_20231_, _20230_, word_in[24]);
  and (_36754_, _20231_, _20229_);
  not (_20232_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_20233_, _20216_, _20232_);
  and (_20234_, _20216_, _19112_);
  nor (_20235_, _20234_, _20233_);
  nor (_20236_, _20235_, _20215_);
  and (_20237_, _20215_, word_in[9]);
  nor (_20238_, _20237_, _20236_);
  nor (_20239_, _20238_, _20214_);
  and (_20240_, _20214_, _19119_);
  or (_20241_, _20240_, _20239_);
  and (_20242_, _20241_, _20230_);
  and (_20243_, _20213_, word_in[25]);
  or (_36755_, _20243_, _20242_);
  and (_20244_, _20216_, _19125_);
  not (_20245_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_20246_, _20216_, _20245_);
  nor (_20247_, _20246_, _20244_);
  nor (_20248_, _20247_, _20215_);
  and (_20249_, _20215_, word_in[10]);
  nor (_20250_, _20249_, _20248_);
  nor (_20251_, _20250_, _20214_);
  and (_20252_, _20214_, _19132_);
  or (_20253_, _20252_, _20251_);
  and (_20254_, _20253_, _20230_);
  and (_20255_, _20213_, word_in[26]);
  or (_36756_, _20255_, _20254_);
  and (_20256_, _20216_, word_in[3]);
  not (_20257_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_20258_, _20216_, _20257_);
  nor (_20259_, _20258_, _20256_);
  nor (_20260_, _20259_, _20215_);
  and (_20261_, _20215_, word_in[11]);
  nor (_20262_, _20261_, _20260_);
  nor (_20263_, _20262_, _20214_);
  and (_20264_, _20214_, _19145_);
  or (_20265_, _20264_, _20263_);
  and (_20266_, _20265_, _20230_);
  and (_20267_, _20213_, word_in[27]);
  or (_36757_, _20267_, _20266_);
  and (_20268_, _20216_, word_in[4]);
  not (_20269_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_20270_, _20216_, _20269_);
  nor (_20271_, _20270_, _20268_);
  nor (_20272_, _20271_, _20215_);
  and (_20273_, _20215_, word_in[12]);
  nor (_20274_, _20273_, _20272_);
  nor (_20275_, _20274_, _20214_);
  and (_20276_, _20214_, _19158_);
  or (_20277_, _20276_, _20275_);
  and (_20278_, _20277_, _20230_);
  and (_20279_, _20213_, word_in[28]);
  or (_36758_, _20279_, _20278_);
  and (_20280_, _20216_, word_in[5]);
  not (_20281_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_20282_, _20216_, _20281_);
  nor (_20283_, _20282_, _20280_);
  nor (_20284_, _20283_, _20215_);
  and (_20285_, _20215_, word_in[13]);
  nor (_20286_, _20285_, _20284_);
  nor (_20287_, _20286_, _20214_);
  and (_20288_, _20214_, _19171_);
  or (_20289_, _20288_, _20287_);
  and (_20290_, _20289_, _20230_);
  and (_20291_, _20213_, word_in[29]);
  or (_36759_, _20291_, _20290_);
  not (_20292_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_20293_, _20216_, _20292_);
  and (_20294_, _20216_, _19177_);
  or (_20295_, _20294_, _20293_);
  or (_20296_, _20295_, _20215_);
  or (_20297_, _20222_, word_in[14]);
  and (_20298_, _20297_, _20296_);
  or (_20299_, _20298_, _20214_);
  or (_20300_, _20226_, _19184_);
  and (_20301_, _20300_, _20299_);
  or (_20302_, _20301_, _20213_);
  or (_20303_, _20230_, word_in[30]);
  and (_36760_, _20303_, _20302_);
  and (_20304_, _20216_, word_in[7]);
  nor (_20305_, _20216_, _18593_);
  nor (_20306_, _20305_, _20304_);
  nor (_20307_, _20306_, _20215_);
  and (_20308_, _20215_, word_in[15]);
  nor (_20309_, _20308_, _20307_);
  nor (_20310_, _20309_, _20214_);
  and (_20311_, _20214_, _18795_);
  or (_20312_, _20311_, _20310_);
  and (_20313_, _20312_, _20230_);
  and (_20314_, _20213_, word_in[31]);
  or (_36761_, _20314_, _20313_);
  and (_20315_, _20212_, _18437_);
  and (_20316_, _19090_, _18778_);
  and (_20317_, _18782_, _18414_);
  not (_20318_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_20319_, _18785_, _18966_);
  nor (_20320_, _20319_, _20318_);
  and (_20321_, _19096_, _18966_);
  or (_20322_, _20321_, _20320_);
  or (_20323_, _20322_, _20317_);
  not (_20324_, _20317_);
  or (_20325_, _20324_, _19407_);
  and (_20326_, _20325_, _20323_);
  or (_20327_, _20326_, _20316_);
  not (_20328_, _20316_);
  or (_20329_, _20328_, _19104_);
  and (_20330_, _20329_, _20327_);
  or (_20331_, _20330_, _20315_);
  not (_20332_, _20315_);
  or (_20333_, _20332_, _19414_);
  and (_36762_, _20333_, _20331_);
  not (_20334_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_20335_, _20319_, _20334_);
  and (_20336_, _19112_, _18966_);
  nor (_20337_, _20336_, _20335_);
  nor (_20338_, _20337_, _20317_);
  and (_20339_, _20317_, _19001_);
  or (_20340_, _20339_, _20338_);
  or (_20341_, _20340_, _20316_);
  or (_20342_, _20328_, _19119_);
  and (_20343_, _20342_, _20332_);
  and (_20344_, _20343_, _20341_);
  and (_20345_, _20315_, _19426_);
  or (_36763_, _20345_, _20344_);
  not (_20346_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_20347_, _20319_, _20346_);
  and (_20348_, _19125_, _18966_);
  or (_20349_, _20348_, _20347_);
  or (_20350_, _20349_, _20317_);
  or (_20351_, _20324_, _19432_);
  and (_20352_, _20351_, _20350_);
  or (_20353_, _20352_, _20316_);
  or (_20354_, _20328_, _19132_);
  and (_20355_, _20354_, _20353_);
  or (_20356_, _20355_, _20315_);
  or (_20357_, _20332_, _19439_);
  and (_36764_, _20357_, _20356_);
  or (_20358_, _20324_, _19445_);
  not (_20359_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_20360_, _20319_, _20359_);
  and (_20361_, _20319_, word_in[3]);
  or (_20362_, _20361_, _20360_);
  or (_20363_, _20362_, _20317_);
  and (_20364_, _20363_, _20358_);
  or (_20365_, _20364_, _20316_);
  or (_20366_, _20328_, _19145_);
  and (_20367_, _20366_, _20365_);
  or (_20368_, _20367_, _20315_);
  or (_20369_, _20332_, _19452_);
  and (_36765_, _20369_, _20368_);
  or (_20370_, _20324_, _19454_);
  and (_20371_, _20319_, word_in[4]);
  not (_20372_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_20373_, _20319_, _20372_);
  or (_20374_, _20373_, _20371_);
  or (_20375_, _20374_, _20317_);
  and (_20376_, _20375_, _20370_);
  or (_20377_, _20376_, _20316_);
  or (_20378_, _20328_, _19158_);
  and (_20379_, _20378_, _20332_);
  and (_20380_, _20379_, _20377_);
  and (_20381_, _20315_, _19038_);
  or (_36766_, _20381_, _20380_);
  not (_20382_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_20383_, _20319_, _20382_);
  and (_20384_, _20319_, _19163_);
  or (_20385_, _20384_, _20383_);
  or (_20386_, _20385_, _20317_);
  or (_20387_, _20324_, _19472_);
  and (_20388_, _20387_, _20386_);
  or (_20389_, _20388_, _20316_);
  or (_20390_, _20328_, _19171_);
  and (_20391_, _20390_, _20332_);
  and (_20392_, _20391_, _20389_);
  and (_20393_, _20315_, _19479_);
  or (_36767_, _20393_, _20392_);
  and (_20394_, _20317_, _19485_);
  not (_20395_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  or (_20396_, _20319_, _20395_);
  nand (_20397_, _20319_, _19177_);
  and (_20398_, _20397_, _20396_);
  nor (_20399_, _20398_, _20317_);
  nor (_20400_, _20399_, _20394_);
  nor (_20401_, _20400_, _20316_);
  and (_20402_, _20316_, _19184_);
  or (_20403_, _20402_, _20401_);
  and (_20404_, _20403_, _20332_);
  and (_20405_, _20315_, _19492_);
  or (_36768_, _20405_, _20404_);
  nor (_20406_, _20319_, _18478_);
  and (_20407_, _20319_, _19189_);
  or (_20408_, _20407_, _20406_);
  or (_20409_, _20408_, _20317_);
  or (_20410_, _20324_, _18791_);
  and (_20411_, _20410_, _20409_);
  or (_20412_, _20411_, _20316_);
  or (_20413_, _20328_, _18795_);
  and (_20414_, _20413_, _20332_);
  and (_20415_, _20414_, _20412_);
  and (_20416_, _20315_, _18768_);
  or (_36769_, _20416_, _20415_);
  and (_20417_, _20212_, _18404_);
  and (_20418_, _19205_, _18778_);
  and (_20419_, _18782_, _18426_);
  not (_20420_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_20421_, _18785_, _18804_);
  nor (_20422_, _20421_, _20420_);
  and (_20423_, _20421_, _19096_);
  or (_20424_, _20423_, _20422_);
  or (_20425_, _20424_, _20419_);
  not (_20426_, _20419_);
  or (_20427_, _20426_, _19407_);
  and (_20428_, _20427_, _20425_);
  or (_20429_, _20428_, _20418_);
  not (_20430_, _20418_);
  or (_20431_, _20430_, _19104_);
  and (_20432_, _20431_, _20429_);
  or (_20433_, _20432_, _20417_);
  not (_20434_, _20417_);
  or (_20435_, _20434_, word_in[24]);
  and (_36770_, _20435_, _20433_);
  or (_20436_, _20426_, _19001_);
  and (_20437_, _20421_, word_in[1]);
  not (_20438_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_20439_, _20421_, _20438_);
  or (_20440_, _20439_, _20437_);
  or (_20441_, _20440_, _20419_);
  and (_20442_, _20441_, _20436_);
  or (_20443_, _20442_, _20418_);
  or (_20444_, _20430_, _19119_);
  and (_20445_, _20444_, _20443_);
  or (_20446_, _20445_, _20417_);
  or (_20447_, _20434_, word_in[25]);
  and (_36771_, _20447_, _20446_);
  or (_20448_, _20426_, _19432_);
  and (_20449_, _20421_, word_in[2]);
  not (_20450_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_20451_, _20421_, _20450_);
  or (_20452_, _20451_, _20449_);
  or (_20453_, _20452_, _20419_);
  and (_20454_, _20453_, _20448_);
  or (_20455_, _20454_, _20418_);
  or (_20456_, _20430_, _19132_);
  and (_20457_, _20456_, _20434_);
  and (_20458_, _20457_, _20455_);
  and (_20459_, _20417_, _19439_);
  or (_36772_, _20459_, _20458_);
  and (_20460_, _20418_, _19145_);
  not (_20461_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_20462_, _20421_, _20461_);
  and (_20463_, _20421_, word_in[3]);
  nor (_20464_, _20463_, _20462_);
  nor (_20465_, _20464_, _20419_);
  and (_20466_, _20419_, _19445_);
  nor (_20467_, _20466_, _20465_);
  nor (_20468_, _20467_, _20418_);
  or (_20469_, _20468_, _20460_);
  and (_20470_, _20469_, _20434_);
  and (_20471_, _20417_, word_in[27]);
  or (_36773_, _20471_, _20470_);
  or (_20472_, _20430_, _19158_);
  not (_20473_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_20474_, _20421_, _20473_);
  and (_20475_, _20421_, _19151_);
  or (_20476_, _20475_, _20474_);
  or (_20477_, _20476_, _20419_);
  or (_20478_, _20426_, _19454_);
  and (_20479_, _20478_, _20477_);
  or (_20480_, _20479_, _20418_);
  and (_20481_, _20480_, _20472_);
  or (_20482_, _20481_, _20417_);
  or (_20483_, _20434_, word_in[28]);
  and (_36774_, _20483_, _20482_);
  or (_20484_, _20426_, _19472_);
  and (_20485_, _20421_, word_in[5]);
  not (_20486_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_20487_, _20421_, _20486_);
  or (_20488_, _20487_, _20485_);
  or (_20489_, _20488_, _20419_);
  and (_20490_, _20489_, _20484_);
  or (_20491_, _20490_, _20418_);
  or (_20492_, _20430_, _19171_);
  and (_20493_, _20492_, _20434_);
  and (_20494_, _20493_, _20491_);
  and (_20495_, _20417_, _19479_);
  or (_36775_, _20495_, _20494_);
  or (_20496_, _20426_, _19485_);
  and (_20497_, _20421_, word_in[6]);
  not (_20498_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_20499_, _20421_, _20498_);
  or (_20500_, _20499_, _20497_);
  or (_20501_, _20500_, _20419_);
  and (_20502_, _20501_, _20496_);
  or (_20503_, _20502_, _20418_);
  or (_20504_, _20430_, _19184_);
  and (_20505_, _20504_, _20503_);
  or (_20506_, _20505_, _20417_);
  or (_20507_, _20434_, word_in[30]);
  and (_36776_, _20507_, _20506_);
  and (_20508_, _20421_, word_in[7]);
  nor (_20509_, _20421_, _18598_);
  nor (_20510_, _20509_, _20508_);
  nor (_20511_, _20510_, _20419_);
  and (_20512_, _20419_, _18791_);
  nor (_20513_, _20512_, _20511_);
  nor (_20514_, _20513_, _20418_);
  and (_20515_, _20418_, _18795_);
  or (_20516_, _20515_, _20514_);
  and (_20517_, _20516_, _20434_);
  and (_20518_, _20417_, word_in[31]);
  or (_36777_, _20518_, _20517_);
  and (_20519_, _19414_, _18770_);
  and (_20520_, _18786_, word_in[0]);
  not (_20521_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_20522_, _18786_, _20521_);
  nor (_20523_, _20522_, _20520_);
  nor (_20524_, _20523_, _18783_);
  and (_20525_, _19407_, _18783_);
  nor (_20526_, _20525_, _20524_);
  nor (_20527_, _20526_, _18779_);
  and (_20528_, _19104_, _18779_);
  or (_20529_, _20528_, _20527_);
  and (_20530_, _20529_, _18772_);
  or (_36778_, _20530_, _20519_);
  not (_20531_, _18783_);
  or (_20532_, _19001_, _20531_);
  and (_20533_, _18786_, word_in[1]);
  not (_20534_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_20535_, _18786_, _20534_);
  or (_20536_, _20535_, _20533_);
  or (_20537_, _20536_, _18783_);
  and (_20538_, _20537_, _20532_);
  or (_20539_, _20538_, _18779_);
  not (_20540_, _18779_);
  or (_20541_, _19119_, _20540_);
  and (_20542_, _20541_, _18772_);
  and (_20543_, _20542_, _20539_);
  and (_20544_, _19426_, _18770_);
  or (_36779_, _20544_, _20543_);
  and (_20545_, _19439_, _18770_);
  and (_20546_, _18786_, word_in[2]);
  not (_20547_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_20548_, _18786_, _20547_);
  nor (_20549_, _20548_, _20546_);
  nor (_20550_, _20549_, _18783_);
  and (_20551_, _19432_, _18783_);
  nor (_20552_, _20551_, _20550_);
  nor (_20553_, _20552_, _18779_);
  and (_20554_, _19132_, _18779_);
  or (_20555_, _20554_, _20553_);
  and (_20556_, _20555_, _18772_);
  or (_36780_, _20556_, _20545_);
  or (_20557_, _19445_, _20531_);
  and (_20558_, _18786_, word_in[3]);
  not (_20559_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_20560_, _18786_, _20559_);
  or (_20561_, _20560_, _20558_);
  or (_20562_, _20561_, _18783_);
  and (_20563_, _20562_, _20557_);
  or (_20564_, _20563_, _18779_);
  or (_20565_, _19145_, _20540_);
  and (_20566_, _20565_, _20564_);
  or (_20567_, _20566_, _18770_);
  or (_20568_, _18772_, word_in[27]);
  and (_36781_, _20568_, _20567_);
  and (_20569_, _19038_, _18770_);
  and (_20570_, _18786_, word_in[4]);
  not (_20571_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_20572_, _18786_, _20571_);
  nor (_20573_, _20572_, _20570_);
  nor (_20574_, _20573_, _18783_);
  and (_20575_, _19454_, _18783_);
  nor (_20576_, _20575_, _20574_);
  nor (_20577_, _20576_, _18779_);
  and (_20578_, _19158_, _18779_);
  or (_20579_, _20578_, _20577_);
  and (_20580_, _20579_, _18772_);
  or (_36782_, _20580_, _20569_);
  and (_20581_, _18770_, word_in[29]);
  or (_20582_, _19472_, _20531_);
  and (_20583_, _18786_, word_in[5]);
  not (_20584_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_20585_, _18786_, _20584_);
  or (_20586_, _20585_, _20583_);
  or (_20587_, _20586_, _18783_);
  and (_20588_, _20587_, _20582_);
  or (_20589_, _20588_, _18779_);
  or (_20590_, _19171_, _20540_);
  and (_20591_, _20590_, _18772_);
  and (_20592_, _20591_, _20589_);
  or (_36783_, _20592_, _20581_);
  not (_20593_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_20594_, _18786_, _20593_);
  and (_20595_, _19177_, _18786_);
  or (_20596_, _20595_, _20594_);
  or (_20597_, _20596_, _18783_);
  or (_20598_, _19485_, _20531_);
  and (_20599_, _20598_, _20597_);
  or (_20600_, _20599_, _18779_);
  or (_20601_, _19184_, _20540_);
  and (_20602_, _20601_, _18772_);
  and (_20603_, _20602_, _20600_);
  and (_20604_, _18770_, word_in[30]);
  or (_36784_, _20604_, _20603_);
  and (_20605_, _18441_, word_in[0]);
  not (_20606_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand (_20607_, _18400_, _20606_);
  or (_20608_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_20609_, _20608_, _20607_);
  and (_20610_, _20609_, _18447_);
  nor (_20611_, _20610_, _18385_);
  not (_20612_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_20613_, _18400_, _20612_);
  or (_20614_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_20615_, _20614_, _20613_);
  and (_20616_, _20615_, _18456_);
  nand (_20617_, _18400_, _19705_);
  or (_20618_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_20619_, _20618_, _20617_);
  and (_20620_, _20619_, _18450_);
  not (_20621_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_20622_, _18400_, _20621_);
  or (_20623_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_20624_, _20623_, _20622_);
  and (_20625_, _20624_, _18466_);
  or (_20626_, _20625_, _20620_);
  nor (_20627_, _20626_, _20616_);
  and (_20628_, _20627_, _20611_);
  nand (_20629_, _18400_, _19913_);
  or (_20630_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_20631_, _20630_, _20629_);
  and (_20632_, _20631_, _18447_);
  nor (_20633_, _20632_, _18471_);
  nand (_20634_, _18400_, _20318_);
  or (_20635_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_20636_, _20635_, _20634_);
  and (_20637_, _20636_, _18456_);
  nand (_20638_, _18400_, _20521_);
  or (_20639_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_20640_, _20639_, _20638_);
  and (_20641_, _20640_, _18450_);
  nand (_20642_, _18400_, _20116_);
  or (_20643_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_20644_, _20643_, _20642_);
  and (_20645_, _20644_, _18466_);
  or (_20646_, _20645_, _20641_);
  nor (_20647_, _20646_, _20637_);
  and (_20648_, _20647_, _20633_);
  or (_20649_, _20648_, _20628_);
  nor (_20650_, _20649_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _20650_, _20605_);
  and (_20651_, _18441_, word_in[1]);
  not (_20652_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nand (_20653_, _18400_, _20652_);
  or (_20654_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_20655_, _20654_, _20653_);
  and (_20656_, _20655_, _18447_);
  nor (_20657_, _20656_, _18385_);
  not (_20658_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nand (_20659_, _18400_, _20658_);
  or (_20660_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_20661_, _20660_, _20659_);
  and (_20662_, _20661_, _18456_);
  nand (_20663_, _18400_, _19721_);
  or (_20664_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_20665_, _20664_, _20663_);
  and (_20666_, _20665_, _18450_);
  not (_20667_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand (_20668_, _18400_, _20667_);
  or (_20669_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_20670_, _20669_, _20668_);
  and (_20671_, _20670_, _18466_);
  or (_20672_, _20671_, _20666_);
  nor (_20673_, _20672_, _20662_);
  and (_20674_, _20673_, _20657_);
  nand (_20675_, _18400_, _19925_);
  or (_20676_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_20677_, _20676_, _20675_);
  and (_20678_, _20677_, _18447_);
  nor (_20679_, _20678_, _18471_);
  nand (_20680_, _18400_, _20334_);
  or (_20681_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_20682_, _20681_, _20680_);
  and (_20683_, _20682_, _18456_);
  nand (_20684_, _18400_, _20534_);
  or (_20685_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_20686_, _20685_, _20684_);
  and (_20687_, _20686_, _18450_);
  nand (_20688_, _18400_, _20127_);
  or (_20689_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_20690_, _20689_, _20688_);
  and (_20691_, _20690_, _18466_);
  or (_20692_, _20691_, _20687_);
  nor (_20693_, _20692_, _20683_);
  and (_20694_, _20693_, _20679_);
  or (_20695_, _20694_, _20674_);
  nor (_20696_, _20695_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _20696_, _20651_);
  and (_20697_, _18441_, word_in[2]);
  not (_20698_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_20699_, _18400_, _20698_);
  or (_20700_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_20701_, _20700_, _20699_);
  and (_20702_, _20701_, _18447_);
  nor (_20703_, _20702_, _18385_);
  not (_20704_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_20705_, _18400_, _20704_);
  or (_20706_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_20707_, _20706_, _20705_);
  and (_20708_, _20707_, _18456_);
  nand (_20709_, _18400_, _19735_);
  or (_20710_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_20711_, _20710_, _20709_);
  and (_20712_, _20711_, _18450_);
  not (_20713_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand (_20714_, _18400_, _20713_);
  or (_20715_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_20716_, _20715_, _20714_);
  and (_20717_, _20716_, _18466_);
  or (_20718_, _20717_, _20712_);
  nor (_20719_, _20718_, _20708_);
  and (_20720_, _20719_, _20703_);
  nand (_20721_, _18400_, _19937_);
  or (_20722_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_20723_, _20722_, _20721_);
  and (_20724_, _20723_, _18447_);
  nor (_20725_, _20724_, _18471_);
  nand (_20726_, _18400_, _20547_);
  or (_20727_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_20728_, _20727_, _20726_);
  and (_20729_, _20728_, _18450_);
  nand (_20730_, _18400_, _20346_);
  or (_20731_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_20732_, _20731_, _20730_);
  and (_20733_, _20732_, _18456_);
  or (_20734_, _20733_, _20729_);
  nand (_20735_, _18400_, _20142_);
  or (_20736_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_20737_, _20736_, _20735_);
  and (_20738_, _20737_, _18466_);
  nor (_20739_, _20738_, _20734_);
  and (_20740_, _20739_, _20725_);
  or (_20741_, _20740_, _20720_);
  nor (_20742_, _20741_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _20742_, _20697_);
  and (_20743_, _18441_, word_in[3]);
  not (_20744_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nand (_20745_, _18400_, _20744_);
  or (_20746_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_20747_, _20746_, _20745_);
  and (_20748_, _20747_, _18447_);
  nor (_20749_, _20748_, _18385_);
  not (_20750_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nand (_20751_, _18400_, _20750_);
  or (_20752_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_20753_, _20752_, _20751_);
  and (_20754_, _20753_, _18456_);
  nand (_20755_, _18400_, _19745_);
  or (_20756_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_20757_, _20756_, _20755_);
  and (_20758_, _20757_, _18450_);
  not (_20759_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nand (_20760_, _18400_, _20759_);
  or (_20761_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_20762_, _20761_, _20760_);
  and (_20763_, _20762_, _18466_);
  or (_20764_, _20763_, _20758_);
  nor (_20765_, _20764_, _20754_);
  and (_20766_, _20765_, _20749_);
  nand (_20767_, _18400_, _19951_);
  or (_20768_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_20769_, _20768_, _20767_);
  and (_20770_, _20769_, _18447_);
  nor (_20771_, _20770_, _18471_);
  nand (_20772_, _18400_, _20359_);
  or (_20773_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_20774_, _20773_, _20772_);
  and (_20775_, _20774_, _18456_);
  nand (_20776_, _18400_, _20559_);
  or (_20777_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_20778_, _20777_, _20776_);
  and (_20779_, _20778_, _18450_);
  nand (_20780_, _18400_, _20154_);
  or (_20781_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_20782_, _20781_, _20780_);
  and (_20783_, _20782_, _18466_);
  or (_20784_, _20783_, _20779_);
  nor (_20785_, _20784_, _20775_);
  and (_20786_, _20785_, _20771_);
  or (_20787_, _20786_, _20766_);
  nor (_20788_, _20787_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _20788_, _20743_);
  and (_20789_, _18441_, word_in[4]);
  not (_20790_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand (_20791_, _18400_, _20790_);
  or (_20792_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_20793_, _20792_, _20791_);
  and (_20794_, _20793_, _18447_);
  nor (_20795_, _20794_, _18385_);
  not (_20796_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nand (_20797_, _18400_, _20796_);
  or (_20798_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_20799_, _20798_, _20797_);
  and (_20800_, _20799_, _18456_);
  nand (_20801_, _18400_, _19759_);
  or (_20802_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_20803_, _20802_, _20801_);
  and (_20804_, _20803_, _18450_);
  not (_20805_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nand (_20806_, _18400_, _20805_);
  or (_20807_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_20808_, _20807_, _20806_);
  and (_20809_, _20808_, _18466_);
  or (_20810_, _20809_, _20804_);
  nor (_20811_, _20810_, _20800_);
  and (_20812_, _20811_, _20795_);
  nand (_20813_, _18400_, _19963_);
  or (_20814_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_20815_, _20814_, _20813_);
  and (_20816_, _20815_, _18447_);
  nor (_20817_, _20816_, _18471_);
  nand (_20818_, _18400_, _20372_);
  or (_20819_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_20820_, _20819_, _20818_);
  and (_20821_, _20820_, _18456_);
  nand (_20822_, _18400_, _20571_);
  or (_20823_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_20824_, _20823_, _20822_);
  and (_20825_, _20824_, _18450_);
  nand (_20826_, _18400_, _20165_);
  or (_20827_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_20828_, _20827_, _20826_);
  and (_20829_, _20828_, _18466_);
  or (_20830_, _20829_, _20825_);
  nor (_20831_, _20830_, _20821_);
  and (_20832_, _20831_, _20817_);
  or (_20833_, _20832_, _20812_);
  nor (_20834_, _20833_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _20834_, _20789_);
  and (_20835_, _18441_, word_in[5]);
  not (_20836_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nand (_20837_, _18400_, _20836_);
  or (_20838_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_20839_, _20838_, _20837_);
  and (_20840_, _20839_, _18447_);
  nor (_20841_, _20840_, _18385_);
  not (_20842_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nand (_20843_, _18400_, _20842_);
  or (_20844_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_20845_, _20844_, _20843_);
  and (_20846_, _20845_, _18456_);
  nand (_20847_, _18400_, _19770_);
  or (_20848_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_20849_, _20848_, _20847_);
  and (_20850_, _20849_, _18450_);
  not (_20851_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand (_20852_, _18400_, _20851_);
  or (_20853_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_20854_, _20853_, _20852_);
  and (_20855_, _20854_, _18466_);
  or (_20856_, _20855_, _20850_);
  nor (_20857_, _20856_, _20846_);
  and (_20858_, _20857_, _20841_);
  nand (_20859_, _18400_, _19975_);
  or (_20860_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_20861_, _20860_, _20859_);
  and (_20862_, _20861_, _18447_);
  nor (_20863_, _20862_, _18471_);
  nand (_20864_, _18400_, _20382_);
  or (_20865_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_20866_, _20865_, _20864_);
  and (_20867_, _20866_, _18456_);
  nand (_20868_, _18400_, _20584_);
  or (_20869_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_20870_, _20869_, _20868_);
  and (_20871_, _20870_, _18450_);
  nand (_20872_, _18400_, _20178_);
  or (_20873_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_20874_, _20873_, _20872_);
  and (_20875_, _20874_, _18466_);
  or (_20876_, _20875_, _20871_);
  nor (_20877_, _20876_, _20867_);
  and (_20878_, _20877_, _20863_);
  or (_20879_, _20878_, _20858_);
  nor (_20880_, _20879_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _20880_, _20835_);
  and (_20881_, _18441_, word_in[6]);
  not (_20882_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nand (_20883_, _18400_, _20882_);
  or (_20884_, _18400_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_20885_, _20884_, _20883_);
  and (_20886_, _20885_, _18447_);
  nor (_20887_, _20886_, _18385_);
  not (_20888_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nand (_20889_, _18400_, _20888_);
  or (_20890_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_20891_, _20890_, _20889_);
  and (_20892_, _20891_, _18456_);
  nand (_20893_, _18400_, _19782_);
  or (_20894_, _18400_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_20895_, _20894_, _20893_);
  and (_20896_, _20895_, _18450_);
  not (_20897_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nand (_20898_, _18400_, _20897_);
  or (_20899_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_20900_, _20899_, _20898_);
  and (_20901_, _20900_, _18466_);
  or (_20902_, _20901_, _20896_);
  nor (_20903_, _20902_, _20892_);
  and (_20904_, _20903_, _20887_);
  nand (_20905_, _18400_, _19988_);
  or (_20906_, _18400_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_20907_, _20906_, _20905_);
  and (_20908_, _20907_, _18447_);
  nor (_20909_, _20908_, _18471_);
  nand (_20910_, _18400_, _20593_);
  or (_20911_, _18400_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_20912_, _20911_, _20910_);
  and (_20913_, _20912_, _18450_);
  nand (_20914_, _18400_, _20395_);
  or (_20915_, _18400_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_20916_, _20915_, _20914_);
  and (_20917_, _20916_, _18456_);
  or (_20918_, _20917_, _20913_);
  nand (_20919_, _18400_, _20190_);
  or (_20920_, _18400_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_20921_, _20920_, _20919_);
  and (_20922_, _20921_, _18466_);
  nor (_20923_, _20922_, _20918_);
  and (_20924_, _20923_, _20909_);
  or (_20925_, _20924_, _20904_);
  nor (_20926_, _20925_, _18441_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _20926_, _20881_);
  and (_20927_, _18553_, word_in[8]);
  nand (_20928_, _18400_, _18987_);
  or (_20929_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_20930_, _20929_, _20928_);
  and (_20931_, _20930_, _18555_);
  and (_20932_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_20933_, _18400_, _20621_);
  or (_20934_, _20933_, _20932_);
  and (_20935_, _20934_, _18561_);
  nor (_20936_, _20935_, _20931_);
  nor (_20937_, _20936_, _18500_);
  and (_20938_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_20939_, _18400_, _20612_);
  or (_20940_, _20939_, _20938_);
  and (_20941_, _20940_, _18555_);
  nand (_20942_, _18400_, _19604_);
  or (_20943_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_20944_, _20943_, _20942_);
  and (_20945_, _20944_, _18561_);
  or (_20946_, _20945_, _20941_);
  and (_20947_, _20946_, _18500_);
  or (_20948_, _20947_, _20937_);
  and (_20949_, _20948_, _18504_);
  nand (_20950_, _18400_, _19807_);
  or (_20951_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_20952_, _20951_, _20950_);
  and (_20953_, _20952_, _18555_);
  nand (_20954_, _18400_, _20016_);
  or (_20955_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_20956_, _20955_, _20954_);
  and (_20957_, _20956_, _18561_);
  nor (_20958_, _20957_, _20953_);
  nor (_20959_, _20958_, _18500_);
  nand (_20960_, _18400_, _20218_);
  or (_20961_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_20962_, _20961_, _20960_);
  and (_20963_, _20962_, _18555_);
  nand (_20964_, _18400_, _20420_);
  or (_20965_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_20966_, _20965_, _20964_);
  and (_20967_, _20966_, _18561_);
  or (_20968_, _20967_, _20963_);
  and (_20969_, _20968_, _18500_);
  nor (_20970_, _20969_, _20959_);
  nor (_20971_, _20970_, _18504_);
  nor (_20972_, _20971_, _20949_);
  nor (_20973_, _20972_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _20973_, _20927_);
  and (_20974_, _18553_, word_in[9]);
  nand (_20975_, _18400_, _19003_);
  or (_20976_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_20977_, _20976_, _20975_);
  and (_20978_, _20977_, _18555_);
  and (_20979_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_20980_, _18400_, _20667_);
  or (_20981_, _20980_, _20979_);
  and (_20982_, _20981_, _18561_);
  nor (_20983_, _20982_, _20978_);
  nor (_20984_, _20983_, _18500_);
  and (_20985_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_20986_, _18400_, _20658_);
  or (_20987_, _20986_, _20985_);
  and (_20988_, _20987_, _18555_);
  nand (_20989_, _18400_, _19618_);
  or (_20990_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_20991_, _20990_, _20989_);
  and (_20992_, _20991_, _18561_);
  or (_20993_, _20992_, _20988_);
  and (_20994_, _20993_, _18500_);
  or (_20995_, _20994_, _20984_);
  and (_20996_, _20995_, _18504_);
  nand (_20997_, _18400_, _19825_);
  or (_20998_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_20999_, _20998_, _20997_);
  and (_21000_, _20999_, _18555_);
  nand (_21001_, _18400_, _20028_);
  or (_21002_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_21003_, _21002_, _21001_);
  and (_21004_, _21003_, _18561_);
  nor (_21005_, _21004_, _21000_);
  nor (_21006_, _21005_, _18500_);
  nand (_21007_, _18400_, _20232_);
  or (_21008_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_21009_, _21008_, _21007_);
  and (_21010_, _21009_, _18555_);
  nand (_21011_, _18400_, _20438_);
  or (_21012_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_21013_, _21012_, _21011_);
  and (_21014_, _21013_, _18561_);
  or (_21015_, _21014_, _21010_);
  and (_21016_, _21015_, _18500_);
  nor (_21017_, _21016_, _21006_);
  nor (_21018_, _21017_, _18504_);
  nor (_21019_, _21018_, _20996_);
  nor (_21020_, _21019_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _21020_, _20974_);
  and (_21021_, _18553_, word_in[10]);
  nand (_21022_, _18400_, _19016_);
  or (_21023_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_21024_, _21023_, _21022_);
  and (_21025_, _21024_, _18555_);
  and (_21026_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_21027_, _18400_, _20713_);
  or (_21028_, _21027_, _21026_);
  and (_21029_, _21028_, _18561_);
  nor (_21030_, _21029_, _21025_);
  nor (_21031_, _21030_, _18500_);
  and (_21032_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_21033_, _18400_, _20704_);
  or (_21034_, _21033_, _21032_);
  and (_21035_, _21034_, _18555_);
  nand (_21036_, _18400_, _19632_);
  or (_21037_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_21038_, _21037_, _21036_);
  and (_21039_, _21038_, _18561_);
  or (_21040_, _21039_, _21035_);
  and (_21041_, _21040_, _18500_);
  or (_21042_, _21041_, _21031_);
  and (_21043_, _21042_, _18504_);
  nand (_21044_, _18400_, _19837_);
  or (_21045_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_21046_, _21045_, _21044_);
  and (_21047_, _21046_, _18555_);
  nand (_21048_, _18400_, _20040_);
  or (_21049_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_21050_, _21049_, _21048_);
  and (_21051_, _21050_, _18561_);
  nor (_21052_, _21051_, _21047_);
  nor (_21053_, _21052_, _18500_);
  nand (_21054_, _18400_, _20245_);
  or (_21055_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_21056_, _21055_, _21054_);
  and (_21057_, _21056_, _18555_);
  nand (_21058_, _18400_, _20450_);
  or (_21059_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _18561_);
  or (_21062_, _21061_, _21057_);
  and (_21063_, _21062_, _18500_);
  nor (_21064_, _21063_, _21053_);
  nor (_21065_, _21064_, _18504_);
  nor (_21066_, _21065_, _21043_);
  nor (_21067_, _21066_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _21067_, _21021_);
  and (_21068_, _18553_, word_in[11]);
  nand (_21069_, _18400_, _19027_);
  or (_21070_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_21071_, _21070_, _21069_);
  and (_21072_, _21071_, _18555_);
  and (_21073_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_21074_, _18400_, _20759_);
  or (_21075_, _21074_, _21073_);
  and (_21076_, _21075_, _18561_);
  nor (_21077_, _21076_, _21072_);
  nor (_21078_, _21077_, _18500_);
  and (_21079_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_21080_, _18400_, _20750_);
  or (_21081_, _21080_, _21079_);
  and (_21082_, _21081_, _18555_);
  nand (_21083_, _18400_, _19645_);
  or (_21084_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_21085_, _21084_, _21083_);
  and (_21086_, _21085_, _18561_);
  or (_21087_, _21086_, _21082_);
  and (_21088_, _21087_, _18500_);
  or (_21089_, _21088_, _21078_);
  and (_21090_, _21089_, _18504_);
  nand (_21091_, _18400_, _19849_);
  or (_21092_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_21093_, _21092_, _21091_);
  and (_21094_, _21093_, _18555_);
  nand (_21095_, _18400_, _20052_);
  or (_21096_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_21097_, _21096_, _21095_);
  and (_21098_, _21097_, _18561_);
  nor (_21099_, _21098_, _21094_);
  nor (_21100_, _21099_, _18500_);
  nand (_21101_, _18400_, _20257_);
  or (_21102_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_21103_, _21102_, _21101_);
  and (_21104_, _21103_, _18555_);
  nand (_21105_, _18400_, _20461_);
  or (_21106_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_21107_, _21106_, _21105_);
  and (_21108_, _21107_, _18561_);
  or (_21109_, _21108_, _21104_);
  and (_21110_, _21109_, _18500_);
  nor (_21111_, _21110_, _21100_);
  nor (_21112_, _21111_, _18504_);
  nor (_21113_, _21112_, _21090_);
  nor (_21114_, _21113_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _21114_, _21068_);
  and (_21115_, _18553_, word_in[12]);
  nand (_21116_, _18400_, _19042_);
  or (_21117_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_21118_, _21117_, _21116_);
  and (_21119_, _21118_, _18555_);
  and (_21120_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_21121_, _18400_, _20805_);
  or (_21122_, _21121_, _21120_);
  and (_21123_, _21122_, _18561_);
  nor (_21124_, _21123_, _21119_);
  nor (_21125_, _21124_, _18500_);
  and (_21126_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_21127_, _18400_, _20796_);
  or (_21128_, _21127_, _21126_);
  and (_21129_, _21128_, _18555_);
  nand (_21130_, _18400_, _19657_);
  or (_21131_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_21132_, _21131_, _21130_);
  and (_21133_, _21132_, _18561_);
  or (_21134_, _21133_, _21129_);
  and (_21135_, _21134_, _18500_);
  or (_21136_, _21135_, _21125_);
  and (_21137_, _21136_, _18504_);
  nand (_21138_, _18400_, _19860_);
  or (_21139_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_21140_, _21139_, _21138_);
  and (_21141_, _21140_, _18555_);
  nand (_21142_, _18400_, _20064_);
  or (_21143_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_21144_, _21143_, _21142_);
  and (_21145_, _21144_, _18561_);
  nor (_21146_, _21145_, _21141_);
  nor (_21147_, _21146_, _18500_);
  nand (_21148_, _18400_, _20269_);
  or (_21149_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_21150_, _21149_, _21148_);
  and (_21151_, _21150_, _18555_);
  nand (_21152_, _18400_, _20473_);
  or (_21153_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_21154_, _21153_, _21152_);
  and (_21155_, _21154_, _18561_);
  or (_21156_, _21155_, _21151_);
  and (_21157_, _21156_, _18500_);
  nor (_21158_, _21157_, _21147_);
  nor (_21159_, _21158_, _18504_);
  nor (_21160_, _21159_, _21137_);
  nor (_21161_, _21160_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _21161_, _21115_);
  and (_21162_, _18553_, word_in[13]);
  nand (_21163_, _18400_, _19054_);
  or (_21164_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_21165_, _21164_, _21163_);
  and (_21166_, _21165_, _18555_);
  and (_21167_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_21168_, _18400_, _20851_);
  or (_21169_, _21168_, _21167_);
  and (_21170_, _21169_, _18561_);
  nor (_21171_, _21170_, _21166_);
  nor (_21172_, _21171_, _18500_);
  and (_21173_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_21174_, _18400_, _20842_);
  or (_21175_, _21174_, _21173_);
  and (_21176_, _21175_, _18555_);
  nand (_21177_, _18400_, _19667_);
  or (_21178_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_21179_, _21178_, _21177_);
  and (_21180_, _21179_, _18561_);
  or (_21181_, _21180_, _21176_);
  and (_21182_, _21181_, _18500_);
  or (_21183_, _21182_, _21172_);
  and (_21184_, _21183_, _18504_);
  nand (_21185_, _18400_, _19873_);
  or (_21186_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_21187_, _21186_, _21185_);
  and (_21188_, _21187_, _18555_);
  nand (_21189_, _18400_, _20076_);
  or (_21190_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_21191_, _21190_, _21189_);
  and (_21192_, _21191_, _18561_);
  nor (_21193_, _21192_, _21188_);
  nor (_21194_, _21193_, _18500_);
  nand (_21195_, _18400_, _20281_);
  or (_21196_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_21197_, _21196_, _21195_);
  and (_21198_, _21197_, _18555_);
  nand (_21199_, _18400_, _20486_);
  or (_21200_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_21201_, _21200_, _21199_);
  and (_21202_, _21201_, _18561_);
  or (_21203_, _21202_, _21198_);
  and (_21204_, _21203_, _18500_);
  nor (_21205_, _21204_, _21194_);
  nor (_21206_, _21205_, _18504_);
  nor (_21207_, _21206_, _21184_);
  nor (_21208_, _21207_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _21208_, _21162_);
  and (_21209_, _18553_, word_in[14]);
  nand (_21210_, _18400_, _19065_);
  or (_21211_, _18400_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_21212_, _21211_, _21210_);
  and (_21213_, _21212_, _18555_);
  and (_21214_, _18400_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_21215_, _18400_, _20897_);
  or (_21216_, _21215_, _21214_);
  and (_21217_, _21216_, _18561_);
  nor (_21218_, _21217_, _21213_);
  nor (_21219_, _21218_, _18500_);
  and (_21220_, _18400_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_21221_, _18400_, _20888_);
  or (_21222_, _21221_, _21220_);
  and (_21223_, _21222_, _18555_);
  nand (_21224_, _18400_, _19679_);
  or (_21225_, _18400_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_21226_, _21225_, _21224_);
  and (_21227_, _21226_, _18561_);
  or (_21228_, _21227_, _21223_);
  and (_21229_, _21228_, _18500_);
  or (_21230_, _21229_, _21219_);
  and (_21231_, _21230_, _18504_);
  nand (_21232_, _18400_, _19885_);
  or (_21233_, _18400_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_21234_, _21233_, _21232_);
  and (_21235_, _21234_, _18555_);
  nand (_21236_, _18400_, _20087_);
  or (_21237_, _18400_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_21238_, _21237_, _21236_);
  and (_21239_, _21238_, _18561_);
  nor (_21240_, _21239_, _21235_);
  nor (_21241_, _21240_, _18500_);
  nand (_21242_, _18400_, _20292_);
  or (_21243_, _18400_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_21244_, _21243_, _21242_);
  and (_21245_, _21244_, _18555_);
  nand (_21246_, _18400_, _20498_);
  or (_21247_, _18400_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_21248_, _21247_, _21246_);
  and (_21249_, _21248_, _18561_);
  or (_21250_, _21249_, _21245_);
  and (_21251_, _21250_, _18500_);
  nor (_21252_, _21251_, _21241_);
  nor (_21253_, _21252_, _18504_);
  nor (_21254_, _21253_, _21231_);
  nor (_21255_, _21254_, _18553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _21255_, _21209_);
  and (_21256_, _18672_, word_in[16]);
  and (_21257_, _20636_, _18466_);
  and (_21258_, _20640_, _18456_);
  or (_21259_, _21258_, _21257_);
  and (_21260_, _20631_, _18450_);
  and (_21261_, _20644_, _18447_);
  or (_21262_, _21261_, _21260_);
  or (_21263_, _21262_, _21259_);
  or (_21264_, _21263_, _18613_);
  and (_21265_, _20615_, _18466_);
  and (_21266_, _20619_, _18456_);
  or (_21267_, _21266_, _21265_);
  and (_21268_, _20609_, _18450_);
  and (_21269_, _20624_, _18447_);
  or (_21270_, _21269_, _21268_);
  nor (_21271_, _21270_, _21267_);
  nand (_21272_, _21271_, _18613_);
  and (_21273_, _21272_, _21264_);
  and (_21274_, _21273_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _21274_, _21256_);
  and (_21275_, _18672_, word_in[17]);
  and (_21276_, _20686_, _18456_);
  and (_21277_, _20682_, _18466_);
  or (_21278_, _21277_, _21276_);
  and (_21279_, _20690_, _18447_);
  and (_21280_, _20677_, _18450_);
  or (_21281_, _21280_, _21279_);
  or (_21282_, _21281_, _21278_);
  or (_21283_, _21282_, _18613_);
  and (_21284_, _20665_, _18456_);
  and (_21285_, _20661_, _18466_);
  or (_21286_, _21285_, _21284_);
  and (_21287_, _20670_, _18447_);
  and (_21288_, _20655_, _18450_);
  or (_21289_, _21288_, _21287_);
  nor (_21290_, _21289_, _21286_);
  nand (_21291_, _21290_, _18613_);
  and (_21292_, _21291_, _21283_);
  and (_21293_, _21292_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _21293_, _21275_);
  and (_21294_, _18672_, word_in[18]);
  and (_21295_, _20732_, _18466_);
  and (_21296_, _20728_, _18456_);
  or (_21297_, _21296_, _21295_);
  and (_21298_, _20723_, _18450_);
  and (_21299_, _20737_, _18447_);
  or (_21300_, _21299_, _21298_);
  or (_21301_, _21300_, _21297_);
  or (_21302_, _21301_, _18613_);
  and (_21303_, _20707_, _18466_);
  and (_21304_, _20711_, _18456_);
  or (_21305_, _21304_, _21303_);
  and (_21306_, _20701_, _18450_);
  and (_21307_, _20716_, _18447_);
  or (_21308_, _21307_, _21306_);
  nor (_21309_, _21308_, _21305_);
  nand (_21310_, _21309_, _18613_);
  and (_21311_, _21310_, _21302_);
  and (_21312_, _21311_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _21312_, _21294_);
  and (_21313_, _18672_, word_in[19]);
  and (_21314_, _20774_, _18466_);
  and (_21315_, _20778_, _18456_);
  or (_21316_, _21315_, _21314_);
  and (_21317_, _20769_, _18450_);
  and (_21318_, _20782_, _18447_);
  or (_21319_, _21318_, _21317_);
  or (_21320_, _21319_, _21316_);
  or (_21321_, _21320_, _18613_);
  and (_21322_, _20757_, _18456_);
  and (_21323_, _20753_, _18466_);
  or (_21324_, _21323_, _21322_);
  and (_21325_, _20762_, _18447_);
  and (_21326_, _20747_, _18450_);
  or (_21327_, _21326_, _21325_);
  nor (_21328_, _21327_, _21324_);
  nand (_21329_, _21328_, _18613_);
  and (_21330_, _21329_, _21321_);
  and (_21331_, _21330_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _21331_, _21313_);
  and (_21332_, _18672_, word_in[20]);
  and (_21333_, _20824_, _18456_);
  and (_21334_, _20820_, _18466_);
  or (_21335_, _21334_, _21333_);
  and (_21336_, _20828_, _18447_);
  and (_21337_, _20815_, _18450_);
  or (_21338_, _21337_, _21336_);
  or (_21339_, _21338_, _21335_);
  or (_21340_, _21339_, _18613_);
  and (_21341_, _20799_, _18466_);
  and (_21342_, _20803_, _18456_);
  or (_21343_, _21342_, _21341_);
  and (_21344_, _20793_, _18450_);
  and (_21345_, _20808_, _18447_);
  or (_21346_, _21345_, _21344_);
  nor (_21347_, _21346_, _21343_);
  nand (_21348_, _21347_, _18613_);
  and (_21349_, _21348_, _21340_);
  and (_21350_, _21349_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _21350_, _21332_);
  and (_21351_, _18672_, word_in[21]);
  and (_21352_, _20866_, _18466_);
  and (_21353_, _20870_, _18456_);
  or (_21354_, _21353_, _21352_);
  and (_21355_, _20861_, _18450_);
  and (_21356_, _20874_, _18447_);
  or (_21357_, _21356_, _21355_);
  or (_21358_, _21357_, _21354_);
  or (_21359_, _21358_, _18613_);
  and (_21360_, _20845_, _18466_);
  and (_21361_, _20849_, _18456_);
  or (_21362_, _21361_, _21360_);
  and (_21363_, _20839_, _18450_);
  and (_21364_, _20854_, _18447_);
  or (_21365_, _21364_, _21363_);
  nor (_21366_, _21365_, _21362_);
  nand (_21367_, _21366_, _18613_);
  and (_21368_, _21367_, _21359_);
  and (_21369_, _21368_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _21369_, _21351_);
  and (_21370_, _18672_, word_in[22]);
  and (_21371_, _20916_, _18466_);
  and (_21372_, _20912_, _18456_);
  or (_21373_, _21372_, _21371_);
  and (_21374_, _20907_, _18450_);
  and (_21375_, _20921_, _18447_);
  or (_21376_, _21375_, _21374_);
  or (_21377_, _21376_, _21373_);
  or (_21378_, _21377_, _18613_);
  and (_21379_, _20895_, _18456_);
  and (_21380_, _20891_, _18466_);
  or (_21381_, _21380_, _21379_);
  and (_21382_, _20900_, _18447_);
  and (_21383_, _20885_, _18450_);
  or (_21384_, _21383_, _21382_);
  nor (_21385_, _21384_, _21381_);
  nand (_21386_, _21385_, _18613_);
  and (_21387_, _21386_, _21378_);
  and (_21388_, _21387_, _18671_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _21388_, _21370_);
  and (_21389_, _18741_, word_in[24]);
  and (_21390_, _20966_, _18555_);
  and (_21391_, _20962_, _18561_);
  or (_21392_, _21391_, _21390_);
  and (_21393_, _21392_, _18699_);
  and (_21394_, _20956_, _18555_);
  and (_21395_, _20952_, _18561_);
  nor (_21396_, _21395_, _21394_);
  nor (_21397_, _21396_, _18699_);
  or (_21398_, _21397_, _21393_);
  and (_21399_, _21398_, _18695_);
  and (_21400_, _20944_, _18555_);
  and (_21401_, _20940_, _18561_);
  or (_21402_, _21401_, _21400_);
  and (_21403_, _21402_, _18699_);
  and (_21404_, _20930_, _18561_);
  and (_21405_, _20934_, _18555_);
  nor (_21406_, _21405_, _21404_);
  nor (_21407_, _21406_, _18699_);
  or (_21408_, _21407_, _21403_);
  and (_21409_, _21408_, _18752_);
  nor (_21410_, _21409_, _21399_);
  nor (_21411_, _21410_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _21411_, _21389_);
  and (_21412_, _18741_, word_in[25]);
  and (_21413_, _21013_, _18555_);
  and (_21414_, _21009_, _18561_);
  or (_21415_, _21414_, _21413_);
  and (_21416_, _21415_, _18699_);
  and (_21417_, _20999_, _18561_);
  and (_21418_, _21003_, _18555_);
  nor (_21419_, _21418_, _21417_);
  nor (_21420_, _21419_, _18699_);
  or (_21421_, _21420_, _21416_);
  and (_21422_, _21421_, _18695_);
  and (_21423_, _20991_, _18555_);
  and (_21424_, _20987_, _18561_);
  or (_21425_, _21424_, _21423_);
  and (_21426_, _21425_, _18699_);
  and (_21427_, _20977_, _18561_);
  and (_21428_, _20981_, _18555_);
  nor (_21429_, _21428_, _21427_);
  nor (_21430_, _21429_, _18699_);
  or (_21431_, _21430_, _21426_);
  and (_21432_, _21431_, _18752_);
  nor (_21433_, _21432_, _21422_);
  nor (_21434_, _21433_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _21434_, _21412_);
  and (_21435_, _18741_, word_in[26]);
  and (_21436_, _21060_, _18555_);
  and (_21437_, _21056_, _18561_);
  or (_21438_, _21437_, _21436_);
  and (_21439_, _21438_, _18699_);
  and (_21440_, _21046_, _18561_);
  and (_21441_, _21050_, _18555_);
  nor (_21442_, _21441_, _21440_);
  nor (_21443_, _21442_, _18699_);
  or (_21444_, _21443_, _21439_);
  and (_21445_, _21444_, _18695_);
  and (_21446_, _21038_, _18555_);
  and (_21447_, _21034_, _18561_);
  or (_21448_, _21447_, _21446_);
  and (_21449_, _21448_, _18699_);
  and (_21450_, _21024_, _18561_);
  and (_21451_, _21028_, _18555_);
  nor (_21452_, _21451_, _21450_);
  nor (_21453_, _21452_, _18699_);
  or (_21454_, _21453_, _21449_);
  and (_21455_, _21454_, _18752_);
  nor (_21456_, _21455_, _21445_);
  nor (_21457_, _21456_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _21457_, _21435_);
  and (_21458_, _18741_, word_in[27]);
  and (_21459_, _21107_, _18555_);
  and (_21460_, _21103_, _18561_);
  or (_21461_, _21460_, _21459_);
  and (_21462_, _21461_, _18699_);
  and (_21463_, _21093_, _18561_);
  and (_21464_, _21097_, _18555_);
  nor (_21465_, _21464_, _21463_);
  nor (_21466_, _21465_, _18699_);
  or (_21467_, _21466_, _21462_);
  and (_21468_, _21467_, _18695_);
  and (_21469_, _21075_, _18555_);
  and (_21470_, _21071_, _18561_);
  nor (_21471_, _21470_, _21469_);
  nor (_21472_, _21471_, _18699_);
  and (_21473_, _21085_, _18555_);
  and (_21474_, _21081_, _18561_);
  or (_21475_, _21474_, _21473_);
  and (_21476_, _21475_, _18699_);
  or (_21477_, _21476_, _21472_);
  and (_21478_, _21477_, _18752_);
  nor (_21479_, _21478_, _21468_);
  nor (_21480_, _21479_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _21480_, _21458_);
  and (_21481_, _18741_, word_in[28]);
  and (_21482_, _21154_, _18555_);
  and (_21483_, _21150_, _18561_);
  or (_21484_, _21483_, _21482_);
  and (_21485_, _21484_, _18699_);
  and (_21486_, _21140_, _18561_);
  and (_21487_, _21144_, _18555_);
  nor (_21488_, _21487_, _21486_);
  nor (_21489_, _21488_, _18699_);
  or (_21490_, _21489_, _21485_);
  and (_21491_, _21490_, _18695_);
  and (_21492_, _21132_, _18555_);
  and (_21493_, _21128_, _18561_);
  or (_21494_, _21493_, _21492_);
  and (_21495_, _21494_, _18699_);
  and (_21496_, _21118_, _18561_);
  and (_21497_, _21122_, _18555_);
  nor (_21498_, _21497_, _21496_);
  nor (_21499_, _21498_, _18699_);
  or (_21500_, _21499_, _21495_);
  and (_21501_, _21500_, _18752_);
  nor (_21502_, _21501_, _21491_);
  nor (_21503_, _21502_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _21503_, _21481_);
  and (_21504_, _18741_, word_in[29]);
  and (_21505_, _21201_, _18555_);
  and (_21506_, _21197_, _18561_);
  or (_21507_, _21506_, _21505_);
  and (_21508_, _21507_, _18699_);
  and (_21509_, _21187_, _18561_);
  and (_21510_, _21191_, _18555_);
  nor (_21511_, _21510_, _21509_);
  nor (_21512_, _21511_, _18699_);
  or (_21513_, _21512_, _21508_);
  and (_21514_, _21513_, _18695_);
  and (_21515_, _21179_, _18555_);
  and (_21516_, _21175_, _18561_);
  or (_21517_, _21516_, _21515_);
  and (_21518_, _21517_, _18699_);
  and (_21519_, _21165_, _18561_);
  and (_21520_, _21169_, _18555_);
  nor (_21521_, _21520_, _21519_);
  nor (_21522_, _21521_, _18699_);
  or (_21523_, _21522_, _21518_);
  and (_21524_, _21523_, _18752_);
  nor (_21525_, _21524_, _21514_);
  nor (_21526_, _21525_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _21526_, _21504_);
  and (_21527_, _18741_, word_in[30]);
  and (_21528_, _21248_, _18555_);
  and (_21529_, _21244_, _18561_);
  or (_21530_, _21529_, _21528_);
  and (_21531_, _21530_, _18699_);
  and (_21532_, _21238_, _18555_);
  and (_21533_, _21234_, _18561_);
  nor (_21534_, _21533_, _21532_);
  nor (_21535_, _21534_, _18699_);
  or (_21536_, _21535_, _21531_);
  and (_21537_, _21536_, _18695_);
  and (_21538_, _21226_, _18555_);
  and (_21539_, _21222_, _18561_);
  or (_21540_, _21539_, _21538_);
  and (_21541_, _21540_, _18699_);
  and (_21542_, _21212_, _18561_);
  and (_21543_, _21216_, _18555_);
  nor (_21544_, _21543_, _21542_);
  nor (_21545_, _21544_, _18699_);
  or (_21546_, _21545_, _21541_);
  and (_21547_, _21546_, _18752_);
  nor (_21548_, _21547_, _21537_);
  nor (_21549_, _21548_, _18741_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _21549_, _21527_);
  and (_21550_, _15585_, iram_op1[6]);
  and (_21551_, _15589_, iram_op1_reg[6]);
  or (_21552_, _21551_, _21550_);
  and (_00004_[6], _21552_, _38997_);
  and (_21553_, _15585_, iram_op1[5]);
  and (_21554_, _15589_, iram_op1_reg[5]);
  or (_21555_, _21554_, _21553_);
  and (_00004_[5], _21555_, _38997_);
  and (_21556_, _15585_, iram_op1[4]);
  and (_21557_, _15589_, iram_op1_reg[4]);
  or (_21558_, _21557_, _21556_);
  and (_00004_[4], _21558_, _38997_);
  and (_21559_, _15585_, iram_op1[3]);
  and (_21560_, _15589_, iram_op1_reg[3]);
  or (_21561_, _21560_, _21559_);
  and (_00004_[3], _21561_, _38997_);
  and (_21562_, _15585_, iram_op1[2]);
  and (_21563_, _15589_, iram_op1_reg[2]);
  or (_21564_, _21563_, _21562_);
  and (_00004_[2], _21564_, _38997_);
  and (_21565_, _15585_, iram_op1[1]);
  not (_21566_, iram_op1_reg[1]);
  nor (_21567_, _15585_, _21566_);
  or (_21568_, _21567_, _21565_);
  and (_00004_[1], _21568_, _38997_);
  and (_21569_, _15585_, iram_op1[0]);
  not (_21570_, iram_op1_reg[0]);
  nor (_21571_, _15585_, _21570_);
  or (_21572_, _21571_, _21569_);
  and (_00004_[0], _21572_, _38997_);
  and (_21573_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not (_21574_, pc_change_r);
  and (_21575_, _21574_, acc_reg[6]);
  or (_21576_, _21575_, _21573_);
  and (_00000_[6], _21576_, _38997_);
  and (_21577_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_21578_, _21574_, acc_reg[5]);
  or (_21579_, _21578_, _21577_);
  and (_00000_[5], _21579_, _38997_);
  and (_21580_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_21581_, _21574_, acc_reg[4]);
  or (_21582_, _21581_, _21580_);
  and (_00000_[4], _21582_, _38997_);
  and (_21583_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_21584_, _21574_, acc_reg[3]);
  or (_21585_, _21584_, _21583_);
  and (_00000_[3], _21585_, _38997_);
  and (_21586_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_21587_, _21574_, acc_reg[2]);
  or (_21588_, _21587_, _21586_);
  and (_00000_[2], _21588_, _38997_);
  and (_21589_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_21590_, _21574_, acc_reg[1]);
  or (_21591_, _21590_, _21589_);
  and (_00000_[1], _21591_, _38997_);
  and (_21592_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_21593_, _21574_, acc_reg[0]);
  or (_21594_, _21593_, _21592_);
  and (_00000_[0], _21594_, _38997_);
  and (_21595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_21596_, _21595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21597_, _21596_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21598_, _21596_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21599_, _21598_, _21597_);
  not (_21600_, _21599_);
  nor (_21601_, _21595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_21602_, _21596_, _21601_);
  and (_21603_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _16190_);
  and (_21604_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_21605_, _16194_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_21606_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_21607_, _21606_, _21604_);
  nor (_21608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_21609_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_21610_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_21611_, _21610_, _21609_);
  and (_21612_, _21611_, _21607_);
  nor (_21613_, _21612_, _21602_);
  not (_21614_, _21602_);
  and (_21615_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_21616_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_21617_, _21616_, _21615_);
  and (_21618_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_21619_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_21620_, _21619_, _21618_);
  and (_21621_, _21620_, _21617_);
  nor (_21622_, _21621_, _21614_);
  or (_21623_, _21622_, _21613_);
  and (_21624_, _21623_, _21600_);
  and (_21625_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_21626_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_21627_, _21626_, _21625_);
  and (_21628_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_21629_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_21630_, _21629_, _21628_);
  and (_21631_, _21630_, _21627_);
  nor (_21632_, _21631_, _21602_);
  and (_21633_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_21634_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_21635_, _21634_, _21633_);
  and (_21636_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_21637_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_21638_, _21637_, _21636_);
  and (_21639_, _21638_, _21635_);
  nor (_21640_, _21639_, _21614_);
  nor (_21641_, _21640_, _21632_);
  nor (_21642_, _21641_, _21600_);
  nor (_21643_, _21642_, _21624_);
  not (_21644_, _21643_);
  not (_21645_, _21603_);
  nor (_21646_, _21599_, _18609_);
  and (_21647_, _21599_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_21648_, _21647_, _21646_);
  nor (_21649_, _21648_, _21645_);
  or (_21650_, _21649_, _21602_);
  not (_21651_, _21595_);
  nor (_21652_, _21599_, _18657_);
  and (_21653_, _21599_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_21654_, _21653_, _21652_);
  nor (_21655_, _21654_, _21651_);
  not (_21656_, _21608_);
  nor (_21657_, _21599_, _18635_);
  and (_21658_, _21599_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_21659_, _21658_, _21657_);
  nor (_21660_, _21659_, _21656_);
  not (_21661_, _21605_);
  nor (_21662_, _21599_, _18644_);
  and (_21663_, _21599_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_21664_, _21663_, _21662_);
  nor (_21665_, _21664_, _21661_);
  or (_21666_, _21665_, _21660_);
  or (_21667_, _21666_, _21655_);
  or (_21668_, _21667_, _21650_);
  and (_21669_, _21599_, _18622_);
  nor (_21670_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21671_, _21670_, _21645_);
  nor (_21672_, _21671_, _21669_);
  or (_21673_, _21672_, _21614_);
  and (_21674_, _21599_, _18663_);
  nor (_21675_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21676_, _21675_, _21651_);
  nor (_21677_, _21676_, _21674_);
  and (_21678_, _21599_, _18630_);
  nor (_21679_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21680_, _21679_, _21656_);
  nor (_21681_, _21680_, _21678_);
  and (_21682_, _21599_, _18651_);
  nor (_21683_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21684_, _21683_, _21661_);
  nor (_21685_, _21684_, _21682_);
  or (_21686_, _21685_, _21681_);
  or (_21687_, _21686_, _21677_);
  or (_21688_, _21687_, _21673_);
  and (_21689_, _21688_, _21668_);
  and (_21690_, _21689_, _21644_);
  or (_21691_, _21690_, _15589_);
  or (_21692_, _15585_, op1_out_r[6]);
  and (_21693_, _21692_, _38997_);
  and (_00005_[6], _21693_, _21691_);
  and (_21694_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_21695_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_21696_, _21695_, _21694_);
  and (_21697_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_21698_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_21699_, _21698_, _21697_);
  and (_21700_, _21699_, _21696_);
  and (_21701_, _21700_, _21614_);
  and (_21702_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_21703_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_21704_, _21703_, _21702_);
  and (_21705_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_21706_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_21707_, _21706_, _21705_);
  and (_21708_, _21707_, _21704_);
  and (_21709_, _21708_, _21602_);
  or (_21710_, _21709_, _21599_);
  nor (_21711_, _21710_, _21701_);
  and (_21712_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_21713_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_21714_, _21713_, _21712_);
  and (_21715_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_21716_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_21717_, _21716_, _21715_);
  and (_21718_, _21717_, _21714_);
  nor (_21719_, _21718_, _21602_);
  and (_21720_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_21721_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_21722_, _21721_, _21720_);
  and (_21723_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_21724_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_21725_, _21724_, _21723_);
  and (_21726_, _21725_, _21722_);
  nor (_21727_, _21726_, _21614_);
  or (_21728_, _21727_, _21719_);
  and (_21729_, _21728_, _21599_);
  nor (_21730_, _21729_, _21711_);
  not (_21731_, _21730_);
  and (_21732_, _21731_, _21689_);
  or (_21733_, _21732_, _15589_);
  or (_21734_, _15585_, op1_out_r[5]);
  and (_21735_, _21734_, _38997_);
  and (_00005_[5], _21735_, _21733_);
  and (_21736_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_21737_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_21738_, _21737_, _21736_);
  and (_21739_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_21740_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_21741_, _21740_, _21739_);
  and (_21742_, _21741_, _21738_);
  and (_21743_, _21742_, _21614_);
  and (_21744_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_21745_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_21746_, _21745_, _21744_);
  and (_21747_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_21748_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_21749_, _21748_, _21747_);
  and (_21750_, _21749_, _21746_);
  and (_21751_, _21750_, _21602_);
  or (_21752_, _21751_, _21599_);
  nor (_21753_, _21752_, _21743_);
  and (_21754_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_21755_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_21756_, _21755_, _21754_);
  and (_21757_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_21758_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_21759_, _21758_, _21757_);
  and (_21760_, _21759_, _21756_);
  and (_21761_, _21760_, _21614_);
  and (_21762_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_21763_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_21764_, _21763_, _21762_);
  and (_21765_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_21766_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_21767_, _21766_, _21765_);
  and (_21768_, _21767_, _21764_);
  and (_21769_, _21768_, _21602_);
  or (_21770_, _21769_, _21600_);
  nor (_21771_, _21770_, _21761_);
  nor (_21772_, _21771_, _21753_);
  not (_21773_, _21772_);
  and (_21774_, _21773_, _21689_);
  or (_21775_, _21774_, _15589_);
  or (_21776_, _15585_, op1_out_r[4]);
  and (_21777_, _21776_, _38997_);
  and (_00005_[4], _21777_, _21775_);
  and (_21778_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_21779_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_21780_, _21779_, _21778_);
  and (_21781_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_21782_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_21783_, _21782_, _21781_);
  and (_21784_, _21783_, _21780_);
  nor (_21785_, _21784_, _21602_);
  and (_21786_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_21787_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_21788_, _21787_, _21786_);
  and (_21789_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_21790_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_21791_, _21790_, _21789_);
  and (_21792_, _21791_, _21788_);
  nor (_21793_, _21792_, _21614_);
  or (_21794_, _21793_, _21785_);
  and (_21795_, _21794_, _21600_);
  and (_21796_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_21797_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_21798_, _21797_, _21796_);
  and (_21799_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_21800_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_21801_, _21800_, _21799_);
  and (_21802_, _21801_, _21798_);
  nor (_21803_, _21802_, _21602_);
  and (_21804_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_21805_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_21806_, _21805_, _21804_);
  and (_21807_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_21808_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_21809_, _21808_, _21807_);
  and (_21810_, _21809_, _21806_);
  nor (_21811_, _21810_, _21614_);
  or (_21812_, _21811_, _21803_);
  and (_21813_, _21812_, _21599_);
  nor (_21814_, _21813_, _21795_);
  not (_21815_, _21814_);
  and (_21816_, _21815_, _21689_);
  or (_21817_, _21816_, _15589_);
  or (_21818_, _15585_, op1_out_r[3]);
  and (_21819_, _21818_, _38997_);
  and (_00005_[3], _21819_, _21817_);
  and (_21820_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_21821_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_21822_, _21821_, _21820_);
  and (_21823_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_21824_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_21825_, _21824_, _21823_);
  and (_21826_, _21825_, _21822_);
  and (_21827_, _21826_, _21602_);
  and (_21828_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_21829_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_21830_, _21829_, _21828_);
  and (_21831_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_21832_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_21833_, _21832_, _21831_);
  and (_21834_, _21833_, _21830_);
  and (_21835_, _21834_, _21614_);
  nor (_21836_, _21835_, _21827_);
  nor (_21837_, _21836_, _21600_);
  and (_21838_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_21839_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_21840_, _21839_, _21838_);
  and (_21841_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_21842_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_21843_, _21842_, _21841_);
  and (_21844_, _21843_, _21840_);
  and (_21845_, _21844_, _21614_);
  and (_21846_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_21847_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_21848_, _21847_, _21846_);
  and (_21849_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_21850_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_21851_, _21850_, _21849_);
  and (_21852_, _21851_, _21848_);
  and (_21853_, _21852_, _21602_);
  nor (_21854_, _21853_, _21845_);
  nor (_21855_, _21854_, _21599_);
  nor (_21856_, _21855_, _21837_);
  and (_21857_, _21856_, _21689_);
  or (_21858_, _21857_, _15589_);
  or (_21859_, _15585_, op1_out_r[2]);
  and (_21860_, _21859_, _38997_);
  and (_00005_[2], _21860_, _21858_);
  and (_21861_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_21862_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_21863_, _21862_, _21861_);
  and (_21864_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_21865_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_21866_, _21865_, _21864_);
  and (_21867_, _21866_, _21863_);
  and (_21868_, _21867_, _21614_);
  and (_21869_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_21870_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_21871_, _21870_, _21869_);
  and (_21872_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_21873_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_21874_, _21873_, _21872_);
  and (_21875_, _21874_, _21871_);
  and (_21876_, _21875_, _21602_);
  nor (_21877_, _21876_, _21868_);
  nor (_21878_, _21877_, _21600_);
  and (_21879_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_21880_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_21881_, _21880_, _21879_);
  and (_21882_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_21883_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_21884_, _21883_, _21882_);
  and (_21885_, _21884_, _21881_);
  and (_21886_, _21885_, _21614_);
  and (_21887_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_21888_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_21889_, _21888_, _21887_);
  and (_21890_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_21891_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_21892_, _21891_, _21890_);
  and (_21893_, _21892_, _21889_);
  and (_21894_, _21893_, _21602_);
  nor (_21895_, _21894_, _21886_);
  nor (_21896_, _21895_, _21599_);
  nor (_21897_, _21896_, _21878_);
  and (_21898_, _21897_, _21689_);
  or (_21899_, _21898_, _15589_);
  or (_21900_, _15585_, op1_out_r[1]);
  and (_21901_, _21900_, _38997_);
  and (_00005_[1], _21901_, _21899_);
  and (_21902_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_21903_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_21904_, _21903_, _21902_);
  and (_21905_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_21906_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_21907_, _21906_, _21905_);
  and (_21908_, _21907_, _21904_);
  and (_21909_, _21908_, _21614_);
  and (_21910_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_21911_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_21912_, _21911_, _21910_);
  and (_21913_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_21914_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_21915_, _21914_, _21913_);
  and (_21916_, _21915_, _21912_);
  and (_21917_, _21916_, _21602_);
  or (_21918_, _21917_, _21599_);
  nor (_21919_, _21918_, _21909_);
  and (_21920_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_21921_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_21922_, _21921_, _21920_);
  and (_21923_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_21924_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_21925_, _21924_, _21923_);
  and (_21926_, _21925_, _21922_);
  and (_21927_, _21926_, _21614_);
  and (_21928_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_21929_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_21930_, _21929_, _21928_);
  and (_21931_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_21932_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_21933_, _21932_, _21931_);
  and (_21934_, _21933_, _21930_);
  and (_21935_, _21934_, _21602_);
  or (_21936_, _21935_, _21600_);
  nor (_21937_, _21936_, _21927_);
  nor (_21938_, _21937_, _21919_);
  not (_21939_, _21938_);
  and (_21940_, _21939_, _21689_);
  or (_21941_, _21940_, _15589_);
  or (_21942_, _15585_, op1_out_r[0]);
  and (_21943_, _21942_, _38997_);
  and (_00005_[0], _21943_, _21941_);
  and (_21944_, _15589_, iram_op1[6]);
  and (_21945_, _21774_, _21732_);
  and (_21946_, _21605_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_21947_, _21595_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_21948_, _21947_, _21946_);
  and (_21949_, _21603_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_21950_, _21608_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_21951_, _21950_, _21949_);
  and (_21952_, _21951_, _21948_);
  and (_21953_, _21952_, _21614_);
  and (_21954_, _21605_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_21955_, _21595_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_21956_, _21955_, _21954_);
  and (_21957_, _21603_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_21958_, _21608_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_21959_, _21958_, _21957_);
  and (_21960_, _21959_, _21956_);
  and (_21961_, _21960_, _21602_);
  nor (_21962_, _21961_, _21953_);
  nor (_21963_, _21962_, _21600_);
  and (_21964_, _21605_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_21965_, _21603_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_21966_, _21965_, _21964_);
  and (_21967_, _21608_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_21968_, _21595_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_21969_, _21968_, _21967_);
  and (_21970_, _21969_, _21966_);
  and (_21971_, _21970_, _21614_);
  and (_21972_, _21603_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_21973_, _21608_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_21974_, _21973_, _21972_);
  and (_21975_, _21605_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_21976_, _21595_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_21977_, _21976_, _21975_);
  and (_21978_, _21977_, _21974_);
  and (_21979_, _21978_, _21602_);
  nor (_21980_, _21979_, _21971_);
  nor (_21981_, _21980_, _21599_);
  nor (_21982_, _21981_, _21963_);
  and (_21983_, _21982_, _21689_);
  and (_21984_, _21983_, _21690_);
  and (_21985_, _21984_, _21945_);
  nor (_21986_, _21857_, _21816_);
  and (_21987_, _21938_, _21898_);
  and (_21988_, _21987_, _21986_);
  and (_21989_, _21988_, _21985_);
  and (_21990_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  not (_21991_, _21898_);
  and (_21992_, _21940_, _21991_);
  and (_21993_, _21986_, _21992_);
  and (_21994_, _21993_, _21985_);
  and (_21995_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_21996_, _21995_, _21990_);
  nor (_21997_, _21940_, _21898_);
  and (_21998_, _21986_, _21997_);
  and (_21999_, _21998_, _21985_);
  and (_22000_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_22001_, _21857_, _21816_);
  and (_22002_, _21940_, _21898_);
  and (_22003_, _22002_, _22001_);
  and (_22004_, _21772_, _21732_);
  and (_22005_, _22004_, _21984_);
  and (_22006_, _22005_, _22003_);
  and (_22007_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or (_22008_, _22007_, _22000_);
  or (_22009_, _22008_, _21996_);
  not (_22010_, _21816_);
  and (_22011_, _21857_, _22010_);
  and (_22012_, _22011_, _21992_);
  and (_22013_, _22012_, _21985_);
  and (_22014_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and (_22015_, _21987_, _22011_);
  and (_22016_, _22015_, _21985_);
  and (_22017_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_22018_, _22017_, _22014_);
  and (_22019_, _22011_, _21997_);
  and (_22020_, _22019_, _21985_);
  and (_22021_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_22022_, _21986_, _22002_);
  and (_22023_, _22022_, _21985_);
  and (_22024_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or (_22025_, _22024_, _22021_);
  or (_22026_, _22025_, _22018_);
  or (_22027_, _22026_, _22009_);
  and (_22028_, _21987_, _22001_);
  and (_22029_, _22028_, _21985_);
  and (_22030_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_22031_, _21992_, _22001_);
  and (_22032_, _22031_, _21985_);
  and (_22033_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or (_22034_, _22033_, _22030_);
  and (_22035_, _22001_, _21997_);
  and (_22036_, _22035_, _21985_);
  and (_22037_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor (_22038_, _21857_, _22010_);
  and (_22039_, _22002_, _22038_);
  and (_22040_, _22039_, _21985_);
  and (_22041_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_22042_, _22041_, _22037_);
  or (_22043_, _22042_, _22034_);
  and (_22044_, _21987_, _22038_);
  and (_22045_, _22044_, _21985_);
  and (_22046_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_22047_, _21992_, _22038_);
  and (_22048_, _22047_, _21985_);
  and (_22049_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or (_22050_, _22049_, _22046_);
  and (_22051_, _22038_, _21997_);
  and (_22052_, _22051_, _21985_);
  and (_22053_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  and (_22054_, _22011_, _22002_);
  and (_22055_, _22054_, _21985_);
  and (_22056_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or (_22057_, _22056_, _22053_);
  or (_22058_, _22057_, _22050_);
  or (_22059_, _22058_, _22043_);
  or (_22060_, _22059_, _22027_);
  and (_22061_, _22005_, _21993_);
  and (_22062_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_22063_, _22005_, _21988_);
  and (_22064_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or (_22065_, _22064_, _22062_);
  and (_22066_, _21774_, _21730_);
  and (_22067_, _22066_, _21984_);
  and (_22068_, _22067_, _22003_);
  and (_22069_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and (_22070_, _22005_, _21998_);
  and (_22071_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_22072_, _22071_, _22069_);
  or (_22073_, _22072_, _22065_);
  and (_22074_, _22005_, _22015_);
  and (_22075_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_22076_, _22005_, _22012_);
  and (_22077_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or (_22078_, _22077_, _22075_);
  and (_22079_, _22005_, _22022_);
  and (_22080_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  and (_22081_, _22005_, _22019_);
  and (_22082_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_22083_, _22082_, _22080_);
  or (_22084_, _22083_, _22078_);
  or (_22085_, _22084_, _22073_);
  and (_22086_, _22005_, _22031_);
  and (_22087_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  and (_22088_, _22005_, _22028_);
  and (_22089_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_22090_, _22089_, _22087_);
  and (_22091_, _22005_, _22039_);
  and (_22092_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_22093_, _22005_, _22035_);
  and (_22094_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or (_22095_, _22094_, _22092_);
  or (_22096_, _22095_, _22090_);
  and (_22097_, _22005_, _22044_);
  and (_22098_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  and (_22099_, _22005_, _22047_);
  and (_22100_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_22101_, _22100_, _22098_);
  and (_22102_, _22005_, _22051_);
  and (_22103_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_22104_, _22005_, _22054_);
  and (_22105_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_22106_, _22105_, _22103_);
  or (_22107_, _22106_, _22101_);
  or (_22108_, _22107_, _22096_);
  or (_22109_, _22108_, _22085_);
  or (_22110_, _22109_, _22060_);
  and (_22111_, _22067_, _22028_);
  and (_22112_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_22113_, _22067_, _22031_);
  and (_22114_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  or (_22115_, _22114_, _22112_);
  and (_22116_, _22067_, _22039_);
  and (_22117_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and (_22118_, _22067_, _22035_);
  and (_22119_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_22120_, _22119_, _22117_);
  or (_22121_, _22120_, _22115_);
  and (_22122_, _22067_, _22044_);
  and (_22123_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_22124_, _22067_, _22047_);
  and (_22125_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  or (_22126_, _22125_, _22123_);
  and (_22127_, _22067_, _22051_);
  and (_22128_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and (_22129_, _22067_, _22054_);
  and (_22130_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  or (_22131_, _22130_, _22128_);
  or (_22132_, _22131_, _22126_);
  or (_22133_, _22132_, _22121_);
  and (_22134_, _22067_, _21993_);
  and (_22135_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and (_22136_, _22067_, _21988_);
  and (_22137_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_22138_, _22137_, _22135_);
  nor (_22139_, _21774_, _21732_);
  and (_22140_, _22139_, _21984_);
  and (_22141_, _22003_, _22140_);
  and (_22142_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_22143_, _22067_, _21998_);
  and (_22144_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  or (_22145_, _22144_, _22142_);
  or (_22146_, _22145_, _22138_);
  and (_22147_, _22067_, _22015_);
  and (_22148_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and (_22149_, _22067_, _22012_);
  and (_22150_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_22151_, _22150_, _22148_);
  and (_22152_, _22067_, _22019_);
  and (_22153_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_22154_, _22067_, _22022_);
  and (_22155_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  or (_22156_, _22155_, _22153_);
  or (_22157_, _22156_, _22151_);
  or (_22158_, _22157_, _22146_);
  or (_22159_, _22158_, _22133_);
  and (_22160_, _22031_, _22140_);
  and (_22161_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and (_22162_, _22028_, _22140_);
  and (_22163_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_22164_, _22163_, _22161_);
  and (_22165_, _22039_, _22140_);
  and (_22166_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_22167_, _22140_, _22035_);
  and (_22168_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_22169_, _22168_, _22166_);
  or (_22170_, _22169_, _22164_);
  and (_22171_, _22047_, _22140_);
  and (_22172_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  and (_22173_, _22044_, _22140_);
  and (_22174_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_22175_, _22174_, _22172_);
  and (_22176_, _22140_, _22051_);
  and (_22177_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_22178_, _22054_, _22140_);
  and (_22179_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_22180_, _22179_, _22177_);
  or (_22181_, _22180_, _22175_);
  or (_22182_, _22181_, _22170_);
  and (_22183_, _22015_, _22140_);
  and (_22184_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_22185_, _22012_, _22140_);
  and (_22186_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_22187_, _22186_, _22184_);
  and (_22188_, _22022_, _22140_);
  and (_22189_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  and (_22190_, _22019_, _22140_);
  and (_22191_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_22192_, _22191_, _22189_);
  or (_22193_, _22192_, _22187_);
  and (_22194_, _21988_, _22140_);
  and (_22195_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_22196_, _21993_, _22140_);
  and (_22197_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_22198_, _22197_, _22195_);
  not (_22199_, _21983_);
  nor (_22200_, _22199_, _21690_);
  and (_22201_, _22200_, _21945_);
  and (_22202_, _22201_, _22003_);
  and (_22203_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  and (_22204_, _21998_, _22140_);
  and (_22205_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_22206_, _22205_, _22203_);
  or (_22207_, _22206_, _22198_);
  or (_22208_, _22207_, _22193_);
  or (_22209_, _22208_, _22182_);
  or (_22210_, _22209_, _22159_);
  or (_22211_, _22210_, _22110_);
  and (_22212_, _22201_, _22012_);
  and (_22213_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  and (_22214_, _22201_, _22015_);
  and (_22215_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_22216_, _22215_, _22213_);
  and (_22217_, _22201_, _22019_);
  and (_22218_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_22219_, _22201_, _22022_);
  and (_22220_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or (_22221_, _22220_, _22218_);
  or (_22222_, _22221_, _22216_);
  and (_22223_, _22201_, _21993_);
  and (_22224_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  and (_22225_, _22201_, _21988_);
  and (_22226_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_22227_, _22226_, _22224_);
  and (_22228_, _22004_, _22200_);
  and (_22229_, _22003_, _22228_);
  and (_22230_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_22231_, _22201_, _21998_);
  and (_22232_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or (_22233_, _22232_, _22230_);
  or (_22234_, _22233_, _22227_);
  or (_22235_, _22234_, _22222_);
  and (_22236_, _22201_, _22044_);
  and (_22237_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_22238_, _22201_, _22047_);
  and (_22239_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or (_22240_, _22239_, _22237_);
  and (_22241_, _22201_, _22051_);
  and (_22242_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  and (_22243_, _22201_, _22054_);
  and (_22244_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or (_22245_, _22244_, _22242_);
  or (_22246_, _22245_, _22240_);
  and (_22247_, _22201_, _22028_);
  and (_22248_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_22249_, _22201_, _22031_);
  and (_22250_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or (_22251_, _22250_, _22248_);
  and (_22252_, _22201_, _22039_);
  and (_22253_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  and (_22254_, _22201_, _22035_);
  and (_22255_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_22256_, _22255_, _22253_);
  or (_22257_, _22256_, _22251_);
  or (_22258_, _22257_, _22246_);
  or (_22259_, _22258_, _22235_);
  and (_22260_, _22047_, _22228_);
  and (_22261_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and (_22262_, _22044_, _22228_);
  and (_22263_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_22264_, _22263_, _22261_);
  and (_22265_, _22054_, _22228_);
  and (_22266_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_22267_, _22228_, _22051_);
  and (_22268_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  or (_22269_, _22268_, _22266_);
  or (_22270_, _22269_, _22264_);
  and (_22271_, _22228_, _22031_);
  and (_22272_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and (_22273_, _22028_, _22228_);
  and (_22274_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_22275_, _22274_, _22272_);
  and (_22276_, _22228_, _22039_);
  and (_22277_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_22278_, _22228_, _22035_);
  and (_22279_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  or (_22280_, _22279_, _22277_);
  or (_22281_, _22280_, _22275_);
  or (_22282_, _22281_, _22270_);
  and (_22283_, _22012_, _22228_);
  and (_22284_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_22285_, _22015_, _22228_);
  and (_22286_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  or (_22287_, _22286_, _22284_);
  and (_22288_, _22022_, _22228_);
  and (_22289_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and (_22290_, _22019_, _22228_);
  and (_22291_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_22292_, _22291_, _22289_);
  or (_22293_, _22292_, _22287_);
  and (_22294_, _21988_, _22228_);
  and (_22295_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_22296_, _21993_, _22228_);
  and (_22297_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  or (_22298_, _22297_, _22295_);
  and (_22299_, _22066_, _22200_);
  and (_22300_, _22299_, _22003_);
  and (_22301_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  and (_22302_, _21998_, _22228_);
  and (_22303_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_22304_, _22303_, _22301_);
  or (_22305_, _22304_, _22298_);
  or (_22306_, _22305_, _22293_);
  or (_22307_, _22306_, _22282_);
  or (_22308_, _22307_, _22259_);
  and (_22309_, _22299_, _21988_);
  and (_22310_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  and (_22311_, _22299_, _21993_);
  and (_22312_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_22313_, _22312_, _22310_);
  and (_22314_, _22299_, _21998_);
  and (_22315_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_22316_, _22200_, _22139_);
  and (_22317_, _22003_, _22316_);
  and (_22318_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or (_22319_, _22318_, _22315_);
  or (_22320_, _22319_, _22313_);
  and (_22321_, _22299_, _22015_);
  and (_22322_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  and (_22323_, _22299_, _22012_);
  and (_22324_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_22325_, _22324_, _22322_);
  and (_22326_, _22299_, _22019_);
  and (_22327_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_22328_, _22299_, _22022_);
  and (_22329_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or (_22330_, _22329_, _22327_);
  or (_22331_, _22330_, _22325_);
  or (_22332_, _22331_, _22320_);
  and (_22333_, _22299_, _22031_);
  and (_22334_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_22335_, _22299_, _22028_);
  and (_22336_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or (_22337_, _22336_, _22334_);
  and (_22338_, _22299_, _22035_);
  and (_22339_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and (_22340_, _22299_, _22039_);
  and (_22341_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_22342_, _22341_, _22339_);
  or (_22343_, _22342_, _22337_);
  and (_22344_, _22299_, _22047_);
  and (_22345_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_22346_, _22299_, _22044_);
  and (_22347_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or (_22348_, _22347_, _22345_);
  and (_22349_, _22299_, _22051_);
  and (_22350_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and (_22351_, _22299_, _22054_);
  and (_22352_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or (_22353_, _22352_, _22350_);
  or (_22354_, _22353_, _22348_);
  or (_22355_, _22354_, _22343_);
  or (_22356_, _22355_, _22332_);
  and (_22357_, _21993_, _22316_);
  and (_22358_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  and (_22359_, _21988_, _22316_);
  and (_22360_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or (_22361_, _22360_, _22358_);
  and (_22362_, _21998_, _22316_);
  and (_22363_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and (_22364_, _22199_, _21690_);
  and (_22365_, _22364_, _21945_);
  and (_22366_, _22003_, _22365_);
  and (_22367_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_22368_, _22367_, _22363_);
  or (_22369_, _22368_, _22361_);
  and (_22370_, _22015_, _22316_);
  and (_22371_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  and (_22372_, _22012_, _22316_);
  and (_22373_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or (_22374_, _22373_, _22371_);
  and (_22375_, _22019_, _22316_);
  and (_22376_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and (_22377_, _22022_, _22316_);
  and (_22378_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_22379_, _22378_, _22376_);
  or (_22380_, _22379_, _22374_);
  or (_22381_, _22380_, _22369_);
  and (_22382_, _22031_, _22316_);
  and (_22383_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and (_22384_, _22028_, _22316_);
  and (_22385_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_22386_, _22385_, _22383_);
  and (_22387_, _22316_, _22035_);
  and (_22388_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  and (_22389_, _22039_, _22316_);
  and (_22390_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or (_22391_, _22390_, _22388_);
  or (_22392_, _22391_, _22386_);
  and (_22393_, _22044_, _22316_);
  and (_22394_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and (_22395_, _22047_, _22316_);
  and (_22396_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_22397_, _22396_, _22394_);
  and (_22398_, _22054_, _22316_);
  and (_22399_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and (_22400_, _22316_, _22051_);
  and (_22401_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or (_22402_, _22401_, _22399_);
  or (_22403_, _22402_, _22397_);
  or (_22404_, _22403_, _22392_);
  or (_22405_, _22404_, _22381_);
  or (_22406_, _22405_, _22356_);
  or (_22407_, _22406_, _22308_);
  or (_22408_, _22407_, _22211_);
  and (_22409_, _22365_, _22012_);
  and (_22410_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  and (_22411_, _22365_, _22015_);
  and (_22412_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_22413_, _22412_, _22410_);
  and (_22414_, _22365_, _22019_);
  and (_22415_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_22416_, _22365_, _22022_);
  and (_22417_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or (_22418_, _22417_, _22415_);
  or (_22419_, _22418_, _22413_);
  and (_22420_, _22365_, _21993_);
  and (_22421_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  and (_22422_, _21988_, _22365_);
  and (_22423_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_22424_, _22423_, _22421_);
  and (_22425_, _22364_, _22004_);
  and (_22426_, _22003_, _22425_);
  and (_22427_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_22428_, _22365_, _21998_);
  and (_22429_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or (_22430_, _22429_, _22427_);
  or (_22431_, _22430_, _22424_);
  or (_22432_, _22431_, _22419_);
  and (_22433_, _22365_, _22044_);
  and (_22434_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_22435_, _22365_, _22047_);
  and (_22436_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or (_22437_, _22436_, _22434_);
  and (_22438_, _22365_, _22054_);
  and (_22439_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_22440_, _22365_, _22051_);
  and (_22441_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_22442_, _22441_, _22439_);
  or (_22443_, _22442_, _22437_);
  and (_22444_, _22365_, _22028_);
  and (_22445_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_22446_, _22365_, _22031_);
  and (_22447_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or (_22448_, _22447_, _22445_);
  and (_22449_, _22365_, _22039_);
  and (_22450_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  and (_22451_, _22365_, _22035_);
  and (_22452_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_22453_, _22452_, _22450_);
  or (_22454_, _22453_, _22448_);
  or (_22455_, _22454_, _22443_);
  or (_22456_, _22455_, _22432_);
  and (_22457_, _22425_, _22028_);
  and (_22458_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  and (_22459_, _22425_, _22031_);
  and (_22460_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_22461_, _22460_, _22458_);
  and (_22462_, _22425_, _22035_);
  and (_22463_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_22464_, _22425_, _22039_);
  and (_22465_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_22466_, _22465_, _22463_);
  or (_22467_, _22466_, _22461_);
  and (_22468_, _22425_, _22044_);
  and (_22469_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  and (_22470_, _22425_, _22047_);
  and (_22471_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_22472_, _22471_, _22469_);
  and (_22473_, _22425_, _22051_);
  and (_22474_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_22475_, _22425_, _22054_);
  and (_22476_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_22477_, _22476_, _22474_);
  or (_22478_, _22477_, _22472_);
  or (_22479_, _22478_, _22467_);
  and (_22480_, _22425_, _22012_);
  and (_22481_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_22482_, _22425_, _22015_);
  and (_22483_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_22484_, _22483_, _22481_);
  and (_22485_, _22019_, _22425_);
  and (_22486_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  and (_22487_, _22425_, _22022_);
  and (_22488_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_22489_, _22488_, _22486_);
  or (_22490_, _22489_, _22484_);
  and (_22491_, _21988_, _22425_);
  and (_22492_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_22493_, _22425_, _21993_);
  and (_22494_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_22495_, _22494_, _22492_);
  and (_22496_, _21998_, _22425_);
  and (_22497_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  and (_22498_, _22364_, _22066_);
  and (_22499_, _22003_, _22498_);
  and (_22500_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_22501_, _22500_, _22497_);
  or (_22502_, _22501_, _22495_);
  or (_22503_, _22502_, _22490_);
  or (_22504_, _22503_, _22479_);
  or (_22505_, _22504_, _22456_);
  and (_22506_, _22012_, _22498_);
  and (_22507_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  and (_22508_, _22015_, _22498_);
  and (_22509_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_22510_, _22509_, _22507_);
  and (_22511_, _22019_, _22498_);
  and (_22512_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_22513_, _22022_, _22498_);
  and (_22514_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_22515_, _22514_, _22512_);
  or (_22516_, _22515_, _22510_);
  and (_22517_, _21988_, _22498_);
  and (_22518_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  and (_22519_, _21993_, _22498_);
  and (_22520_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_22521_, _22520_, _22518_);
  and (_22522_, _21998_, _22498_);
  and (_22523_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_22524_, _22364_, _22139_);
  and (_22525_, _22003_, _22524_);
  and (_22526_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_22527_, _22526_, _22523_);
  or (_22528_, _22527_, _22521_);
  or (_22529_, _22528_, _22516_);
  and (_22530_, _22044_, _22498_);
  and (_22531_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_22532_, _22047_, _22498_);
  and (_22533_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_22534_, _22533_, _22531_);
  and (_22535_, _22498_, _22054_);
  and (_22536_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_22537_, _22498_, _22051_);
  and (_22538_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_22539_, _22538_, _22536_);
  or (_22540_, _22539_, _22534_);
  and (_22541_, _22498_, _22039_);
  and (_22542_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  and (_22543_, _22498_, _22035_);
  and (_22544_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_22545_, _22544_, _22542_);
  and (_22546_, _22498_, _22031_);
  and (_22547_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_22548_, _22028_, _22498_);
  and (_22549_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_22550_, _22549_, _22547_);
  or (_22551_, _22550_, _22545_);
  or (_22552_, _22551_, _22540_);
  or (_22553_, _22552_, _22529_);
  and (_22554_, _22524_, _21993_);
  and (_22555_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_22556_, _22524_, _21988_);
  and (_22557_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_22558_, _22557_, _22555_);
  nor (_22559_, _21983_, _21690_);
  and (_22560_, _22559_, _21945_);
  and (_22561_, _22003_, _22560_);
  and (_22562_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  and (_22563_, _22524_, _21998_);
  and (_22564_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_22565_, _22564_, _22562_);
  or (_22566_, _22565_, _22558_);
  and (_22567_, _22524_, _22015_);
  and (_22568_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_22569_, _22524_, _22012_);
  and (_22570_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_22571_, _22570_, _22568_);
  and (_22572_, _22524_, _22022_);
  and (_22573_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  and (_22574_, _22524_, _22019_);
  and (_22575_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_22576_, _22575_, _22573_);
  or (_22577_, _22576_, _22571_);
  or (_22578_, _22577_, _22566_);
  and (_22579_, _22524_, _22044_);
  and (_22580_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  and (_22581_, _22524_, _22047_);
  and (_22582_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_22583_, _22582_, _22580_);
  and (_22584_, _22524_, _22054_);
  and (_22585_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and (_22586_, _22524_, _22051_);
  and (_22587_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_22588_, _22587_, _22585_);
  or (_22589_, _22588_, _22583_);
  and (_22590_, _22524_, _22031_);
  and (_22591_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  and (_22592_, _22524_, _22028_);
  and (_22593_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_22594_, _22593_, _22591_);
  and (_22595_, _22524_, _22035_);
  and (_22596_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_22597_, _22524_, _22039_);
  and (_22598_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_22599_, _22598_, _22596_);
  or (_22600_, _22599_, _22594_);
  or (_22601_, _22600_, _22589_);
  or (_22602_, _22601_, _22578_);
  or (_22603_, _22602_, _22553_);
  or (_22604_, _22603_, _22505_);
  and (_22605_, _22047_, _22560_);
  and (_22606_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_22607_, _22044_, _22560_);
  and (_22608_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_22609_, _22608_, _22606_);
  and (_22610_, _22560_, _22054_);
  and (_22611_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_22612_, _22560_, _22051_);
  and (_22613_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_22614_, _22613_, _22611_);
  or (_22615_, _22614_, _22609_);
  and (_22616_, _22028_, _22560_);
  and (_22617_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_22618_, _22560_, _22031_);
  and (_22619_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_22620_, _22619_, _22617_);
  and (_22621_, _22560_, _22039_);
  and (_22622_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  and (_22623_, _22560_, _22035_);
  and (_22624_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_22625_, _22624_, _22622_);
  or (_22626_, _22625_, _22620_);
  or (_22627_, _22626_, _22615_);
  and (_22628_, _22012_, _22560_);
  and (_22629_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  and (_22630_, _22015_, _22560_);
  and (_22631_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_22632_, _22631_, _22629_);
  and (_22633_, _22019_, _22560_);
  and (_22634_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_22635_, _22560_, _22022_);
  and (_22636_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_22637_, _22636_, _22634_);
  or (_22638_, _22637_, _22632_);
  and (_22639_, _21988_, _22560_);
  and (_22640_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  and (_22641_, _22560_, _21993_);
  and (_22642_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_22643_, _22642_, _22640_);
  and (_22644_, _21998_, _22560_);
  and (_22645_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_22646_, _22559_, _22004_);
  and (_22647_, _22003_, _22646_);
  and (_22648_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_22649_, _22648_, _22645_);
  or (_22650_, _22649_, _22643_);
  or (_22651_, _22650_, _22638_);
  or (_22652_, _22651_, _22627_);
  and (_22653_, _22646_, _22028_);
  and (_22654_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  and (_22655_, _22646_, _22031_);
  and (_22656_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_22657_, _22656_, _22654_);
  and (_22658_, _22646_, _22035_);
  and (_22659_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_22660_, _22646_, _22039_);
  and (_22661_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_22662_, _22661_, _22659_);
  or (_22663_, _22662_, _22657_);
  and (_22664_, _22047_, _22646_);
  and (_22665_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  and (_22666_, _22044_, _22646_);
  and (_22667_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_22668_, _22667_, _22665_);
  and (_22669_, _22646_, _22051_);
  and (_22670_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_22671_, _22646_, _22054_);
  and (_22672_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_22673_, _22672_, _22670_);
  or (_22674_, _22673_, _22668_);
  or (_22675_, _22674_, _22663_);
  and (_22676_, _22015_, _22646_);
  and (_22677_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_22678_, _22012_, _22646_);
  and (_22679_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_22680_, _22679_, _22677_);
  and (_22681_, _22019_, _22646_);
  and (_22682_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  and (_22683_, _22646_, _22022_);
  and (_22684_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_22685_, _22684_, _22682_);
  or (_22686_, _22685_, _22680_);
  and (_22687_, _21988_, _22646_);
  and (_22688_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_22689_, _22646_, _21993_);
  and (_22690_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_22691_, _22690_, _22688_);
  and (_22692_, _22559_, _22066_);
  and (_22693_, _22003_, _22692_);
  and (_22694_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  and (_22695_, _21998_, _22646_);
  and (_22696_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_22697_, _22696_, _22694_);
  or (_22698_, _22697_, _22691_);
  or (_22699_, _22698_, _22686_);
  or (_22700_, _22699_, _22675_);
  or (_22701_, _22700_, _22652_);
  and (_22702_, _22559_, _22139_);
  and (_22703_, _22012_, _22702_);
  and (_22704_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_22705_, _22015_, _22702_);
  and (_22706_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_22707_, _22706_, _22704_);
  and (_22708_, _22019_, _22702_);
  and (_22709_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_22710_, _22709_, _22707_);
  and (_22711_, _21988_, _22702_);
  and (_22712_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_22713_, _21998_, _22702_);
  and (_22714_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_22715_, _22714_, _22712_);
  and (_22716_, _22702_, _21993_);
  and (_22717_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_22718_, _22702_, _22022_);
  and (_22719_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_22720_, _22719_, _22717_);
  or (_22721_, _22720_, _22715_);
  or (_22722_, _22721_, _22710_);
  and (_22723_, _22044_, _22702_);
  and (_22724_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_22725_, _22047_, _22702_);
  and (_22726_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_22727_, _22726_, _22724_);
  and (_22728_, _22702_, _22051_);
  and (_22729_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_22730_, _22702_, _22054_);
  and (_22731_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_22732_, _22731_, _22729_);
  or (_22733_, _22732_, _22727_);
  and (_22734_, _22702_, _22031_);
  and (_22735_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_22736_, _22028_, _22702_);
  and (_22737_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_22738_, _22737_, _22735_);
  and (_22739_, _22702_, _22039_);
  and (_22740_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_22741_, _22702_, _22035_);
  and (_22742_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_22743_, _22742_, _22740_);
  or (_22744_, _22743_, _22738_);
  or (_22745_, _22744_, _22733_);
  or (_22746_, _22745_, _22722_);
  and (_22747_, _22692_, _22028_);
  and (_22748_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_22749_, _22692_, _22031_);
  and (_22750_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_22751_, _22750_, _22748_);
  and (_22752_, _22692_, _22035_);
  and (_22753_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  and (_22754_, _22692_, _22039_);
  and (_22755_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_22756_, _22755_, _22753_);
  or (_22757_, _22756_, _22751_);
  and (_22758_, _22692_, _22044_);
  and (_22759_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_22760_, _22692_, _22047_);
  and (_22761_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_22762_, _22761_, _22759_);
  and (_22763_, _22692_, _22051_);
  and (_22764_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  and (_22765_, _22692_, _22054_);
  and (_22766_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_22767_, _22766_, _22764_);
  or (_22768_, _22767_, _22762_);
  or (_22769_, _22768_, _22757_);
  and (_22770_, _22692_, _22015_);
  and (_22771_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  and (_22772_, _22692_, _22012_);
  and (_22773_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_22774_, _22773_, _22771_);
  and (_22775_, _22692_, _22022_);
  and (_22776_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_22777_, _22692_, _22019_);
  and (_22778_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_22779_, _22778_, _22776_);
  or (_22780_, _22779_, _22774_);
  and (_22781_, _22003_, _22702_);
  and (_22782_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_22783_, _22692_, _21998_);
  and (_22784_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_22785_, _22784_, _22782_);
  and (_22786_, _21988_, _22692_);
  and (_22787_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  and (_22788_, _22692_, _21993_);
  and (_22789_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_22790_, _22789_, _22787_);
  or (_22791_, _22790_, _22785_);
  or (_22792_, _22791_, _22780_);
  or (_22793_, _22792_, _22769_);
  or (_22794_, _22793_, _22746_);
  or (_22795_, _22794_, _22701_);
  or (_22796_, _22795_, _22604_);
  or (_22797_, _22796_, _22408_);
  nor (_22798_, _22032_, _22029_);
  nor (_22799_, _22040_, _22036_);
  and (_22800_, _22799_, _22798_);
  nor (_22801_, _22055_, _22052_);
  nor (_22802_, _22048_, _22045_);
  and (_22803_, _22802_, _22801_);
  and (_22804_, _22803_, _22800_);
  nor (_22805_, _22006_, _21999_);
  nor (_22806_, _21994_, _21989_);
  and (_22807_, _22806_, _22805_);
  nor (_22808_, _22016_, _22013_);
  nor (_22809_, _22023_, _22020_);
  and (_22810_, _22809_, _22808_);
  and (_22811_, _22810_, _22807_);
  and (_22812_, _22811_, _22804_);
  nor (_22813_, _22070_, _22061_);
  nor (_22814_, _22068_, _22063_);
  and (_22815_, _22814_, _22813_);
  nor (_22816_, _22081_, _22079_);
  nor (_22817_, _22076_, _22074_);
  and (_22818_, _22817_, _22816_);
  and (_22819_, _22818_, _22815_);
  nor (_22820_, _22099_, _22097_);
  nor (_22821_, _22104_, _22102_);
  and (_22822_, _22821_, _22820_);
  nor (_22823_, _22088_, _22086_);
  nor (_22824_, _22093_, _22091_);
  and (_22825_, _22824_, _22823_);
  and (_22826_, _22825_, _22822_);
  and (_22827_, _22826_, _22819_);
  and (_22828_, _22827_, _22812_);
  nor (_22829_, _22154_, _22152_);
  nor (_22830_, _22149_, _22147_);
  and (_22831_, _22830_, _22829_);
  nor (_22832_, _22136_, _22134_);
  nor (_22833_, _22143_, _22141_);
  and (_22834_, _22833_, _22832_);
  and (_22835_, _22834_, _22831_);
  nor (_22836_, _22129_, _22127_);
  nor (_22837_, _22124_, _22122_);
  and (_22838_, _22837_, _22836_);
  nor (_22839_, _22118_, _22116_);
  nor (_22840_, _22113_, _22111_);
  and (_22841_, _22840_, _22839_);
  and (_22842_, _22841_, _22838_);
  and (_22843_, _22842_, _22835_);
  nor (_22844_, _22196_, _22204_);
  nor (_22845_, _22202_, _22194_);
  and (_22846_, _22845_, _22844_);
  nor (_22847_, _22185_, _22183_);
  nor (_22848_, _22190_, _22188_);
  and (_22849_, _22848_, _22847_);
  and (_22850_, _22849_, _22846_);
  nor (_22851_, _22178_, _22176_);
  nor (_22852_, _22173_, _22171_);
  and (_22853_, _22852_, _22851_);
  nor (_22854_, _22167_, _22165_);
  nor (_22855_, _22162_, _22160_);
  and (_22856_, _22855_, _22854_);
  and (_22857_, _22856_, _22853_);
  and (_22858_, _22857_, _22850_);
  and (_22859_, _22858_, _22843_);
  and (_22860_, _22859_, _22828_);
  nor (_22861_, _22231_, _22229_);
  nor (_22862_, _22225_, _22223_);
  and (_22863_, _22862_, _22861_);
  nor (_22864_, _22214_, _22212_);
  nor (_22865_, _22219_, _22217_);
  and (_22866_, _22865_, _22864_);
  and (_22867_, _22866_, _22863_);
  nor (_22868_, _22249_, _22247_);
  nor (_22869_, _22254_, _22252_);
  and (_22870_, _22869_, _22868_);
  nor (_22871_, _22243_, _22241_);
  nor (_22872_, _22238_, _22236_);
  and (_22873_, _22872_, _22871_);
  and (_22874_, _22873_, _22870_);
  and (_22875_, _22874_, _22867_);
  nor (_22876_, _22296_, _22302_);
  nor (_22877_, _22300_, _22294_);
  and (_22878_, _22877_, _22876_);
  nor (_22879_, _22285_, _22283_);
  nor (_22880_, _22290_, _22288_);
  and (_22881_, _22880_, _22879_);
  and (_22882_, _22881_, _22878_);
  nor (_22883_, _22273_, _22271_);
  nor (_22884_, _22278_, _22276_);
  and (_22885_, _22884_, _22883_);
  nor (_22886_, _22267_, _22265_);
  nor (_22887_, _22262_, _22260_);
  and (_22888_, _22887_, _22886_);
  and (_22889_, _22888_, _22885_);
  and (_22890_, _22889_, _22882_);
  and (_22891_, _22890_, _22875_);
  nor (_22892_, _22335_, _22333_);
  nor (_22893_, _22340_, _22338_);
  and (_22894_, _22893_, _22892_);
  nor (_22895_, _22351_, _22349_);
  nor (_22896_, _22346_, _22344_);
  and (_22897_, _22896_, _22895_);
  and (_22898_, _22897_, _22894_);
  nor (_22899_, _22317_, _22314_);
  nor (_22900_, _22311_, _22309_);
  and (_22901_, _22900_, _22899_);
  nor (_22902_, _22323_, _22321_);
  nor (_22903_, _22328_, _22326_);
  and (_22904_, _22903_, _22902_);
  and (_22905_, _22904_, _22901_);
  and (_22906_, _22905_, _22898_);
  nor (_22907_, _22384_, _22382_);
  nor (_22908_, _22389_, _22387_);
  and (_22909_, _22908_, _22907_);
  nor (_22910_, _22400_, _22398_);
  nor (_22911_, _22395_, _22393_);
  and (_22912_, _22911_, _22910_);
  and (_22913_, _22912_, _22909_);
  nor (_22914_, _22366_, _22362_);
  nor (_22915_, _22359_, _22357_);
  and (_22916_, _22915_, _22914_);
  nor (_22917_, _22372_, _22370_);
  nor (_22918_, _22377_, _22375_);
  and (_22919_, _22918_, _22917_);
  and (_22920_, _22919_, _22916_);
  and (_22921_, _22920_, _22913_);
  and (_22922_, _22921_, _22906_);
  and (_22923_, _22922_, _22891_);
  and (_22924_, _22923_, _22860_);
  nor (_22925_, _22428_, _22420_);
  nor (_22926_, _22422_, _22426_);
  and (_22927_, _22926_, _22925_);
  nor (_22928_, _22416_, _22414_);
  nor (_22929_, _22411_, _22409_);
  and (_22930_, _22929_, _22928_);
  and (_22931_, _22930_, _22927_);
  nor (_22932_, _22440_, _22438_);
  nor (_22933_, _22435_, _22433_);
  and (_22934_, _22933_, _22932_);
  nor (_22935_, _22446_, _22444_);
  nor (_22936_, _22451_, _22449_);
  and (_22937_, _22936_, _22935_);
  and (_22938_, _22937_, _22934_);
  and (_22939_, _22938_, _22931_);
  nor (_22940_, _22493_, _22491_);
  nor (_22941_, _22499_, _22496_);
  and (_22942_, _22941_, _22940_);
  nor (_22943_, _22487_, _22485_);
  nor (_22944_, _22482_, _22480_);
  and (_22945_, _22944_, _22943_);
  and (_22946_, _22945_, _22942_);
  nor (_22947_, _22470_, _22468_);
  nor (_22948_, _22475_, _22473_);
  and (_22949_, _22948_, _22947_);
  nor (_22950_, _22459_, _22457_);
  nor (_22951_, _22464_, _22462_);
  and (_22952_, _22951_, _22950_);
  and (_22953_, _22952_, _22949_);
  and (_22954_, _22953_, _22946_);
  and (_22955_, _22954_, _22939_);
  nor (_22956_, _22519_, _22517_);
  nor (_22957_, _22525_, _22522_);
  and (_22958_, _22957_, _22956_);
  nor (_22959_, _22508_, _22506_);
  nor (_22960_, _22513_, _22511_);
  and (_22961_, _22960_, _22959_);
  and (_22962_, _22961_, _22958_);
  nor (_22963_, _22548_, _22546_);
  nor (_22964_, _22543_, _22541_);
  and (_22965_, _22964_, _22963_);
  nor (_22966_, _22532_, _22530_);
  nor (_22967_, _22537_, _22535_);
  and (_22968_, _22967_, _22966_);
  and (_22969_, _22968_, _22965_);
  and (_22970_, _22969_, _22962_);
  nor (_22971_, _22563_, _22554_);
  nor (_22972_, _22556_, _22561_);
  and (_22973_, _22972_, _22971_);
  nor (_22974_, _22574_, _22572_);
  nor (_22975_, _22569_, _22567_);
  and (_22976_, _22975_, _22974_);
  and (_22977_, _22976_, _22973_);
  nor (_22978_, _22592_, _22590_);
  nor (_22979_, _22597_, _22595_);
  and (_22980_, _22979_, _22978_);
  nor (_22981_, _22581_, _22579_);
  nor (_22982_, _22586_, _22584_);
  and (_22983_, _22982_, _22981_);
  and (_22984_, _22983_, _22980_);
  and (_22985_, _22984_, _22977_);
  and (_22986_, _22985_, _22970_);
  and (_22987_, _22986_, _22955_);
  nor (_22988_, _22644_, _22641_);
  nor (_22989_, _22647_, _22639_);
  and (_22990_, _22989_, _22988_);
  nor (_22991_, _22635_, _22633_);
  nor (_22992_, _22630_, _22628_);
  and (_22993_, _22992_, _22991_);
  and (_22994_, _22993_, _22990_);
  nor (_22995_, _22607_, _22605_);
  nor (_22996_, _22612_, _22610_);
  and (_22997_, _22996_, _22995_);
  nor (_22998_, _22618_, _22616_);
  nor (_22999_, _22623_, _22621_);
  and (_23000_, _22999_, _22998_);
  and (_23001_, _23000_, _22997_);
  and (_23002_, _23001_, _22994_);
  nor (_23003_, _22695_, _22689_);
  nor (_23004_, _22687_, _22693_);
  and (_23005_, _23004_, _23003_);
  nor (_23006_, _22678_, _22676_);
  nor (_23007_, _22683_, _22681_);
  and (_23008_, _23007_, _23006_);
  and (_23009_, _23008_, _23005_);
  nor (_23010_, _22671_, _22669_);
  nor (_23011_, _22666_, _22664_);
  and (_23012_, _23011_, _23010_);
  nor (_23013_, _22655_, _22653_);
  nor (_23014_, _22660_, _22658_);
  and (_23015_, _23014_, _23013_);
  and (_23016_, _23015_, _23012_);
  and (_23017_, _23016_, _23009_);
  and (_23018_, _23017_, _23002_);
  nor (_23019_, _22788_, _22786_);
  nor (_23020_, _22783_, _22781_);
  and (_23021_, _23020_, _23019_);
  nor (_23022_, _22772_, _22770_);
  nor (_23023_, _22777_, _22775_);
  and (_23024_, _23023_, _23022_);
  and (_23025_, _23024_, _23021_);
  nor (_23026_, _22754_, _22752_);
  nor (_23027_, _22749_, _22747_);
  and (_23028_, _23027_, _23026_);
  nor (_23029_, _22765_, _22763_);
  nor (_23030_, _22760_, _22758_);
  and (_23031_, _23030_, _23029_);
  and (_23032_, _23031_, _23028_);
  and (_23033_, _23032_, _23025_);
  nor (_23034_, _22012_, _22015_);
  nor (_23035_, _22019_, _21986_);
  nand (_23036_, _23035_, _23034_);
  nand (_23037_, _23036_, _22702_);
  nor (_23038_, _22725_, _22723_);
  nor (_23039_, _22730_, _22728_);
  and (_23040_, _23039_, _23038_);
  nor (_23041_, _22741_, _22739_);
  nor (_23042_, _22736_, _22734_);
  and (_23043_, _23042_, _23041_);
  and (_23044_, _23043_, _23040_);
  and (_23045_, _23044_, _23037_);
  and (_23046_, _23045_, _23033_);
  and (_23047_, _23046_, _23018_);
  and (_23048_, _23047_, _22987_);
  and (_23049_, _23048_, _22924_);
  and (_23050_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_23051_, _23050_, _22797_);
  and (_23052_, _23051_, _00006_);
  or (_23053_, _23052_, _21944_);
  and (_00003_[6], _23053_, _38997_);
  and (_23054_, _15589_, iram_op1[5]);
  and (_23055_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  and (_23056_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_23057_, _23056_, _23055_);
  and (_23058_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_23059_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_23060_, _23059_, _23058_);
  or (_23061_, _23060_, _23057_);
  and (_23062_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and (_23063_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_23064_, _23063_, _23062_);
  and (_23065_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_23066_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or (_23067_, _23066_, _23065_);
  or (_23068_, _23067_, _23064_);
  or (_23069_, _23068_, _23061_);
  and (_23070_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_23071_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or (_23072_, _23071_, _23070_);
  and (_23073_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  and (_23074_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_23075_, _23074_, _23073_);
  or (_23076_, _23075_, _23072_);
  and (_23077_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_23078_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or (_23079_, _23078_, _23077_);
  and (_23080_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_23081_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_23082_, _23081_, _23080_);
  or (_23083_, _23082_, _23079_);
  or (_23084_, _23083_, _23076_);
  or (_23085_, _23084_, _23069_);
  and (_23086_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_23087_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or (_23088_, _23087_, _23086_);
  and (_23089_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  and (_23090_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_23091_, _23090_, _23089_);
  or (_23092_, _23091_, _23088_);
  and (_23093_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_23094_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_23095_, _23094_, _23093_);
  and (_23096_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  and (_23097_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_23098_, _23097_, _23096_);
  or (_23099_, _23098_, _23095_);
  or (_23100_, _23099_, _23092_);
  and (_23101_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  and (_23102_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or (_23103_, _23102_, _23101_);
  and (_23104_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  and (_23105_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_23106_, _23105_, _23104_);
  or (_23107_, _23106_, _23103_);
  and (_23108_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  and (_23109_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_23110_, _23109_, _23108_);
  and (_23111_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_23112_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_23113_, _23112_, _23111_);
  or (_23114_, _23113_, _23110_);
  or (_23115_, _23114_, _23107_);
  or (_23116_, _23115_, _23100_);
  or (_23117_, _23116_, _23085_);
  and (_23118_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_23119_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or (_23120_, _23119_, _23118_);
  and (_23121_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and (_23122_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_23123_, _23122_, _23121_);
  or (_23124_, _23123_, _23120_);
  and (_23125_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_23126_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or (_23127_, _23126_, _23125_);
  and (_23128_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_23129_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_23130_, _23129_, _23128_);
  or (_23131_, _23130_, _23127_);
  or (_23132_, _23131_, _23124_);
  and (_23133_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_23134_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or (_23135_, _23134_, _23133_);
  and (_23136_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and (_23137_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_23138_, _23137_, _23136_);
  or (_23139_, _23138_, _23135_);
  and (_23140_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and (_23141_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_23142_, _23141_, _23140_);
  and (_23143_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_23144_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_23145_, _23144_, _23143_);
  or (_23146_, _23145_, _23142_);
  or (_23147_, _23146_, _23139_);
  or (_23148_, _23147_, _23132_);
  and (_23149_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  and (_23150_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_23151_, _23150_, _23149_);
  and (_23152_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_23153_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_23154_, _23153_, _23152_);
  or (_23155_, _23154_, _23151_);
  and (_23156_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and (_23157_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_23158_, _23157_, _23156_);
  and (_23159_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_23160_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_23161_, _23160_, _23159_);
  or (_23162_, _23161_, _23158_);
  or (_23163_, _23162_, _23155_);
  and (_23164_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_23165_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_23166_, _23165_, _23164_);
  and (_23167_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  and (_23168_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_23169_, _23168_, _23167_);
  or (_23170_, _23169_, _23166_);
  and (_23171_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_23172_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_23173_, _23172_, _23171_);
  and (_23174_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  and (_23175_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_23176_, _23175_, _23174_);
  or (_23177_, _23176_, _23173_);
  or (_23178_, _23177_, _23170_);
  or (_23179_, _23178_, _23163_);
  or (_23180_, _23179_, _23148_);
  or (_23181_, _23180_, _23117_);
  and (_23182_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_23183_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_23184_, _23183_, _23182_);
  and (_23185_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  and (_23186_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_23187_, _23186_, _23185_);
  or (_23188_, _23187_, _23184_);
  and (_23189_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_23190_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or (_23191_, _23190_, _23189_);
  and (_23192_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_23193_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_23194_, _23193_, _23192_);
  or (_23195_, _23194_, _23191_);
  or (_23196_, _23195_, _23188_);
  and (_23197_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  and (_23198_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_23199_, _23198_, _23197_);
  and (_23200_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_23201_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or (_23202_, _23201_, _23200_);
  or (_23203_, _23202_, _23199_);
  and (_23204_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_23205_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_23206_, _23205_, _23204_);
  and (_23207_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  and (_23208_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_23209_, _23208_, _23207_);
  or (_23210_, _23209_, _23206_);
  or (_23211_, _23210_, _23203_);
  or (_23212_, _23211_, _23196_);
  and (_23213_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_23214_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_23215_, _23214_, _23213_);
  and (_23216_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_23217_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  or (_23218_, _23217_, _23216_);
  or (_23219_, _23218_, _23215_);
  and (_23220_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_23221_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_23222_, _23221_, _23220_);
  and (_23223_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_23224_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_23225_, _23224_, _23223_);
  or (_23226_, _23225_, _23222_);
  or (_23227_, _23226_, _23219_);
  and (_23228_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_23229_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  or (_23230_, _23229_, _23228_);
  and (_23231_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_23232_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_23233_, _23232_, _23231_);
  or (_23234_, _23233_, _23230_);
  and (_23235_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_23236_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  or (_23237_, _23236_, _23235_);
  and (_23238_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  and (_23239_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_23240_, _23239_, _23238_);
  or (_23241_, _23240_, _23237_);
  or (_23242_, _23241_, _23234_);
  or (_23243_, _23242_, _23227_);
  or (_23244_, _23243_, _23212_);
  and (_23245_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and (_23246_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_23247_, _23246_, _23245_);
  and (_23248_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_23249_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or (_23250_, _23249_, _23248_);
  or (_23251_, _23250_, _23247_);
  and (_23252_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_23253_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or (_23254_, _23253_, _23252_);
  and (_23255_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and (_23256_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_23257_, _23256_, _23255_);
  or (_23258_, _23257_, _23254_);
  or (_23259_, _23258_, _23251_);
  and (_23260_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_23261_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or (_23262_, _23261_, _23260_);
  and (_23263_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  and (_23264_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_23265_, _23264_, _23263_);
  or (_23266_, _23265_, _23262_);
  and (_23267_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_23268_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or (_23269_, _23268_, _23267_);
  and (_23270_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_23271_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_23272_, _23271_, _23270_);
  or (_23273_, _23272_, _23269_);
  or (_23274_, _23273_, _23266_);
  or (_23275_, _23274_, _23259_);
  and (_23276_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  and (_23277_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_23278_, _23277_, _23276_);
  and (_23279_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and (_23280_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or (_23281_, _23280_, _23279_);
  or (_23282_, _23281_, _23278_);
  and (_23283_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_23284_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or (_23285_, _23284_, _23283_);
  and (_23286_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and (_23287_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_23288_, _23287_, _23286_);
  or (_23289_, _23288_, _23285_);
  or (_23290_, _23289_, _23282_);
  and (_23291_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_23292_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or (_23293_, _23292_, _23291_);
  and (_23294_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and (_23295_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_23296_, _23295_, _23294_);
  or (_23297_, _23296_, _23293_);
  and (_23298_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_23299_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or (_23300_, _23299_, _23298_);
  and (_23301_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and (_23302_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_23303_, _23302_, _23301_);
  or (_23304_, _23303_, _23300_);
  or (_23305_, _23304_, _23297_);
  or (_23306_, _23305_, _23290_);
  or (_23307_, _23306_, _23275_);
  or (_23308_, _23307_, _23244_);
  or (_23309_, _23308_, _23181_);
  and (_23310_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  and (_23311_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_23312_, _23311_, _23310_);
  and (_23313_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_23314_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or (_23315_, _23314_, _23313_);
  or (_23316_, _23315_, _23312_);
  and (_23317_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  and (_23318_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_23319_, _23318_, _23317_);
  and (_23320_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_23321_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_23322_, _23321_, _23320_);
  or (_23323_, _23322_, _23319_);
  or (_23324_, _23323_, _23316_);
  and (_23325_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_23326_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or (_23327_, _23326_, _23325_);
  and (_23328_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_23329_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_23330_, _23329_, _23328_);
  or (_23331_, _23330_, _23327_);
  and (_23332_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_23333_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_23334_, _23333_, _23332_);
  and (_23335_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  and (_23336_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_23337_, _23336_, _23335_);
  or (_23338_, _23337_, _23334_);
  or (_23339_, _23338_, _23331_);
  or (_23340_, _23339_, _23324_);
  and (_23341_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  and (_23342_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_23343_, _23342_, _23341_);
  and (_23344_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_23345_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_23346_, _23345_, _23344_);
  or (_23347_, _23346_, _23343_);
  and (_23348_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  and (_23349_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_23350_, _23349_, _23348_);
  and (_23351_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_23352_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_23353_, _23352_, _23351_);
  or (_23354_, _23353_, _23350_);
  or (_23355_, _23354_, _23347_);
  and (_23356_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_23357_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_23358_, _23357_, _23356_);
  and (_23359_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  and (_23360_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_23361_, _23360_, _23359_);
  or (_23362_, _23361_, _23358_);
  and (_23363_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_23364_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_23365_, _23364_, _23363_);
  and (_23366_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  and (_23367_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_23368_, _23367_, _23366_);
  or (_23369_, _23368_, _23365_);
  or (_23370_, _23369_, _23362_);
  or (_23371_, _23370_, _23355_);
  or (_23372_, _23371_, _23340_);
  and (_23373_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  and (_23374_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_23375_, _23374_, _23373_);
  and (_23376_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_23377_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_23378_, _23377_, _23376_);
  or (_23379_, _23378_, _23375_);
  and (_23380_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  and (_23381_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_23382_, _23381_, _23380_);
  and (_23383_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_23384_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_23385_, _23384_, _23383_);
  or (_23386_, _23385_, _23382_);
  or (_23387_, _23386_, _23379_);
  and (_23388_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_23389_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_23390_, _23389_, _23388_);
  and (_23391_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  and (_23392_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_23393_, _23392_, _23391_);
  or (_23394_, _23393_, _23390_);
  and (_23395_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_23396_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_23397_, _23396_, _23395_);
  and (_23398_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  and (_23399_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_23400_, _23399_, _23398_);
  or (_23401_, _23400_, _23397_);
  or (_23402_, _23401_, _23394_);
  or (_23403_, _23402_, _23387_);
  and (_23404_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and (_23405_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_23406_, _23405_, _23404_);
  and (_23407_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_23408_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_23409_, _23408_, _23407_);
  or (_23410_, _23409_, _23406_);
  and (_23411_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and (_23412_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_23413_, _23412_, _23411_);
  and (_23414_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  and (_23415_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_23416_, _23415_, _23414_);
  or (_23417_, _23416_, _23413_);
  or (_23418_, _23417_, _23410_);
  and (_23419_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_23420_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_23421_, _23420_, _23419_);
  and (_23422_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  and (_23423_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_23424_, _23423_, _23422_);
  or (_23425_, _23424_, _23421_);
  and (_23426_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_23427_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_23428_, _23427_, _23426_);
  and (_23429_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  and (_23430_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_23431_, _23430_, _23429_);
  or (_23432_, _23431_, _23428_);
  or (_23433_, _23432_, _23425_);
  or (_23434_, _23433_, _23418_);
  or (_23435_, _23434_, _23403_);
  or (_23436_, _23435_, _23372_);
  and (_23437_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  and (_23438_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_23439_, _23438_, _23437_);
  and (_23440_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_23441_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_23442_, _23441_, _23440_);
  or (_23443_, _23442_, _23439_);
  and (_23444_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  and (_23445_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_23446_, _23445_, _23444_);
  and (_23447_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_23448_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_23449_, _23448_, _23447_);
  or (_23450_, _23449_, _23446_);
  or (_23451_, _23450_, _23443_);
  and (_23452_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_23453_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_23454_, _23453_, _23452_);
  and (_23455_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  and (_23456_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_23457_, _23456_, _23455_);
  or (_23458_, _23457_, _23454_);
  and (_23459_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_23460_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_23461_, _23460_, _23459_);
  and (_23462_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  and (_23463_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_23464_, _23463_, _23462_);
  or (_23465_, _23464_, _23461_);
  or (_23466_, _23465_, _23458_);
  or (_23467_, _23466_, _23451_);
  and (_23468_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_23469_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_23470_, _23469_, _23468_);
  and (_23471_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  and (_23472_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_23473_, _23472_, _23471_);
  or (_23474_, _23473_, _23470_);
  and (_23475_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_23476_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_23477_, _23476_, _23475_);
  and (_23478_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  and (_23479_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_23480_, _23479_, _23478_);
  or (_23481_, _23480_, _23477_);
  or (_23482_, _23481_, _23474_);
  and (_23483_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  and (_23484_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_23485_, _23484_, _23483_);
  and (_23486_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_23487_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_23488_, _23487_, _23486_);
  or (_23489_, _23488_, _23485_);
  and (_23490_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  and (_23491_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_23492_, _23491_, _23490_);
  and (_23493_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  and (_23494_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_23495_, _23494_, _23493_);
  or (_23496_, _23495_, _23492_);
  or (_23497_, _23496_, _23489_);
  or (_23498_, _23497_, _23482_);
  or (_23499_, _23498_, _23467_);
  and (_23500_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_23501_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_23502_, _23501_, _23500_);
  and (_23503_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  and (_23504_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_23505_, _23504_, _23503_);
  or (_23506_, _23505_, _23502_);
  and (_23507_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_23508_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_23509_, _23508_, _23507_);
  and (_23510_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  and (_23511_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_23512_, _23511_, _23510_);
  or (_23513_, _23512_, _23509_);
  or (_23514_, _23513_, _23506_);
  and (_23515_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  and (_23516_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_23517_, _23516_, _23515_);
  and (_23518_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_23519_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_23520_, _23519_, _23518_);
  or (_23521_, _23520_, _23517_);
  and (_23522_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  and (_23523_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_23524_, _23523_, _23522_);
  and (_23525_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_23526_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_23527_, _23526_, _23525_);
  or (_23528_, _23527_, _23524_);
  or (_23529_, _23528_, _23521_);
  or (_23530_, _23529_, _23514_);
  and (_23531_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_23532_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_23533_, _23532_, _23531_);
  and (_23534_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_23535_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_23536_, _23535_, _23534_);
  or (_23537_, _23536_, _23533_);
  and (_23538_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_23539_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_23540_, _23539_, _23538_);
  and (_23541_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_23542_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_23543_, _23542_, _23541_);
  or (_23544_, _23543_, _23540_);
  or (_23545_, _23544_, _23537_);
  and (_23546_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_23547_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_23548_, _23547_, _23546_);
  and (_23549_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_23550_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_23551_, _23550_, _23549_);
  or (_23552_, _23551_, _23548_);
  and (_23553_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_23554_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_23555_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_23556_, _23555_, _23554_);
  or (_23557_, _23556_, _23553_);
  or (_23558_, _23557_, _23552_);
  or (_23559_, _23558_, _23545_);
  or (_23560_, _23559_, _23530_);
  or (_23561_, _23560_, _23499_);
  or (_23562_, _23561_, _23436_);
  or (_23563_, _23562_, _23309_);
  and (_23564_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_23565_, _23564_, _23563_);
  and (_23566_, _23565_, _00006_);
  or (_23567_, _23566_, _23054_);
  and (_00003_[5], _23567_, _38997_);
  and (_23568_, _15589_, iram_op1[4]);
  and (_23569_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and (_23570_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_23571_, _23570_, _23569_);
  and (_23572_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_23573_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or (_23574_, _23573_, _23572_);
  or (_23575_, _23574_, _23571_);
  and (_23576_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and (_23577_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_23578_, _23577_, _23576_);
  and (_23579_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_23580_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or (_23581_, _23580_, _23579_);
  or (_23582_, _23581_, _23578_);
  or (_23583_, _23582_, _23575_);
  and (_23584_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_23585_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or (_23586_, _23585_, _23584_);
  and (_23587_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and (_23588_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_23589_, _23588_, _23587_);
  or (_23590_, _23589_, _23586_);
  and (_23591_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_23592_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or (_23593_, _23592_, _23591_);
  and (_23594_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  and (_23595_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or (_23596_, _23595_, _23594_);
  or (_23597_, _23596_, _23593_);
  or (_23598_, _23597_, _23590_);
  or (_23599_, _23598_, _23583_);
  and (_23600_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  and (_23601_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_23602_, _23601_, _23600_);
  and (_23603_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_23604_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or (_23605_, _23604_, _23603_);
  or (_23606_, _23605_, _23602_);
  and (_23607_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  and (_23608_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_23609_, _23608_, _23607_);
  and (_23610_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_23611_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_23612_, _23611_, _23610_);
  or (_23613_, _23612_, _23609_);
  or (_23614_, _23613_, _23606_);
  and (_23615_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_23616_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or (_23617_, _23616_, _23615_);
  and (_23618_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  and (_23619_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_23620_, _23619_, _23618_);
  or (_23621_, _23620_, _23617_);
  and (_23622_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_23623_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or (_23624_, _23623_, _23622_);
  and (_23625_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  and (_23626_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_23627_, _23626_, _23625_);
  or (_23628_, _23627_, _23624_);
  or (_23629_, _23628_, _23621_);
  or (_23630_, _23629_, _23614_);
  or (_23631_, _23630_, _23599_);
  and (_23632_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_23633_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or (_23634_, _23633_, _23632_);
  and (_23635_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  and (_23636_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_23637_, _23636_, _23635_);
  or (_23638_, _23637_, _23634_);
  and (_23639_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_23640_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or (_23641_, _23640_, _23639_);
  and (_23642_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  and (_23643_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_23644_, _23643_, _23642_);
  or (_23645_, _23644_, _23641_);
  or (_23646_, _23645_, _23638_);
  and (_23647_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  and (_23648_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_23649_, _23648_, _23647_);
  and (_23650_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  and (_23651_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or (_23652_, _23651_, _23650_);
  or (_23653_, _23652_, _23649_);
  and (_23654_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_23655_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or (_23656_, _23655_, _23654_);
  and (_23657_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  and (_23658_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_23659_, _23658_, _23657_);
  or (_23660_, _23659_, _23656_);
  or (_23661_, _23660_, _23653_);
  or (_23662_, _23661_, _23646_);
  and (_23663_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_23664_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  or (_23665_, _23664_, _23663_);
  and (_23666_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and (_23667_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_23668_, _23667_, _23666_);
  or (_23669_, _23668_, _23665_);
  and (_23670_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_23671_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  or (_23672_, _23671_, _23670_);
  and (_23673_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and (_23674_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  or (_23675_, _23674_, _23673_);
  or (_23676_, _23675_, _23672_);
  or (_23677_, _23676_, _23669_);
  and (_23678_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and (_23679_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_23680_, _23679_, _23678_);
  and (_23681_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_23682_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  or (_23683_, _23682_, _23681_);
  or (_23684_, _23683_, _23680_);
  and (_23685_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and (_23686_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_23687_, _23686_, _23685_);
  and (_23688_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_23689_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  or (_23690_, _23689_, _23688_);
  or (_23691_, _23690_, _23687_);
  or (_23692_, _23691_, _23684_);
  or (_23693_, _23692_, _23677_);
  or (_23694_, _23693_, _23662_);
  or (_23695_, _23694_, _23631_);
  and (_23696_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_23697_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or (_23698_, _23697_, _23696_);
  and (_23699_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  and (_23700_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_23701_, _23700_, _23699_);
  or (_23702_, _23701_, _23698_);
  and (_23703_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_23704_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or (_23705_, _23704_, _23703_);
  and (_23706_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  and (_23707_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or (_23708_, _23707_, _23706_);
  or (_23709_, _23708_, _23705_);
  or (_23710_, _23709_, _23702_);
  and (_23711_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  and (_23712_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_23713_, _23712_, _23711_);
  and (_23714_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_23715_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or (_23716_, _23715_, _23714_);
  or (_23717_, _23716_, _23713_);
  and (_23718_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  and (_23719_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_23720_, _23719_, _23718_);
  and (_23721_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_23722_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or (_23723_, _23722_, _23721_);
  or (_23724_, _23723_, _23720_);
  or (_23725_, _23724_, _23717_);
  or (_23726_, _23725_, _23710_);
  and (_23727_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and (_23728_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_23729_, _23728_, _23727_);
  and (_23730_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_23731_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  or (_23732_, _23731_, _23730_);
  or (_23733_, _23732_, _23729_);
  and (_23734_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_23735_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_23736_, _23735_, _23734_);
  and (_23737_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_23738_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  or (_23739_, _23738_, _23737_);
  or (_23740_, _23739_, _23736_);
  or (_23741_, _23740_, _23733_);
  and (_23742_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_23743_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_23744_, _23743_, _23742_);
  and (_23745_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_23746_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  or (_23747_, _23746_, _23745_);
  or (_23748_, _23747_, _23744_);
  and (_23749_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_23750_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  or (_23751_, _23750_, _23749_);
  and (_23752_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and (_23753_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_23754_, _23753_, _23752_);
  or (_23755_, _23754_, _23751_);
  or (_23756_, _23755_, _23748_);
  or (_23757_, _23756_, _23741_);
  or (_23758_, _23757_, _23726_);
  and (_23759_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and (_23760_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_23761_, _23760_, _23759_);
  and (_23762_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_23763_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or (_23764_, _23763_, _23762_);
  or (_23765_, _23764_, _23761_);
  and (_23766_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and (_23767_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_23768_, _23767_, _23766_);
  and (_23769_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_23770_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or (_23771_, _23770_, _23769_);
  or (_23772_, _23771_, _23768_);
  or (_23773_, _23772_, _23765_);
  and (_23774_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_23775_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or (_23776_, _23775_, _23774_);
  and (_23777_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  and (_23778_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_23779_, _23778_, _23777_);
  or (_23780_, _23779_, _23776_);
  and (_23781_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_23782_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or (_23783_, _23782_, _23781_);
  and (_23784_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_23785_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_23786_, _23785_, _23784_);
  or (_23787_, _23786_, _23783_);
  or (_23788_, _23787_, _23780_);
  or (_23789_, _23788_, _23773_);
  and (_23790_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  and (_23791_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_23792_, _23791_, _23790_);
  and (_23793_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and (_23794_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or (_23795_, _23794_, _23793_);
  or (_23796_, _23795_, _23792_);
  and (_23797_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and (_23798_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_23799_, _23798_, _23797_);
  and (_23800_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_23801_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or (_23802_, _23801_, _23800_);
  or (_23803_, _23802_, _23799_);
  or (_23804_, _23803_, _23796_);
  and (_23805_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_23806_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or (_23807_, _23806_, _23805_);
  and (_23808_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  and (_23809_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_23810_, _23809_, _23808_);
  or (_23811_, _23810_, _23807_);
  and (_23812_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_23813_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or (_23814_, _23813_, _23812_);
  and (_23815_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  and (_23816_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_23817_, _23816_, _23815_);
  or (_23818_, _23817_, _23814_);
  or (_23819_, _23818_, _23811_);
  or (_23820_, _23819_, _23804_);
  or (_23821_, _23820_, _23789_);
  or (_23822_, _23821_, _23758_);
  or (_23823_, _23822_, _23695_);
  and (_23824_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  and (_23825_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_23826_, _23825_, _23824_);
  and (_23827_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_23828_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or (_23829_, _23828_, _23827_);
  or (_23830_, _23829_, _23826_);
  and (_23831_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  and (_23832_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_23833_, _23832_, _23831_);
  and (_23834_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_23835_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or (_23836_, _23835_, _23834_);
  or (_23837_, _23836_, _23833_);
  or (_23838_, _23837_, _23830_);
  and (_23839_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_23840_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or (_23841_, _23840_, _23839_);
  and (_23842_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_23843_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_23844_, _23843_, _23842_);
  or (_23845_, _23844_, _23841_);
  and (_23846_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_23847_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or (_23848_, _23847_, _23846_);
  and (_23849_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  and (_23850_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_23851_, _23850_, _23849_);
  or (_23852_, _23851_, _23848_);
  or (_23853_, _23852_, _23845_);
  or (_23854_, _23853_, _23838_);
  and (_23855_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  and (_23856_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_23857_, _23856_, _23855_);
  and (_23858_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_23859_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_23860_, _23859_, _23858_);
  or (_23861_, _23860_, _23857_);
  and (_23862_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  and (_23863_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_23864_, _23863_, _23862_);
  and (_23865_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_23866_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_23867_, _23866_, _23865_);
  or (_23868_, _23867_, _23864_);
  or (_23869_, _23868_, _23861_);
  and (_23870_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_23871_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_23872_, _23871_, _23870_);
  and (_23873_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  and (_23874_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_23875_, _23874_, _23873_);
  or (_23876_, _23875_, _23872_);
  and (_23877_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_23878_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_23879_, _23878_, _23877_);
  and (_23880_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  and (_23881_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_23882_, _23881_, _23880_);
  or (_23883_, _23882_, _23879_);
  or (_23884_, _23883_, _23876_);
  or (_23885_, _23884_, _23869_);
  or (_23886_, _23885_, _23854_);
  and (_23887_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_23888_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_23889_, _23888_, _23887_);
  and (_23890_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_23891_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_23892_, _23891_, _23890_);
  or (_23893_, _23892_, _23889_);
  and (_23894_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_23895_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_23896_, _23895_, _23894_);
  and (_23897_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  and (_23898_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_23899_, _23898_, _23897_);
  or (_23900_, _23899_, _23896_);
  or (_23901_, _23900_, _23893_);
  and (_23902_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  and (_23903_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_23904_, _23903_, _23902_);
  and (_23905_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_23906_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_23907_, _23906_, _23905_);
  or (_23908_, _23907_, _23904_);
  and (_23909_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  and (_23910_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_23911_, _23910_, _23909_);
  and (_23912_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_23913_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_23914_, _23913_, _23912_);
  or (_23915_, _23914_, _23911_);
  or (_23916_, _23915_, _23908_);
  or (_23917_, _23916_, _23901_);
  and (_23918_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_23919_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_23920_, _23919_, _23918_);
  and (_23921_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  and (_23922_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_23923_, _23922_, _23921_);
  or (_23924_, _23923_, _23920_);
  and (_23925_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  and (_23926_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_23927_, _23926_, _23925_);
  and (_23928_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_23929_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_23930_, _23929_, _23928_);
  or (_23931_, _23930_, _23927_);
  or (_23932_, _23931_, _23924_);
  and (_23933_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and (_23934_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_23935_, _23934_, _23933_);
  and (_23936_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and (_23937_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_23938_, _23937_, _23936_);
  or (_23939_, _23938_, _23935_);
  and (_23940_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and (_23941_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_23942_, _23941_, _23940_);
  and (_23943_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_23944_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_23945_, _23944_, _23943_);
  or (_23946_, _23945_, _23942_);
  or (_23947_, _23946_, _23939_);
  or (_23948_, _23947_, _23932_);
  or (_23949_, _23948_, _23917_);
  or (_23950_, _23949_, _23886_);
  and (_23951_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  and (_23952_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_23953_, _23952_, _23951_);
  and (_23954_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_23955_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_23956_, _23955_, _23954_);
  or (_23957_, _23956_, _23953_);
  and (_23958_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  and (_23959_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_23960_, _23959_, _23958_);
  and (_23961_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_23962_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_23963_, _23962_, _23961_);
  or (_23964_, _23963_, _23960_);
  or (_23965_, _23964_, _23957_);
  and (_23966_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_23967_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_23968_, _23967_, _23966_);
  and (_23969_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  and (_23970_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_23971_, _23970_, _23969_);
  or (_23972_, _23971_, _23968_);
  and (_23973_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_23974_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_23975_, _23974_, _23973_);
  and (_23976_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  and (_23977_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_23978_, _23977_, _23976_);
  or (_23979_, _23978_, _23975_);
  or (_23980_, _23979_, _23972_);
  or (_23981_, _23980_, _23965_);
  and (_23982_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_23983_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_23984_, _23983_, _23982_);
  and (_23985_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  and (_23986_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_23987_, _23986_, _23985_);
  or (_23988_, _23987_, _23984_);
  and (_23989_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_23990_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_23991_, _23990_, _23989_);
  and (_23992_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  and (_23993_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_23994_, _23993_, _23992_);
  or (_23995_, _23994_, _23991_);
  or (_23996_, _23995_, _23988_);
  and (_23997_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_23998_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_23999_, _23998_, _23997_);
  and (_24000_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  and (_24001_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_24002_, _24001_, _24000_);
  or (_24003_, _24002_, _23999_);
  and (_24004_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_24005_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or (_24006_, _24005_, _24004_);
  and (_24007_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  and (_24008_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_24009_, _24008_, _24007_);
  or (_24010_, _24009_, _24006_);
  or (_24011_, _24010_, _24003_);
  or (_24012_, _24011_, _23996_);
  or (_24013_, _24012_, _23981_);
  and (_24014_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_24015_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_24016_, _24015_, _24014_);
  and (_24017_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  and (_24018_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_24019_, _24018_, _24017_);
  or (_24020_, _24019_, _24016_);
  and (_24021_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_24022_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_24023_, _24022_, _24021_);
  and (_24024_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_24025_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_24026_, _24025_, _24024_);
  or (_24027_, _24026_, _24023_);
  or (_24028_, _24027_, _24020_);
  and (_24029_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  and (_24030_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_24031_, _24030_, _24029_);
  and (_24032_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_24033_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_24034_, _24033_, _24032_);
  or (_24035_, _24034_, _24031_);
  and (_24036_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  and (_24037_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_24038_, _24037_, _24036_);
  and (_24039_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_24040_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_24041_, _24040_, _24039_);
  or (_24042_, _24041_, _24038_);
  or (_24043_, _24042_, _24035_);
  or (_24044_, _24043_, _24028_);
  and (_24045_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_24046_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_24047_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_24048_, _24047_, _24046_);
  or (_24049_, _24048_, _24045_);
  and (_24050_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_24051_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_24052_, _24051_, _24050_);
  and (_24053_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_24054_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_24055_, _24054_, _24053_);
  or (_24056_, _24055_, _24052_);
  or (_24057_, _24056_, _24049_);
  and (_24058_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_24059_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_24060_, _24059_, _24058_);
  and (_24061_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_24062_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_24063_, _24062_, _24061_);
  or (_24064_, _24063_, _24060_);
  and (_24065_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_24066_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_24067_, _24066_, _24065_);
  and (_24068_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_24069_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_24070_, _24069_, _24068_);
  or (_24071_, _24070_, _24067_);
  or (_24072_, _24071_, _24064_);
  or (_24073_, _24072_, _24057_);
  or (_24074_, _24073_, _24044_);
  or (_24075_, _24074_, _24013_);
  or (_24076_, _24075_, _23950_);
  or (_24077_, _24076_, _23823_);
  and (_24078_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_24079_, _24078_, _24077_);
  and (_24080_, _24079_, _00006_);
  or (_24081_, _24080_, _23568_);
  and (_00003_[4], _24081_, _38997_);
  and (_24082_, _15589_, iram_op1[3]);
  and (_24083_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_24084_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or (_24085_, _24084_, _24083_);
  and (_24086_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and (_24087_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_24088_, _24087_, _24086_);
  or (_24089_, _24088_, _24085_);
  and (_24090_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_24091_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or (_24092_, _24091_, _24090_);
  and (_24093_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_24094_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_24095_, _24094_, _24093_);
  or (_24096_, _24095_, _24092_);
  or (_24097_, _24096_, _24089_);
  and (_24098_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and (_24099_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_24100_, _24099_, _24098_);
  and (_24101_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_24102_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or (_24103_, _24102_, _24101_);
  or (_24104_, _24103_, _24100_);
  and (_24105_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  and (_24106_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_24107_, _24106_, _24105_);
  and (_24108_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_24109_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or (_24110_, _24109_, _24108_);
  or (_24111_, _24110_, _24107_);
  or (_24112_, _24111_, _24104_);
  or (_24113_, _24112_, _24097_);
  and (_24114_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  and (_24115_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_24116_, _24115_, _24114_);
  and (_24117_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  and (_24118_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or (_24119_, _24118_, _24117_);
  or (_24120_, _24119_, _24116_);
  and (_24121_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  and (_24122_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_24123_, _24122_, _24121_);
  and (_24124_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_24125_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or (_24126_, _24125_, _24124_);
  or (_24127_, _24126_, _24123_);
  or (_24128_, _24127_, _24120_);
  and (_24129_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_24130_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or (_24131_, _24130_, _24129_);
  and (_24132_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  and (_24133_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_24134_, _24133_, _24132_);
  or (_24135_, _24134_, _24131_);
  and (_24136_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_24137_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or (_24138_, _24137_, _24136_);
  and (_24139_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  and (_24140_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_24141_, _24140_, _24139_);
  or (_24142_, _24141_, _24138_);
  or (_24143_, _24142_, _24135_);
  or (_24144_, _24143_, _24128_);
  or (_24145_, _24144_, _24113_);
  and (_24146_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_24147_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  or (_24148_, _24147_, _24146_);
  and (_24149_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and (_24150_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_24151_, _24150_, _24149_);
  or (_24152_, _24151_, _24148_);
  and (_24153_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_24154_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  or (_24155_, _24154_, _24153_);
  and (_24156_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and (_24157_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  or (_24158_, _24157_, _24156_);
  or (_24159_, _24158_, _24155_);
  or (_24160_, _24159_, _24152_);
  and (_24161_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_24162_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  or (_24163_, _24162_, _24161_);
  and (_24164_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and (_24165_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_24166_, _24165_, _24164_);
  or (_24167_, _24166_, _24163_);
  and (_24168_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and (_24169_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_24170_, _24169_, _24168_);
  and (_24171_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_24172_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  or (_24173_, _24172_, _24171_);
  or (_24174_, _24173_, _24170_);
  or (_24175_, _24174_, _24167_);
  or (_24176_, _24175_, _24160_);
  and (_24177_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_24178_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or (_24179_, _24178_, _24177_);
  and (_24180_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  and (_24181_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_24182_, _24181_, _24180_);
  or (_24183_, _24182_, _24179_);
  and (_24184_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_24185_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or (_24186_, _24185_, _24184_);
  and (_24187_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  and (_24188_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_24189_, _24188_, _24187_);
  or (_24190_, _24189_, _24186_);
  or (_24191_, _24190_, _24183_);
  and (_24192_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  and (_24193_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_24194_, _24193_, _24192_);
  and (_24195_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_24196_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_24197_, _24196_, _24195_);
  or (_24198_, _24197_, _24194_);
  and (_24199_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and (_24200_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_24201_, _24200_, _24199_);
  and (_24202_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_24203_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or (_24204_, _24203_, _24202_);
  or (_24205_, _24204_, _24201_);
  or (_24206_, _24205_, _24198_);
  or (_24207_, _24206_, _24191_);
  or (_24208_, _24207_, _24176_);
  or (_24209_, _24208_, _24145_);
  and (_24210_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_24211_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or (_24212_, _24211_, _24210_);
  and (_24213_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  and (_24214_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_24215_, _24214_, _24213_);
  or (_24216_, _24215_, _24212_);
  and (_24217_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_24218_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or (_24219_, _24218_, _24217_);
  and (_24220_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_24221_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_24222_, _24221_, _24220_);
  or (_24223_, _24222_, _24219_);
  or (_24224_, _24223_, _24216_);
  and (_24225_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  and (_24226_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_24227_, _24226_, _24225_);
  and (_24228_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_24229_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or (_24230_, _24229_, _24228_);
  or (_24231_, _24230_, _24227_);
  and (_24232_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_24233_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  or (_24234_, _24233_, _24232_);
  and (_24235_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  and (_24236_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_24237_, _24236_, _24235_);
  or (_24238_, _24237_, _24234_);
  or (_24239_, _24238_, _24231_);
  or (_24240_, _24239_, _24224_);
  and (_24241_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and (_24242_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_24243_, _24242_, _24241_);
  and (_24244_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_24245_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  or (_24246_, _24245_, _24244_);
  or (_24247_, _24246_, _24243_);
  and (_24248_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and (_24249_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_24250_, _24249_, _24248_);
  and (_24251_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_24252_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_24253_, _24252_, _24251_);
  or (_24254_, _24253_, _24250_);
  or (_24255_, _24254_, _24247_);
  and (_24256_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_24257_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  or (_24258_, _24257_, _24256_);
  and (_24259_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  and (_24260_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_24261_, _24260_, _24259_);
  or (_24262_, _24261_, _24258_);
  and (_24263_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_24264_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  or (_24265_, _24264_, _24263_);
  and (_24266_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and (_24267_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_24268_, _24267_, _24266_);
  or (_24269_, _24268_, _24265_);
  or (_24270_, _24269_, _24262_);
  or (_24271_, _24270_, _24255_);
  or (_24272_, _24271_, _24240_);
  and (_24273_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_24274_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_24275_, _24274_, _24273_);
  and (_24276_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_24277_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or (_24278_, _24277_, _24276_);
  or (_24279_, _24278_, _24275_);
  and (_24280_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_24281_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or (_24282_, _24281_, _24280_);
  and (_24283_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  and (_24284_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_24285_, _24284_, _24283_);
  or (_24286_, _24285_, _24282_);
  or (_24287_, _24286_, _24279_);
  and (_24288_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and (_24289_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_24290_, _24289_, _24288_);
  and (_24291_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_24292_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or (_24293_, _24292_, _24291_);
  or (_24294_, _24293_, _24290_);
  and (_24295_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  and (_24296_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_24297_, _24296_, _24295_);
  and (_24298_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_24299_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or (_24300_, _24299_, _24298_);
  or (_24301_, _24300_, _24297_);
  or (_24302_, _24301_, _24294_);
  or (_24303_, _24302_, _24287_);
  and (_24304_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and (_24305_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_24306_, _24305_, _24304_);
  and (_24307_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_24308_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_24309_, _24308_, _24307_);
  or (_24310_, _24309_, _24306_);
  and (_24311_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and (_24312_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_24313_, _24312_, _24311_);
  and (_24314_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_24315_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or (_24316_, _24315_, _24314_);
  or (_24317_, _24316_, _24313_);
  or (_24318_, _24317_, _24310_);
  and (_24319_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_24320_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or (_24321_, _24320_, _24319_);
  and (_24322_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  and (_24323_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_24324_, _24323_, _24322_);
  or (_24325_, _24324_, _24321_);
  and (_24326_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_24327_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or (_24328_, _24327_, _24326_);
  and (_24329_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  and (_24330_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_24331_, _24330_, _24329_);
  or (_24332_, _24331_, _24328_);
  or (_24333_, _24332_, _24325_);
  or (_24334_, _24333_, _24318_);
  or (_24335_, _24334_, _24303_);
  or (_24336_, _24335_, _24272_);
  or (_24337_, _24336_, _24209_);
  and (_24338_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  and (_24339_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_24340_, _24339_, _24338_);
  and (_24341_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_24342_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or (_24343_, _24342_, _24341_);
  or (_24344_, _24343_, _24340_);
  and (_24345_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  and (_24346_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_24347_, _24346_, _24345_);
  and (_24348_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_24349_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_24350_, _24349_, _24348_);
  or (_24351_, _24350_, _24347_);
  or (_24352_, _24351_, _24344_);
  and (_24353_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_24354_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or (_24355_, _24354_, _24353_);
  and (_24356_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_24357_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_24358_, _24357_, _24356_);
  or (_24359_, _24358_, _24355_);
  and (_24360_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_24361_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or (_24362_, _24361_, _24360_);
  and (_24363_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  and (_24364_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_24365_, _24364_, _24363_);
  or (_24366_, _24365_, _24362_);
  or (_24367_, _24366_, _24359_);
  or (_24368_, _24367_, _24352_);
  and (_24369_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  and (_24370_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_24371_, _24370_, _24369_);
  and (_24372_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_24373_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_24374_, _24373_, _24372_);
  or (_24375_, _24374_, _24371_);
  and (_24376_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  and (_24377_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_24378_, _24377_, _24376_);
  and (_24379_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  and (_24380_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_24381_, _24380_, _24379_);
  or (_24382_, _24381_, _24378_);
  or (_24383_, _24382_, _24375_);
  and (_24384_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_24385_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_24386_, _24385_, _24384_);
  and (_24387_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  and (_24388_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_24389_, _24388_, _24387_);
  or (_24390_, _24389_, _24386_);
  and (_24391_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_24392_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_24393_, _24392_, _24391_);
  and (_24394_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  and (_24395_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_24396_, _24395_, _24394_);
  or (_24397_, _24396_, _24393_);
  or (_24398_, _24397_, _24390_);
  or (_24399_, _24398_, _24383_);
  or (_24400_, _24399_, _24368_);
  and (_24401_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  and (_24402_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_24403_, _24402_, _24401_);
  and (_24404_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_24405_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_24406_, _24405_, _24404_);
  or (_24407_, _24406_, _24403_);
  and (_24408_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_24409_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_24410_, _24409_, _24408_);
  and (_24411_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  and (_24412_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_24413_, _24412_, _24411_);
  or (_24414_, _24413_, _24410_);
  or (_24415_, _24414_, _24407_);
  and (_24416_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  and (_24417_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_24418_, _24417_, _24416_);
  and (_24419_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_24420_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_24421_, _24420_, _24419_);
  or (_24422_, _24421_, _24418_);
  and (_24423_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  and (_24424_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_24425_, _24424_, _24423_);
  and (_24426_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_24427_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_24428_, _24427_, _24426_);
  or (_24429_, _24428_, _24425_);
  or (_24430_, _24429_, _24422_);
  or (_24431_, _24430_, _24415_);
  and (_24432_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_24433_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_24434_, _24433_, _24432_);
  and (_24435_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and (_24436_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_24437_, _24436_, _24435_);
  or (_24438_, _24437_, _24434_);
  and (_24439_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_24440_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_24441_, _24440_, _24439_);
  and (_24442_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and (_24443_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_24444_, _24443_, _24442_);
  or (_24445_, _24444_, _24441_);
  or (_24446_, _24445_, _24438_);
  and (_24447_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_24448_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_24449_, _24448_, _24447_);
  and (_24450_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and (_24451_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_24452_, _24451_, _24450_);
  or (_24453_, _24452_, _24449_);
  and (_24454_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and (_24455_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_24456_, _24455_, _24454_);
  and (_24457_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and (_24458_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_24459_, _24458_, _24457_);
  or (_24460_, _24459_, _24456_);
  or (_24461_, _24460_, _24453_);
  or (_24462_, _24461_, _24446_);
  or (_24463_, _24462_, _24431_);
  or (_24464_, _24463_, _24400_);
  and (_24465_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  and (_24466_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_24467_, _24466_, _24465_);
  and (_24468_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_24469_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_24470_, _24469_, _24468_);
  or (_24471_, _24470_, _24467_);
  and (_24472_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  and (_24473_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_24474_, _24473_, _24472_);
  and (_24475_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_24476_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_24477_, _24476_, _24475_);
  or (_24478_, _24477_, _24474_);
  or (_24479_, _24478_, _24471_);
  and (_24480_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_24481_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_24482_, _24481_, _24480_);
  and (_24483_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  and (_24484_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_24485_, _24484_, _24483_);
  or (_24486_, _24485_, _24482_);
  and (_24487_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_24488_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_24489_, _24488_, _24487_);
  and (_24490_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  and (_24491_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_24492_, _24491_, _24490_);
  or (_24493_, _24492_, _24489_);
  or (_24494_, _24493_, _24486_);
  or (_24495_, _24494_, _24479_);
  and (_24496_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  and (_24497_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_24498_, _24497_, _24496_);
  and (_24499_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_24500_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_24501_, _24500_, _24499_);
  or (_24502_, _24501_, _24498_);
  and (_24503_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  and (_24504_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_24505_, _24504_, _24503_);
  and (_24506_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_24507_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_24508_, _24507_, _24506_);
  or (_24509_, _24508_, _24505_);
  or (_24510_, _24509_, _24502_);
  and (_24511_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_24512_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_24513_, _24512_, _24511_);
  and (_24514_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  and (_24515_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_24516_, _24515_, _24514_);
  or (_24517_, _24516_, _24513_);
  and (_24518_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_24519_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_24520_, _24519_, _24518_);
  and (_24521_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  and (_24522_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_24523_, _24522_, _24521_);
  or (_24524_, _24523_, _24520_);
  or (_24525_, _24524_, _24517_);
  or (_24526_, _24525_, _24510_);
  or (_24527_, _24526_, _24495_);
  and (_24528_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  and (_24529_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_24530_, _24529_, _24528_);
  and (_24531_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_24532_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_24533_, _24532_, _24531_);
  or (_24534_, _24533_, _24530_);
  and (_24535_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  and (_24536_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_24537_, _24536_, _24535_);
  and (_24538_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_24539_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_24540_, _24539_, _24538_);
  or (_24541_, _24540_, _24537_);
  or (_24542_, _24541_, _24534_);
  and (_24543_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_24544_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_24545_, _24544_, _24543_);
  and (_24546_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  and (_24547_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_24548_, _24547_, _24546_);
  or (_24549_, _24548_, _24545_);
  and (_24550_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_24551_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_24552_, _24551_, _24550_);
  and (_24553_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  and (_24554_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_24555_, _24554_, _24553_);
  or (_24556_, _24555_, _24552_);
  or (_24557_, _24556_, _24549_);
  or (_24558_, _24557_, _24542_);
  and (_24559_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_24560_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_24561_, _24560_, _24559_);
  and (_24562_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_24563_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_24564_, _24563_, _24562_);
  or (_24565_, _24564_, _24561_);
  and (_24566_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_24567_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_24568_, _24567_, _24566_);
  and (_24569_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_24570_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_24571_, _24570_, _24569_);
  or (_24572_, _24571_, _24568_);
  or (_24573_, _24572_, _24565_);
  and (_24574_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_24575_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_24576_, _24575_, _24574_);
  and (_24577_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_24578_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_24579_, _24578_, _24577_);
  or (_24580_, _24579_, _24576_);
  and (_24581_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_24582_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_24583_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_24584_, _24583_, _24582_);
  or (_24585_, _24584_, _24581_);
  or (_24586_, _24585_, _24580_);
  or (_24587_, _24586_, _24573_);
  or (_24588_, _24587_, _24558_);
  or (_24589_, _24588_, _24527_);
  or (_24590_, _24589_, _24464_);
  or (_24591_, _24590_, _24337_);
  and (_24592_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_24593_, _24592_, _24591_);
  and (_24594_, _24593_, _00006_);
  or (_24595_, _24594_, _24082_);
  and (_00003_[3], _24595_, _38997_);
  and (_24596_, _15589_, iram_op1[2]);
  and (_24597_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_24598_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or (_24599_, _24598_, _24597_);
  and (_24600_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_24601_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_24602_, _24601_, _24600_);
  or (_24603_, _24602_, _24599_);
  and (_24604_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_24605_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or (_24606_, _24605_, _24604_);
  and (_24607_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  and (_24608_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_24609_, _24608_, _24607_);
  or (_24610_, _24609_, _24606_);
  or (_24611_, _24610_, _24603_);
  and (_24612_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and (_24613_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_24614_, _24613_, _24612_);
  and (_24615_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_24616_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or (_24617_, _24616_, _24615_);
  or (_24618_, _24617_, _24614_);
  and (_24619_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  and (_24620_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_24621_, _24620_, _24619_);
  and (_24622_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_24623_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or (_24624_, _24623_, _24622_);
  or (_24625_, _24624_, _24621_);
  or (_24626_, _24625_, _24618_);
  or (_24627_, _24626_, _24611_);
  and (_24628_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  and (_24629_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_24630_, _24629_, _24628_);
  and (_24631_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_24632_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_24633_, _24632_, _24631_);
  or (_24634_, _24633_, _24630_);
  and (_24635_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  and (_24636_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_24637_, _24636_, _24635_);
  and (_24638_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_24639_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or (_24640_, _24639_, _24638_);
  or (_24641_, _24640_, _24637_);
  or (_24642_, _24641_, _24634_);
  and (_24643_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_24644_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or (_24645_, _24644_, _24643_);
  and (_24646_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and (_24647_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_24648_, _24647_, _24646_);
  or (_24649_, _24648_, _24645_);
  and (_24650_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_24651_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or (_24652_, _24651_, _24650_);
  and (_24653_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  and (_24654_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_24655_, _24654_, _24653_);
  or (_24656_, _24655_, _24652_);
  or (_24657_, _24656_, _24649_);
  or (_24658_, _24657_, _24642_);
  or (_24659_, _24658_, _24627_);
  and (_24660_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_24661_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  or (_24662_, _24661_, _24660_);
  and (_24663_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and (_24664_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_24665_, _24664_, _24663_);
  or (_24666_, _24665_, _24662_);
  and (_24667_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_24668_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  or (_24669_, _24668_, _24667_);
  and (_24670_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and (_24671_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  or (_24672_, _24671_, _24670_);
  or (_24673_, _24672_, _24669_);
  or (_24674_, _24673_, _24666_);
  and (_24675_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and (_24676_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_24677_, _24676_, _24675_);
  and (_24678_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_24679_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  or (_24680_, _24679_, _24678_);
  or (_24681_, _24680_, _24677_);
  and (_24682_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and (_24683_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_24684_, _24683_, _24682_);
  and (_24685_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_24686_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  or (_24687_, _24686_, _24685_);
  or (_24688_, _24687_, _24684_);
  or (_24689_, _24688_, _24681_);
  or (_24690_, _24689_, _24674_);
  and (_24691_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_24692_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_24693_, _24692_, _24691_);
  and (_24694_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  and (_24695_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_24696_, _24695_, _24694_);
  or (_24697_, _24696_, _24693_);
  and (_24698_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  and (_24699_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_24700_, _24699_, _24698_);
  and (_24701_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_24702_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or (_24703_, _24702_, _24701_);
  or (_24704_, _24703_, _24700_);
  or (_24705_, _24704_, _24697_);
  and (_24706_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_24707_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or (_24708_, _24707_, _24706_);
  and (_24709_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  and (_24710_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_24711_, _24710_, _24709_);
  or (_24712_, _24711_, _24708_);
  and (_24713_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_24714_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or (_24715_, _24714_, _24713_);
  and (_24716_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  and (_24717_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_24718_, _24717_, _24716_);
  or (_24719_, _24718_, _24715_);
  or (_24720_, _24719_, _24712_);
  or (_24721_, _24720_, _24705_);
  or (_24722_, _24721_, _24690_);
  or (_24723_, _24722_, _24659_);
  and (_24724_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_24725_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or (_24726_, _24725_, _24724_);
  and (_24727_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  and (_24728_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_24729_, _24728_, _24727_);
  or (_24730_, _24729_, _24726_);
  and (_24731_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_24732_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or (_24733_, _24732_, _24731_);
  and (_24734_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  and (_24735_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or (_24736_, _24735_, _24734_);
  or (_24737_, _24736_, _24733_);
  or (_24738_, _24737_, _24730_);
  and (_24739_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  and (_24740_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_24741_, _24740_, _24739_);
  and (_24742_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_24743_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  or (_24744_, _24743_, _24742_);
  or (_24745_, _24744_, _24741_);
  and (_24746_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  and (_24747_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_24748_, _24747_, _24746_);
  and (_24749_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_24750_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or (_24751_, _24750_, _24749_);
  or (_24752_, _24751_, _24748_);
  or (_24753_, _24752_, _24745_);
  or (_24754_, _24753_, _24738_);
  and (_24755_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and (_24756_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_24757_, _24756_, _24755_);
  and (_24758_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_24759_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  or (_24760_, _24759_, _24758_);
  or (_24761_, _24760_, _24757_);
  and (_24762_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_24763_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_24764_, _24763_, _24762_);
  and (_24765_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_24766_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_24767_, _24766_, _24765_);
  or (_24768_, _24767_, _24764_);
  or (_24769_, _24768_, _24761_);
  and (_24770_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_24771_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  or (_24772_, _24771_, _24770_);
  and (_24773_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_24774_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_24775_, _24774_, _24773_);
  or (_24776_, _24775_, _24772_);
  and (_24777_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_24778_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  or (_24779_, _24778_, _24777_);
  and (_24780_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and (_24781_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_24782_, _24781_, _24780_);
  or (_24783_, _24782_, _24779_);
  or (_24784_, _24783_, _24776_);
  or (_24785_, _24784_, _24769_);
  or (_24786_, _24785_, _24754_);
  and (_24787_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_24788_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or (_24789_, _24788_, _24787_);
  and (_24790_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and (_24791_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_24792_, _24791_, _24790_);
  or (_24793_, _24792_, _24789_);
  and (_24794_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_24795_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or (_24796_, _24795_, _24794_);
  and (_24797_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  and (_24798_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or (_24799_, _24798_, _24797_);
  or (_24800_, _24799_, _24796_);
  or (_24801_, _24800_, _24793_);
  and (_24802_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and (_24803_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_24804_, _24803_, _24802_);
  and (_24805_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_24806_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or (_24807_, _24806_, _24805_);
  or (_24808_, _24807_, _24804_);
  and (_24809_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and (_24810_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_24811_, _24810_, _24809_);
  and (_24812_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_24813_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_24814_, _24813_, _24812_);
  or (_24815_, _24814_, _24811_);
  or (_24816_, _24815_, _24808_);
  or (_24817_, _24816_, _24801_);
  and (_24818_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  and (_24819_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_24820_, _24819_, _24818_);
  and (_24821_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_24822_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_24823_, _24822_, _24821_);
  or (_24824_, _24823_, _24820_);
  and (_24825_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and (_24826_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_24827_, _24826_, _24825_);
  and (_24828_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and (_24829_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_24830_, _24829_, _24828_);
  or (_24831_, _24830_, _24827_);
  or (_24832_, _24831_, _24824_);
  and (_24833_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_24834_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_24835_, _24834_, _24833_);
  and (_24836_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  and (_24837_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_24838_, _24837_, _24836_);
  or (_24839_, _24838_, _24835_);
  and (_24840_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_24841_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_24842_, _24841_, _24840_);
  and (_24843_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  and (_24844_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_24845_, _24844_, _24843_);
  or (_24846_, _24845_, _24842_);
  or (_24847_, _24846_, _24839_);
  or (_24848_, _24847_, _24832_);
  or (_24849_, _24848_, _24817_);
  or (_24850_, _24849_, _24786_);
  or (_24851_, _24850_, _24723_);
  and (_24852_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_24853_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or (_24854_, _24853_, _24852_);
  and (_24855_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  and (_24856_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_24857_, _24856_, _24855_);
  or (_24858_, _24857_, _24854_);
  and (_24859_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_24860_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or (_24861_, _24860_, _24859_);
  and (_24862_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_24863_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_24864_, _24863_, _24862_);
  or (_24865_, _24864_, _24861_);
  or (_24866_, _24865_, _24858_);
  and (_24867_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  and (_24868_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_24869_, _24868_, _24867_);
  and (_24870_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_24871_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or (_24872_, _24871_, _24870_);
  or (_24873_, _24872_, _24869_);
  and (_24874_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_24875_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or (_24876_, _24875_, _24874_);
  and (_24877_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  and (_24878_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_24879_, _24878_, _24877_);
  or (_24880_, _24879_, _24876_);
  or (_24881_, _24880_, _24873_);
  or (_24882_, _24881_, _24866_);
  and (_24883_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  and (_24884_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_24885_, _24884_, _24883_);
  and (_24886_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_24887_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_24888_, _24887_, _24886_);
  or (_24889_, _24888_, _24885_);
  and (_24890_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  and (_24891_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_24892_, _24891_, _24890_);
  and (_24893_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  and (_24894_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_24895_, _24894_, _24893_);
  or (_24896_, _24895_, _24892_);
  or (_24897_, _24896_, _24889_);
  and (_24898_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_24899_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_24900_, _24899_, _24898_);
  and (_24901_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  and (_24902_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_24903_, _24902_, _24901_);
  or (_24904_, _24903_, _24900_);
  and (_24905_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_24906_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_24907_, _24906_, _24905_);
  and (_24908_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  and (_24909_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_24910_, _24909_, _24908_);
  or (_24911_, _24910_, _24907_);
  or (_24912_, _24911_, _24904_);
  or (_24913_, _24912_, _24897_);
  or (_24914_, _24913_, _24882_);
  and (_24915_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_24916_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_24917_, _24916_, _24915_);
  and (_24918_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  and (_24919_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_24920_, _24919_, _24918_);
  or (_24921_, _24920_, _24917_);
  and (_24922_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_24923_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_24924_, _24923_, _24922_);
  and (_24925_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  and (_24926_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_24927_, _24926_, _24925_);
  or (_24928_, _24927_, _24924_);
  or (_24929_, _24928_, _24921_);
  and (_24930_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_24931_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_24932_, _24931_, _24930_);
  and (_24933_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  and (_24934_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_24935_, _24934_, _24933_);
  or (_24936_, _24935_, _24932_);
  and (_24937_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  and (_24938_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_24939_, _24938_, _24937_);
  and (_24940_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_24941_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_24942_, _24941_, _24940_);
  or (_24943_, _24942_, _24939_);
  or (_24944_, _24943_, _24936_);
  or (_24945_, _24944_, _24929_);
  and (_24946_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and (_24947_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_24948_, _24947_, _24946_);
  and (_24949_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_24950_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_24951_, _24950_, _24949_);
  or (_24952_, _24951_, _24948_);
  and (_24953_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and (_24954_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_24955_, _24954_, _24953_);
  and (_24956_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_24957_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_24958_, _24957_, _24956_);
  or (_24959_, _24958_, _24955_);
  or (_24960_, _24959_, _24952_);
  and (_24961_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_24962_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_24963_, _24962_, _24961_);
  and (_24964_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and (_24965_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_24966_, _24965_, _24964_);
  or (_24967_, _24966_, _24963_);
  and (_24968_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_24969_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_24970_, _24969_, _24968_);
  and (_24971_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and (_24972_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_24973_, _24972_, _24971_);
  or (_24974_, _24973_, _24970_);
  or (_24975_, _24974_, _24967_);
  or (_24976_, _24975_, _24960_);
  or (_24977_, _24976_, _24945_);
  or (_24978_, _24977_, _24914_);
  and (_24979_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  and (_24980_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_24981_, _24980_, _24979_);
  and (_24982_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_24983_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or (_24984_, _24983_, _24982_);
  or (_24985_, _24984_, _24981_);
  and (_24986_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_24987_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_24988_, _24987_, _24986_);
  and (_24989_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  and (_24990_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_24991_, _24990_, _24989_);
  or (_24992_, _24991_, _24988_);
  or (_24993_, _24992_, _24985_);
  and (_24994_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_24995_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_24996_, _24995_, _24994_);
  and (_24997_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  and (_24998_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_24999_, _24998_, _24997_);
  or (_25000_, _24999_, _24996_);
  and (_25001_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_25002_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_25003_, _25002_, _25001_);
  and (_25004_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  and (_25005_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_25006_, _25005_, _25004_);
  or (_25007_, _25006_, _25003_);
  or (_25008_, _25007_, _25000_);
  or (_25009_, _25008_, _24993_);
  and (_25010_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  and (_25011_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_25012_, _25011_, _25010_);
  and (_25013_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  and (_25014_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_25015_, _25014_, _25013_);
  or (_25016_, _25015_, _25012_);
  and (_25017_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  and (_25018_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_25019_, _25018_, _25017_);
  and (_25020_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_25021_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_25022_, _25021_, _25020_);
  or (_25023_, _25022_, _25019_);
  or (_25024_, _25023_, _25016_);
  and (_25025_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_25026_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_25027_, _25026_, _25025_);
  and (_25028_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  and (_25029_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_25030_, _25029_, _25028_);
  or (_25031_, _25030_, _25027_);
  and (_25032_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_25033_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_25034_, _25033_, _25032_);
  and (_25035_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  and (_25036_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_25037_, _25036_, _25035_);
  or (_25038_, _25037_, _25034_);
  or (_25039_, _25038_, _25031_);
  or (_25040_, _25039_, _25024_);
  or (_25041_, _25040_, _25009_);
  and (_25042_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_25043_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_25044_, _25043_, _25042_);
  and (_25045_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  and (_25046_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_25047_, _25046_, _25045_);
  or (_25048_, _25047_, _25044_);
  and (_25049_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_25050_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_25051_, _25050_, _25049_);
  and (_25052_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_25053_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_25054_, _25053_, _25052_);
  or (_25055_, _25054_, _25051_);
  or (_25056_, _25055_, _25048_);
  and (_25057_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  and (_25058_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_25059_, _25058_, _25057_);
  and (_25060_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_25061_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_25062_, _25061_, _25060_);
  or (_25063_, _25062_, _25059_);
  and (_25064_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  and (_25065_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_25066_, _25065_, _25064_);
  and (_25067_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_25068_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_25069_, _25068_, _25067_);
  or (_25070_, _25069_, _25066_);
  or (_25071_, _25070_, _25063_);
  or (_25072_, _25071_, _25056_);
  and (_25073_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_25074_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_25075_, _25074_, _25073_);
  and (_25076_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_25077_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_25078_, _25077_, _25076_);
  or (_25079_, _25078_, _25075_);
  and (_25080_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_25081_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_25082_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_25083_, _25082_, _25081_);
  or (_25084_, _25083_, _25080_);
  or (_25085_, _25084_, _25079_);
  and (_25086_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_25087_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_25088_, _25087_, _25086_);
  and (_25089_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_25090_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_25091_, _25090_, _25089_);
  or (_25092_, _25091_, _25088_);
  and (_25093_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_25094_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_25095_, _25094_, _25093_);
  and (_25096_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_25097_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_25098_, _25097_, _25096_);
  or (_25099_, _25098_, _25095_);
  or (_25100_, _25099_, _25092_);
  or (_25101_, _25100_, _25085_);
  or (_25102_, _25101_, _25072_);
  or (_25103_, _25102_, _25041_);
  or (_25104_, _25103_, _24978_);
  or (_25105_, _25104_, _24851_);
  and (_25106_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_25107_, _25106_, _25105_);
  and (_25108_, _25107_, _00006_);
  or (_25109_, _25108_, _24596_);
  and (_00003_[2], _25109_, _38997_);
  and (_25110_, _15589_, iram_op1[1]);
  and (_25111_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  and (_25112_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_25113_, _25112_, _25111_);
  and (_25114_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_25115_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or (_25116_, _25115_, _25114_);
  or (_25117_, _25116_, _25113_);
  and (_25118_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and (_25119_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_25120_, _25119_, _25118_);
  and (_25121_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_25122_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or (_25123_, _25122_, _25121_);
  or (_25124_, _25123_, _25120_);
  or (_25125_, _25124_, _25117_);
  and (_25126_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_25127_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or (_25128_, _25127_, _25126_);
  and (_25129_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  and (_25130_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_25131_, _25130_, _25129_);
  or (_25132_, _25131_, _25128_);
  and (_25133_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_25134_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or (_25135_, _25134_, _25133_);
  and (_25136_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_25137_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_25138_, _25137_, _25136_);
  or (_25139_, _25138_, _25135_);
  or (_25140_, _25139_, _25132_);
  or (_25141_, _25140_, _25125_);
  and (_25142_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  and (_25143_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_25144_, _25143_, _25142_);
  and (_25145_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_25146_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or (_25147_, _25146_, _25145_);
  or (_25148_, _25147_, _25144_);
  and (_25149_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  and (_25150_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_25151_, _25150_, _25149_);
  and (_25152_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_25153_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_25154_, _25153_, _25152_);
  or (_25155_, _25154_, _25151_);
  or (_25156_, _25155_, _25148_);
  and (_25157_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_25158_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or (_25159_, _25158_, _25157_);
  and (_25160_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  and (_25161_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_25162_, _25161_, _25160_);
  or (_25163_, _25162_, _25159_);
  and (_25164_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_25165_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or (_25166_, _25165_, _25164_);
  and (_25167_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  and (_25168_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_25169_, _25168_, _25167_);
  or (_25170_, _25169_, _25166_);
  or (_25171_, _25170_, _25163_);
  or (_25172_, _25171_, _25156_);
  or (_25173_, _25172_, _25141_);
  and (_25174_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_25175_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  or (_25176_, _25175_, _25174_);
  and (_25177_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and (_25178_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_25179_, _25178_, _25177_);
  or (_25180_, _25179_, _25176_);
  and (_25181_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_25182_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  or (_25183_, _25182_, _25181_);
  and (_25184_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_25185_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_25186_, _25185_, _25184_);
  or (_25187_, _25186_, _25183_);
  or (_25188_, _25187_, _25180_);
  and (_25189_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and (_25190_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_25191_, _25190_, _25189_);
  and (_25192_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_25193_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or (_25194_, _25193_, _25192_);
  or (_25195_, _25194_, _25191_);
  and (_25196_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and (_25197_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_25198_, _25197_, _25196_);
  and (_25199_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_25200_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  or (_25201_, _25200_, _25199_);
  or (_25202_, _25201_, _25198_);
  or (_25203_, _25202_, _25195_);
  or (_25204_, _25203_, _25188_);
  and (_25205_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  and (_25206_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_25207_, _25206_, _25205_);
  and (_25208_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_25209_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or (_25210_, _25209_, _25208_);
  or (_25211_, _25210_, _25207_);
  and (_25212_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  and (_25213_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_25214_, _25213_, _25212_);
  and (_25215_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_25216_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_25217_, _25216_, _25215_);
  or (_25218_, _25217_, _25214_);
  or (_25219_, _25218_, _25211_);
  and (_25220_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_25221_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or (_25222_, _25221_, _25220_);
  and (_25223_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  and (_25224_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_25225_, _25224_, _25223_);
  or (_25226_, _25225_, _25222_);
  and (_25227_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_25228_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or (_25229_, _25228_, _25227_);
  and (_25230_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  and (_25231_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_25232_, _25231_, _25230_);
  or (_25233_, _25232_, _25229_);
  or (_25234_, _25233_, _25226_);
  or (_25235_, _25234_, _25219_);
  or (_25236_, _25235_, _25204_);
  or (_25237_, _25236_, _25173_);
  and (_25238_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  and (_25239_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_25240_, _25239_, _25238_);
  and (_25241_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_25242_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  or (_25243_, _25242_, _25241_);
  or (_25244_, _25243_, _25240_);
  and (_25245_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  and (_25246_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_25247_, _25246_, _25245_);
  and (_25248_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_25249_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or (_25250_, _25249_, _25248_);
  or (_25251_, _25250_, _25247_);
  or (_25252_, _25251_, _25244_);
  and (_25253_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_25254_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or (_25255_, _25254_, _25253_);
  and (_25256_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  and (_25257_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or (_25258_, _25257_, _25256_);
  or (_25259_, _25258_, _25255_);
  and (_25260_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_25261_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or (_25262_, _25261_, _25260_);
  and (_25263_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  and (_25264_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_25265_, _25264_, _25263_);
  or (_25266_, _25265_, _25262_);
  or (_25267_, _25266_, _25259_);
  or (_25268_, _25267_, _25252_);
  and (_25269_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and (_25270_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_25271_, _25270_, _25269_);
  and (_25272_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_25273_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  or (_25274_, _25273_, _25272_);
  or (_25275_, _25274_, _25271_);
  and (_25276_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_25277_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_25278_, _25277_, _25276_);
  and (_25279_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_25280_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_25281_, _25280_, _25279_);
  or (_25282_, _25281_, _25278_);
  or (_25283_, _25282_, _25275_);
  and (_25284_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_25285_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  or (_25286_, _25285_, _25284_);
  and (_25287_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_25288_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_25289_, _25288_, _25287_);
  or (_25290_, _25289_, _25286_);
  and (_25291_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_25292_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  or (_25293_, _25292_, _25291_);
  and (_25294_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and (_25295_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_25296_, _25295_, _25294_);
  or (_25297_, _25296_, _25293_);
  or (_25298_, _25297_, _25290_);
  or (_25299_, _25298_, _25283_);
  or (_25300_, _25299_, _25268_);
  and (_25301_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  and (_25302_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_25303_, _25302_, _25301_);
  and (_25304_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_25305_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_25306_, _25305_, _25304_);
  or (_25307_, _25306_, _25303_);
  and (_25308_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and (_25309_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_25310_, _25309_, _25308_);
  and (_25311_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_25312_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_25313_, _25312_, _25311_);
  or (_25314_, _25313_, _25310_);
  or (_25315_, _25314_, _25307_);
  and (_25316_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_25317_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_25318_, _25317_, _25316_);
  and (_25319_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and (_25320_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_25321_, _25320_, _25319_);
  or (_25322_, _25321_, _25318_);
  and (_25323_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_25324_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_25325_, _25324_, _25323_);
  and (_25326_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and (_25327_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_25328_, _25327_, _25326_);
  or (_25329_, _25328_, _25325_);
  or (_25330_, _25329_, _25322_);
  or (_25331_, _25330_, _25315_);
  and (_25332_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_25333_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or (_25334_, _25333_, _25332_);
  and (_25335_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and (_25336_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_25337_, _25336_, _25335_);
  or (_25338_, _25337_, _25334_);
  and (_25339_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_25340_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or (_25341_, _25340_, _25339_);
  and (_25342_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and (_25343_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or (_25344_, _25343_, _25342_);
  or (_25345_, _25344_, _25341_);
  or (_25346_, _25345_, _25338_);
  and (_25347_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  and (_25348_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_25349_, _25348_, _25347_);
  and (_25350_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_25351_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or (_25352_, _25351_, _25350_);
  or (_25353_, _25352_, _25349_);
  and (_25354_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and (_25355_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_25356_, _25355_, _25354_);
  and (_25357_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_25358_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_25359_, _25358_, _25357_);
  or (_25360_, _25359_, _25356_);
  or (_25361_, _25360_, _25353_);
  or (_25362_, _25361_, _25346_);
  or (_25363_, _25362_, _25331_);
  or (_25364_, _25363_, _25300_);
  or (_25365_, _25364_, _25237_);
  and (_25366_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  and (_25367_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_25368_, _25367_, _25366_);
  and (_25369_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_25370_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or (_25371_, _25370_, _25369_);
  or (_25372_, _25371_, _25368_);
  and (_25373_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  and (_25374_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_25375_, _25374_, _25373_);
  and (_25376_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_25377_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or (_25378_, _25377_, _25376_);
  or (_25379_, _25378_, _25375_);
  or (_25380_, _25379_, _25372_);
  and (_25381_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_25382_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or (_25383_, _25382_, _25381_);
  and (_25384_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  and (_25385_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or (_25386_, _25385_, _25384_);
  or (_25387_, _25386_, _25383_);
  and (_25388_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_25389_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or (_25390_, _25389_, _25388_);
  and (_25391_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  and (_25392_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_25393_, _25392_, _25391_);
  or (_25394_, _25393_, _25390_);
  or (_25395_, _25394_, _25387_);
  or (_25396_, _25395_, _25380_);
  and (_25397_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  and (_25398_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_25399_, _25398_, _25397_);
  and (_25400_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_25401_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_25402_, _25401_, _25400_);
  or (_25403_, _25402_, _25399_);
  and (_25404_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  and (_25405_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_25406_, _25405_, _25404_);
  and (_25407_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_25408_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_25409_, _25408_, _25407_);
  or (_25410_, _25409_, _25406_);
  or (_25411_, _25410_, _25403_);
  and (_25412_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_25413_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_25414_, _25413_, _25412_);
  and (_25415_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  and (_25416_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_25417_, _25416_, _25415_);
  or (_25418_, _25417_, _25414_);
  and (_25419_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_25420_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_25421_, _25420_, _25419_);
  and (_25422_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  and (_25423_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_25424_, _25423_, _25422_);
  or (_25425_, _25424_, _25421_);
  or (_25426_, _25425_, _25418_);
  or (_25427_, _25426_, _25411_);
  or (_25428_, _25427_, _25396_);
  and (_25429_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  and (_25430_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_25431_, _25430_, _25429_);
  and (_25432_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and (_25433_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_25434_, _25433_, _25432_);
  or (_25435_, _25434_, _25431_);
  and (_25436_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  and (_25437_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_25438_, _25437_, _25436_);
  and (_25439_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_25440_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_25441_, _25440_, _25439_);
  or (_25442_, _25441_, _25438_);
  or (_25443_, _25442_, _25435_);
  and (_25444_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_25445_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_25446_, _25445_, _25444_);
  and (_25447_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  and (_25448_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_25449_, _25448_, _25447_);
  or (_25450_, _25449_, _25446_);
  and (_25451_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_25452_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_25453_, _25452_, _25451_);
  and (_25454_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  and (_25455_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_25456_, _25455_, _25454_);
  or (_25457_, _25456_, _25453_);
  or (_25458_, _25457_, _25450_);
  or (_25459_, _25458_, _25443_);
  and (_25460_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and (_25461_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_25462_, _25461_, _25460_);
  and (_25463_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_25464_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_25465_, _25464_, _25463_);
  or (_25466_, _25465_, _25462_);
  and (_25467_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and (_25468_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_25469_, _25468_, _25467_);
  and (_25470_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and (_25471_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_25472_, _25471_, _25470_);
  or (_25473_, _25472_, _25469_);
  or (_25474_, _25473_, _25466_);
  and (_25475_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and (_25476_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_25477_, _25476_, _25475_);
  and (_25478_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and (_25479_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_25480_, _25479_, _25478_);
  or (_25481_, _25480_, _25477_);
  and (_25482_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_25483_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_25484_, _25483_, _25482_);
  and (_25485_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  and (_25486_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_25487_, _25486_, _25485_);
  or (_25488_, _25487_, _25484_);
  or (_25489_, _25488_, _25481_);
  or (_25490_, _25489_, _25474_);
  or (_25491_, _25490_, _25459_);
  or (_25492_, _25491_, _25428_);
  and (_25493_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_25494_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_25495_, _25494_, _25493_);
  and (_25496_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  and (_25497_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_25498_, _25497_, _25496_);
  or (_25499_, _25498_, _25495_);
  and (_25500_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_25501_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_25502_, _25501_, _25500_);
  and (_25503_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  and (_25504_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_25505_, _25504_, _25503_);
  or (_25506_, _25505_, _25502_);
  or (_25507_, _25506_, _25499_);
  and (_25508_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  and (_25509_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_25510_, _25509_, _25508_);
  and (_25511_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_25512_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_25513_, _25512_, _25511_);
  or (_25514_, _25513_, _25510_);
  and (_25515_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  and (_25516_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_25517_, _25516_, _25515_);
  and (_25518_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_25519_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_25520_, _25519_, _25518_);
  or (_25521_, _25520_, _25517_);
  or (_25522_, _25521_, _25514_);
  or (_25523_, _25522_, _25507_);
  and (_25524_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  and (_25525_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_25526_, _25525_, _25524_);
  and (_25527_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_25528_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_25529_, _25528_, _25527_);
  or (_25530_, _25529_, _25526_);
  and (_25531_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  and (_25532_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_25533_, _25532_, _25531_);
  and (_25534_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_25535_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_25536_, _25535_, _25534_);
  or (_25537_, _25536_, _25533_);
  or (_25538_, _25537_, _25530_);
  and (_25539_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_25540_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_25541_, _25540_, _25539_);
  and (_25542_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  and (_25543_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_25544_, _25543_, _25542_);
  or (_25545_, _25544_, _25541_);
  and (_25546_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_25547_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_25548_, _25547_, _25546_);
  and (_25549_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  and (_25550_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_25551_, _25550_, _25549_);
  or (_25552_, _25551_, _25548_);
  or (_25553_, _25552_, _25545_);
  or (_25554_, _25553_, _25538_);
  or (_25555_, _25554_, _25523_);
  and (_25556_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  and (_25557_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_25558_, _25557_, _25556_);
  and (_25559_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_25560_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_25561_, _25560_, _25559_);
  or (_25562_, _25561_, _25558_);
  and (_25563_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  and (_25564_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_25565_, _25564_, _25563_);
  and (_25566_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_25567_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_25568_, _25567_, _25566_);
  or (_25569_, _25568_, _25565_);
  or (_25570_, _25569_, _25562_);
  and (_25571_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_25572_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_25573_, _25572_, _25571_);
  and (_25574_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  and (_25575_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_25576_, _25575_, _25574_);
  or (_25577_, _25576_, _25573_);
  and (_25578_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_25579_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_25580_, _25579_, _25578_);
  and (_25581_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  and (_25582_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_25583_, _25582_, _25581_);
  or (_25584_, _25583_, _25580_);
  or (_25585_, _25584_, _25577_);
  or (_25586_, _25585_, _25570_);
  and (_25587_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_25588_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_25589_, _25588_, _25587_);
  and (_25590_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_25591_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_25592_, _25591_, _25590_);
  or (_25593_, _25592_, _25589_);
  and (_25594_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_25595_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_25596_, _25595_, _25594_);
  and (_25597_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_25598_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_25599_, _25598_, _25597_);
  or (_25600_, _25599_, _25596_);
  or (_25601_, _25600_, _25593_);
  and (_25602_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_25603_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_25604_, _25603_, _25602_);
  and (_25605_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_25606_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_25607_, _25606_, _25605_);
  or (_25608_, _25607_, _25604_);
  and (_25609_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_25610_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_25611_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_25612_, _25611_, _25610_);
  or (_25613_, _25612_, _25609_);
  or (_25614_, _25613_, _25608_);
  or (_25615_, _25614_, _25601_);
  or (_25616_, _25615_, _25586_);
  or (_25617_, _25616_, _25555_);
  or (_25618_, _25617_, _25492_);
  or (_25619_, _25618_, _25365_);
  and (_25620_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_25621_, _25620_, _25619_);
  and (_25622_, _25621_, _00006_);
  or (_25623_, _25622_, _25110_);
  and (_00003_[1], _25623_, _38997_);
  and (_25624_, _15589_, iram_op1[0]);
  and (_25625_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_25626_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or (_25627_, _25626_, _25625_);
  and (_25628_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and (_25629_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_25630_, _25629_, _25628_);
  or (_25631_, _25630_, _25627_);
  and (_25632_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_25633_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or (_25634_, _25633_, _25632_);
  and (_25635_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  and (_25636_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_25637_, _25636_, _25635_);
  or (_25638_, _25637_, _25634_);
  or (_25639_, _25638_, _25631_);
  and (_25640_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  and (_25641_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_25642_, _25641_, _25640_);
  and (_25643_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_25644_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_25645_, _25644_, _25643_);
  or (_25646_, _25645_, _25642_);
  and (_25647_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  and (_25648_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_25649_, _25648_, _25647_);
  and (_25650_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_25651_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or (_25652_, _25651_, _25650_);
  or (_25653_, _25652_, _25649_);
  or (_25654_, _25653_, _25646_);
  or (_25655_, _25654_, _25639_);
  and (_25656_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_25657_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or (_25658_, _25657_, _25656_);
  and (_25659_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and (_25660_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_25661_, _25660_, _25659_);
  or (_25662_, _25661_, _25658_);
  and (_25663_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_25664_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or (_25665_, _25664_, _25663_);
  and (_25666_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  and (_25667_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or (_25668_, _25667_, _25666_);
  or (_25669_, _25668_, _25665_);
  or (_25670_, _25669_, _25662_);
  and (_25671_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  and (_25672_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_25673_, _25672_, _25671_);
  and (_25674_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_25675_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or (_25676_, _25675_, _25674_);
  or (_25677_, _25676_, _25673_);
  and (_25678_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  and (_25679_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_25680_, _25679_, _25678_);
  and (_25681_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_25682_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or (_25683_, _25682_, _25681_);
  or (_25684_, _25683_, _25680_);
  or (_25685_, _25684_, _25677_);
  or (_25686_, _25685_, _25670_);
  or (_25687_, _25686_, _25655_);
  and (_25688_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_25689_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  or (_25690_, _25689_, _25688_);
  and (_25691_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_25692_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_25693_, _25692_, _25691_);
  or (_25694_, _25693_, _25690_);
  and (_25695_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_25696_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  or (_25697_, _25696_, _25695_);
  and (_25698_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and (_25699_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_25700_, _25699_, _25698_);
  or (_25701_, _25700_, _25697_);
  or (_25702_, _25701_, _25694_);
  and (_25703_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and (_25704_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_25705_, _25704_, _25703_);
  and (_25706_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_25707_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  or (_25708_, _25707_, _25706_);
  or (_25709_, _25708_, _25705_);
  and (_25710_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and (_25711_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_25712_, _25711_, _25710_);
  and (_25713_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_25714_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_25715_, _25714_, _25713_);
  or (_25716_, _25715_, _25712_);
  or (_25717_, _25716_, _25709_);
  or (_25718_, _25717_, _25702_);
  and (_25719_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_25720_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_25721_, _25720_, _25719_);
  and (_25722_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  and (_25723_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_25724_, _25723_, _25722_);
  or (_25725_, _25724_, _25721_);
  and (_25726_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_25727_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_25728_, _25727_, _25726_);
  and (_25729_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  and (_25730_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_25731_, _25730_, _25729_);
  or (_25732_, _25731_, _25728_);
  or (_25733_, _25732_, _25725_);
  and (_25734_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  and (_25735_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_25736_, _25735_, _25734_);
  and (_25737_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  and (_25738_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_25739_, _25738_, _25737_);
  or (_25740_, _25739_, _25736_);
  and (_25741_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  and (_25742_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_25743_, _25742_, _25741_);
  and (_25744_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_25745_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_25746_, _25745_, _25744_);
  or (_25747_, _25746_, _25743_);
  or (_25748_, _25747_, _25740_);
  or (_25749_, _25748_, _25733_);
  or (_25750_, _25749_, _25718_);
  or (_25751_, _25750_, _25687_);
  and (_25752_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  and (_25753_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_25754_, _25753_, _25752_);
  and (_25755_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_25756_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or (_25757_, _25756_, _25755_);
  or (_25758_, _25757_, _25754_);
  and (_25759_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  and (_25760_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_25761_, _25760_, _25759_);
  and (_25762_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_25763_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or (_25764_, _25763_, _25762_);
  or (_25765_, _25764_, _25761_);
  or (_25766_, _25765_, _25758_);
  and (_25767_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_25768_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or (_25769_, _25768_, _25767_);
  and (_25770_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  and (_25771_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or (_25772_, _25771_, _25770_);
  or (_25773_, _25772_, _25769_);
  and (_25774_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_25775_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or (_25776_, _25775_, _25774_);
  and (_25777_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  and (_25778_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_25779_, _25778_, _25777_);
  or (_25780_, _25779_, _25776_);
  or (_25781_, _25780_, _25773_);
  or (_25782_, _25781_, _25766_);
  and (_25783_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_25784_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_25785_, _25784_, _25783_);
  and (_25786_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_25787_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  or (_25788_, _25787_, _25786_);
  or (_25789_, _25788_, _25785_);
  and (_25790_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_25791_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_25792_, _25791_, _25790_);
  and (_25793_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_25794_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_25795_, _25794_, _25793_);
  or (_25796_, _25795_, _25792_);
  or (_25797_, _25796_, _25789_);
  and (_25798_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_25799_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  or (_25800_, _25799_, _25798_);
  and (_25801_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_25802_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_25803_, _25802_, _25801_);
  or (_25804_, _25803_, _25800_);
  and (_25805_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_25806_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  or (_25807_, _25806_, _25805_);
  and (_25808_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and (_25809_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_25810_, _25809_, _25808_);
  or (_25811_, _25810_, _25807_);
  or (_25812_, _25811_, _25804_);
  or (_25813_, _25812_, _25797_);
  or (_25814_, _25813_, _25782_);
  and (_25815_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  and (_25816_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_25817_, _25816_, _25815_);
  and (_25818_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_25819_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or (_25820_, _25819_, _25818_);
  or (_25821_, _25820_, _25817_);
  and (_25822_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  and (_25823_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_25824_, _25823_, _25822_);
  and (_25825_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_25826_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or (_25827_, _25826_, _25825_);
  or (_25828_, _25827_, _25824_);
  or (_25829_, _25828_, _25821_);
  and (_25830_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_25831_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or (_25832_, _25831_, _25830_);
  and (_25833_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and (_25834_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_25835_, _25834_, _25833_);
  or (_25836_, _25835_, _25832_);
  and (_25837_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_25838_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or (_25839_, _25838_, _25837_);
  and (_25840_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and (_25841_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or (_25842_, _25841_, _25840_);
  or (_25843_, _25842_, _25839_);
  or (_25844_, _25843_, _25836_);
  or (_25845_, _25844_, _25829_);
  and (_25846_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_25847_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or (_25848_, _25847_, _25846_);
  and (_25849_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  and (_25850_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_25851_, _25850_, _25849_);
  or (_25852_, _25851_, _25848_);
  and (_25853_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_25854_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or (_25855_, _25854_, _25853_);
  and (_25856_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and (_25857_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_25858_, _25857_, _25856_);
  or (_25859_, _25858_, _25855_);
  or (_25860_, _25859_, _25852_);
  and (_25861_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  and (_25862_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_25863_, _25862_, _25861_);
  and (_25864_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_25865_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or (_25866_, _25865_, _25864_);
  or (_25867_, _25866_, _25863_);
  and (_25868_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  and (_25869_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_25870_, _25869_, _25868_);
  and (_25871_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_25872_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_25873_, _25872_, _25871_);
  or (_25874_, _25873_, _25870_);
  or (_25875_, _25874_, _25867_);
  or (_25876_, _25875_, _25860_);
  or (_25877_, _25876_, _25845_);
  or (_25878_, _25877_, _25814_);
  or (_25879_, _25878_, _25751_);
  and (_25880_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_25881_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or (_25882_, _25881_, _25880_);
  and (_25883_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  and (_25884_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_25885_, _25884_, _25883_);
  or (_25886_, _25885_, _25882_);
  and (_25887_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_25888_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or (_25889_, _25888_, _25887_);
  and (_25890_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_25891_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_25892_, _25891_, _25890_);
  or (_25893_, _25892_, _25889_);
  or (_25894_, _25893_, _25886_);
  and (_25895_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  and (_25896_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_25897_, _25896_, _25895_);
  and (_25898_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_25899_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or (_25900_, _25899_, _25898_);
  or (_25901_, _25900_, _25897_);
  and (_25902_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  and (_25903_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_25904_, _25903_, _25902_);
  and (_25905_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_25906_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or (_25907_, _25906_, _25905_);
  or (_25908_, _25907_, _25904_);
  or (_25909_, _25908_, _25901_);
  or (_25910_, _25909_, _25894_);
  and (_25911_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  and (_25912_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_25913_, _25912_, _25911_);
  and (_25914_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_25915_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_25916_, _25915_, _25914_);
  or (_25917_, _25916_, _25913_);
  and (_25918_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  and (_25919_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_25920_, _25919_, _25918_);
  and (_25921_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_25922_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_25923_, _25922_, _25921_);
  or (_25924_, _25923_, _25920_);
  or (_25925_, _25924_, _25917_);
  and (_25926_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_25927_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_25928_, _25927_, _25926_);
  and (_25929_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  and (_25930_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_25931_, _25930_, _25929_);
  or (_25932_, _25931_, _25928_);
  and (_25933_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_25934_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_25935_, _25934_, _25933_);
  and (_25936_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  and (_25937_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_25938_, _25937_, _25936_);
  or (_25939_, _25938_, _25935_);
  or (_25940_, _25939_, _25932_);
  or (_25941_, _25940_, _25925_);
  or (_25942_, _25941_, _25910_);
  and (_25943_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_25944_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_25945_, _25944_, _25943_);
  and (_25946_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  and (_25947_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_25948_, _25947_, _25946_);
  or (_25949_, _25948_, _25945_);
  and (_25950_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_25951_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_25952_, _25951_, _25950_);
  and (_25953_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_25954_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_25955_, _25954_, _25953_);
  or (_25956_, _25955_, _25952_);
  or (_25957_, _25956_, _25949_);
  and (_25958_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  and (_25959_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_25960_, _25959_, _25958_);
  and (_25961_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_25962_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_25963_, _25962_, _25961_);
  or (_25964_, _25963_, _25960_);
  and (_25965_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  and (_25966_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_25967_, _25966_, _25965_);
  and (_25968_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_25969_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_25970_, _25969_, _25968_);
  or (_25971_, _25970_, _25967_);
  or (_25972_, _25971_, _25964_);
  or (_25973_, _25972_, _25957_);
  and (_25974_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  and (_25975_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_25976_, _25975_, _25974_);
  and (_25977_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_25978_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_25979_, _25978_, _25977_);
  or (_25980_, _25979_, _25976_);
  and (_25981_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and (_25982_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_25983_, _25982_, _25981_);
  and (_25984_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and (_25985_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_25986_, _25985_, _25984_);
  or (_25987_, _25986_, _25983_);
  or (_25988_, _25987_, _25980_);
  and (_25989_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_25990_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_25991_, _25990_, _25989_);
  and (_25992_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and (_25993_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_25994_, _25993_, _25992_);
  or (_25995_, _25994_, _25991_);
  and (_25996_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_25997_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_25998_, _25997_, _25996_);
  and (_25999_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  and (_26000_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_26001_, _26000_, _25999_);
  or (_26002_, _26001_, _25998_);
  or (_26003_, _26002_, _25995_);
  or (_26004_, _26003_, _25988_);
  or (_26005_, _26004_, _25973_);
  or (_26006_, _26005_, _25942_);
  and (_26007_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_26008_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_26009_, _26008_, _26007_);
  and (_26010_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_26011_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_26012_, _26011_, _26010_);
  or (_26013_, _26012_, _26009_);
  and (_26014_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_26015_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_26016_, _26015_, _26014_);
  and (_26017_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  and (_26018_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_26019_, _26018_, _26017_);
  or (_26020_, _26019_, _26016_);
  or (_26021_, _26020_, _26013_);
  and (_26022_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  and (_26023_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_26024_, _26023_, _26022_);
  and (_26025_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_26026_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or (_26027_, _26026_, _26025_);
  or (_26028_, _26027_, _26024_);
  and (_26029_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  and (_26030_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_26031_, _26030_, _26029_);
  and (_26032_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_26033_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_26034_, _26033_, _26032_);
  or (_26035_, _26034_, _26031_);
  or (_26036_, _26035_, _26028_);
  or (_26037_, _26036_, _26021_);
  and (_26038_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  and (_26039_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_26040_, _26039_, _26038_);
  and (_26041_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  and (_26042_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_26043_, _26042_, _26041_);
  or (_26044_, _26043_, _26040_);
  and (_26045_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  and (_26046_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_26047_, _26046_, _26045_);
  and (_26048_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_26049_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_26050_, _26049_, _26048_);
  or (_26051_, _26050_, _26047_);
  or (_26052_, _26051_, _26044_);
  and (_26053_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_26054_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_26055_, _26054_, _26053_);
  and (_26056_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  and (_26057_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_26058_, _26057_, _26056_);
  or (_26059_, _26058_, _26055_);
  and (_26060_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_26061_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_26062_, _26061_, _26060_);
  and (_26063_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  and (_26064_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_26065_, _26064_, _26063_);
  or (_26066_, _26065_, _26062_);
  or (_26067_, _26066_, _26059_);
  or (_26068_, _26067_, _26052_);
  or (_26069_, _26068_, _26037_);
  and (_26070_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_26071_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_26072_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_26073_, _26072_, _26071_);
  or (_26074_, _26073_, _26070_);
  and (_26075_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_26076_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_26077_, _26076_, _26075_);
  and (_26078_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_26079_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_26080_, _26079_, _26078_);
  or (_26081_, _26080_, _26077_);
  or (_26082_, _26081_, _26074_);
  and (_26083_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_26084_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_26085_, _26084_, _26083_);
  and (_26086_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_26087_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_26088_, _26087_, _26086_);
  or (_26089_, _26088_, _26085_);
  and (_26090_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_26091_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_26092_, _26091_, _26090_);
  and (_26093_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_26094_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_26095_, _26094_, _26093_);
  or (_26096_, _26095_, _26092_);
  or (_26097_, _26096_, _26089_);
  or (_26098_, _26097_, _26082_);
  and (_26099_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_26100_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_26101_, _26100_, _26099_);
  and (_26102_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  and (_26103_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_26104_, _26103_, _26102_);
  or (_26105_, _26104_, _26101_);
  and (_26106_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_26107_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_26108_, _26107_, _26106_);
  and (_26109_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_26110_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_26111_, _26110_, _26109_);
  or (_26112_, _26111_, _26108_);
  or (_26113_, _26112_, _26105_);
  and (_26114_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  and (_26115_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_26116_, _26115_, _26114_);
  and (_26117_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_26118_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_26119_, _26118_, _26117_);
  or (_26120_, _26119_, _26116_);
  and (_26121_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  and (_26122_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_26123_, _26122_, _26121_);
  and (_26124_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_26125_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_26126_, _26125_, _26124_);
  or (_26127_, _26126_, _26123_);
  or (_26128_, _26127_, _26120_);
  or (_26129_, _26128_, _26113_);
  or (_26130_, _26129_, _26098_);
  or (_26131_, _26130_, _26069_);
  or (_26132_, _26131_, _26006_);
  or (_26133_, _26132_, _25879_);
  and (_26134_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_26135_, _26134_, _26133_);
  and (_26136_, _26135_, _00006_);
  or (_26137_, _26136_, _25624_);
  and (_00003_[0], _26137_, _38997_);
  not (_26138_, first_instr);
  nor (_26139_, _15585_, _26138_);
  or (_00002_, _26139_, rst);
  and (_26140_, _15585_, iram_op1[7]);
  and (_26141_, _15589_, iram_op1_reg[7]);
  or (_26142_, _26141_, _26140_);
  and (_00004_[7], _26142_, _38997_);
  and (_26143_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_26144_, _21574_, acc_reg[7]);
  or (_26145_, _26144_, _26143_);
  and (_00000_[7], _26145_, _38997_);
  and (_26146_, pc_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_26147_, cy_reg, _21574_);
  or (_26148_, _26147_, _26146_);
  and (_00001_, _26148_, _38997_);
  and (_26149_, _18651_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26150_, _26149_, _21683_);
  nor (_26151_, _26150_, _16198_);
  nor (_26152_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26153_, _18646_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26154_, _26153_, _26152_);
  nor (_26155_, _26154_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_26156_, _26155_, _26151_);
  and (_26157_, _26156_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_26158_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_26159_, \oc8051_symbolic_cxrom1.regvalid [8], _16202_);
  nor (_26160_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26161_, _26160_, _26159_);
  and (_26162_, _26161_, _26158_);
  and (_26163_, _18663_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26164_, _26163_, _21675_);
  and (_26165_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], _16194_);
  and (_26166_, _26165_, _26164_);
  or (_26167_, _26166_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_26168_, _26167_, _26162_);
  nor (_26169_, _26168_, _26157_);
  and (_26170_, _18622_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_26171_, _26170_);
  nor (_26172_, _21670_, _16198_);
  and (_26173_, _26172_, _26171_);
  nor (_26174_, \oc8051_symbolic_cxrom1.regvalid [11], _16202_);
  nor (_26175_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26176_, _26175_, _26174_);
  and (_26177_, _26176_, _16198_);
  nor (_26178_, _26177_, _26173_);
  nor (_26179_, _26178_, _16194_);
  and (_26180_, _18885_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26181_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26182_, _26181_, _26180_);
  and (_26183_, _26182_, _26158_);
  and (_26184_, _18630_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26185_, _26184_, _21679_);
  and (_26186_, _26185_, _26165_);
  or (_26187_, _26186_, _16190_);
  or (_26188_, _26187_, _26183_);
  nor (_26189_, _26188_, _26179_);
  nor (_26190_, _26189_, _26169_);
  nor (_26191_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26192_, _20612_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26193_, _26192_, _26191_);
  and (_26194_, _26193_, _26165_);
  not (_26195_, _26194_);
  and (_26196_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_26197_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26198_, _19705_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26199_, _26198_, _26197_);
  and (_26200_, _26199_, _26196_);
  nor (_26201_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26202_, _20606_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26203_, _26202_, _26201_);
  and (_26204_, _26203_, _26158_);
  nor (_26205_, _26204_, _26200_);
  and (_26206_, _26205_, _26195_);
  nor (_26207_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26208_, _20621_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26209_, _26208_, _26207_);
  and (_26210_, _16198_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_26211_, _26210_, _26209_);
  nor (_26212_, _26211_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26213_, _26212_, _26206_);
  nor (_26214_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26215_, _20318_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26216_, _26215_, _26214_);
  and (_26217_, _26216_, _26165_);
  not (_26218_, _26217_);
  nor (_26219_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26220_, _20521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26221_, _26220_, _26219_);
  and (_26222_, _26221_, _26196_);
  nor (_26223_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26224_, _19913_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26225_, _26224_, _26223_);
  and (_26226_, _26225_, _26158_);
  nor (_26227_, _26226_, _26222_);
  and (_26228_, _26227_, _26218_);
  nor (_26229_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26230_, _20116_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26231_, _26230_, _26229_);
  and (_26232_, _26231_, _26210_);
  nor (_26233_, _26232_, _16202_);
  and (_26234_, _26233_, _26228_);
  nor (_26235_, _26234_, _26213_);
  and (_26236_, _26235_, _26190_);
  nor (_26237_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26238_, _20704_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26239_, _26238_, _26237_);
  and (_26240_, _26239_, _26165_);
  not (_26241_, _26240_);
  nor (_26242_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26243_, _19735_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26244_, _26243_, _26242_);
  and (_26245_, _26244_, _26196_);
  nor (_26246_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26247_, _20698_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26248_, _26247_, _26246_);
  and (_26249_, _26248_, _26158_);
  nor (_26250_, _26249_, _26245_);
  and (_26251_, _26250_, _26241_);
  nor (_26252_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26253_, _20713_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26254_, _26253_, _26252_);
  and (_26255_, _26254_, _26210_);
  nor (_26256_, _26255_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26257_, _26256_, _26251_);
  nor (_26258_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26259_, _20346_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26260_, _26259_, _26258_);
  and (_26261_, _26260_, _26165_);
  not (_26262_, _26261_);
  nor (_26263_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26264_, _20547_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26265_, _26264_, _26263_);
  and (_26266_, _26265_, _26196_);
  nor (_26267_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26268_, _19937_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26269_, _26268_, _26267_);
  and (_26270_, _26269_, _26158_);
  nor (_26271_, _26270_, _26266_);
  and (_26272_, _26271_, _26262_);
  nor (_26273_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26274_, _20142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26275_, _26274_, _26273_);
  and (_26276_, _26275_, _26210_);
  nor (_26277_, _26276_, _16202_);
  and (_26278_, _26277_, _26272_);
  nor (_26279_, _26278_, _26257_);
  and (_26280_, _26279_, _26190_);
  nor (_26281_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26282_, _20658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26283_, _26282_, _26281_);
  and (_26284_, _26283_, _26165_);
  not (_26285_, _26284_);
  nor (_26286_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26287_, _19721_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26288_, _26287_, _26286_);
  and (_26289_, _26288_, _26196_);
  nor (_26290_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26291_, _20652_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26292_, _26291_, _26290_);
  and (_26293_, _26292_, _26158_);
  nor (_26294_, _26293_, _26289_);
  and (_26295_, _26294_, _26285_);
  nor (_26296_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26297_, _20667_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26298_, _26297_, _26296_);
  and (_26299_, _26298_, _26210_);
  nor (_26300_, _26299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26301_, _26300_, _26295_);
  nor (_26302_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26303_, _20334_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26304_, _26303_, _26302_);
  and (_26305_, _26304_, _26165_);
  not (_26306_, _26305_);
  nor (_26307_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26308_, _20534_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26309_, _26308_, _26307_);
  and (_26310_, _26309_, _26196_);
  nor (_26311_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26312_, _19925_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26313_, _26312_, _26311_);
  and (_26314_, _26313_, _26158_);
  nor (_26315_, _26314_, _26310_);
  and (_26316_, _26315_, _26306_);
  nor (_26317_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26318_, _20127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26319_, _26318_, _26317_);
  and (_26320_, _26319_, _26210_);
  nor (_26321_, _26320_, _16202_);
  and (_26322_, _26321_, _26316_);
  nor (_26323_, _26322_, _26301_);
  nor (_26324_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26325_, _20750_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26326_, _26325_, _26324_);
  and (_26327_, _26326_, _26165_);
  not (_26328_, _26327_);
  nor (_26329_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26330_, _19745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26331_, _26330_, _26329_);
  and (_26332_, _26331_, _26196_);
  nor (_26333_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26334_, _20744_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26335_, _26334_, _26333_);
  and (_26336_, _26335_, _26158_);
  nor (_26337_, _26336_, _26332_);
  and (_26338_, _26337_, _26328_);
  nor (_26339_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26340_, _20759_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26341_, _26340_, _26339_);
  and (_26342_, _26341_, _26210_);
  nor (_26343_, _26342_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26344_, _26343_, _26338_);
  nor (_26345_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26346_, _20359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26347_, _26346_, _26345_);
  and (_26348_, _26347_, _26165_);
  not (_26349_, _26348_);
  nor (_26350_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26351_, _20559_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26352_, _26351_, _26350_);
  and (_26353_, _26352_, _26196_);
  nor (_26354_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26355_, _19951_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26356_, _26355_, _26354_);
  and (_26357_, _26356_, _26158_);
  nor (_26358_, _26357_, _26353_);
  and (_26359_, _26358_, _26349_);
  nor (_26360_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26361_, _20154_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26362_, _26361_, _26360_);
  and (_26363_, _26362_, _26210_);
  nor (_26364_, _26363_, _16202_);
  and (_26365_, _26364_, _26359_);
  nor (_26366_, _26365_, _26344_);
  nor (_26367_, _26366_, _26323_);
  and (_26368_, _26367_, _26280_);
  and (_26369_, _26368_, _26236_);
  nor (_26370_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26371_, _20888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26372_, _26371_, _26370_);
  and (_26373_, _26372_, _26165_);
  not (_26374_, _26373_);
  nor (_26375_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26376_, _19782_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26377_, _26376_, _26375_);
  and (_26378_, _26377_, _26196_);
  nor (_26379_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26380_, _20882_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26381_, _26380_, _26379_);
  and (_26382_, _26381_, _26158_);
  nor (_26383_, _26382_, _26378_);
  and (_26384_, _26383_, _26374_);
  nor (_26385_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26386_, _20897_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26387_, _26386_, _26385_);
  and (_26388_, _26387_, _26210_);
  nor (_26389_, _26388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26390_, _26389_, _26384_);
  nor (_26391_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26392_, _20395_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26393_, _26392_, _26391_);
  and (_26394_, _26393_, _26165_);
  not (_26395_, _26394_);
  nor (_26396_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26397_, _20593_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26398_, _26397_, _26396_);
  and (_26399_, _26398_, _26196_);
  nor (_26400_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26401_, _19988_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26402_, _26401_, _26400_);
  and (_26403_, _26402_, _26158_);
  nor (_26404_, _26403_, _26399_);
  and (_26405_, _26404_, _26395_);
  nor (_26406_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26407_, _20190_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26408_, _26407_, _26406_);
  and (_26409_, _26408_, _26210_);
  nor (_26410_, _26409_, _16202_);
  and (_26411_, _26410_, _26405_);
  nor (_26412_, _26411_, _26390_);
  and (_26413_, _26412_, _26190_);
  nor (_26414_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26415_, _18457_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26416_, _26415_, _26414_);
  and (_26417_, _26416_, _26165_);
  not (_26418_, _26417_);
  nor (_26419_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26420_, _18451_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26421_, _26420_, _26419_);
  and (_26422_, _26421_, _26196_);
  nor (_26423_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26424_, _18443_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26425_, _26424_, _26423_);
  and (_26426_, _26425_, _26158_);
  nor (_26427_, _26426_, _26422_);
  and (_26428_, _26427_, _26418_);
  nor (_26429_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26430_, _18462_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26431_, _26430_, _26429_);
  and (_26432_, _26431_, _26210_);
  nor (_26433_, _26432_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26434_, _26433_, _26428_);
  nor (_26435_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26436_, _18478_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26437_, _26436_, _26435_);
  and (_26438_, _26437_, _26165_);
  not (_26439_, _26438_);
  nor (_26440_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26441_, _18483_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26442_, _26441_, _26440_);
  and (_26443_, _26442_, _26196_);
  nor (_26444_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26445_, _18472_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26446_, _26445_, _26444_);
  and (_26447_, _26446_, _26158_);
  nor (_26448_, _26447_, _26443_);
  and (_26449_, _26448_, _26439_);
  nor (_26450_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26451_, _18489_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26452_, _26451_, _26450_);
  and (_26453_, _26452_, _26210_);
  nor (_26454_, _26453_, _16202_);
  and (_26455_, _26454_, _26449_);
  nor (_26456_, _26455_, _26434_);
  and (_26457_, _26456_, _26190_);
  nor (_26458_, _26457_, _26413_);
  nor (_26459_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26460_, _20796_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26461_, _26460_, _26459_);
  and (_26462_, _26461_, _26165_);
  not (_26463_, _26462_);
  nor (_26464_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26465_, _19759_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26466_, _26465_, _26464_);
  and (_26467_, _26466_, _26196_);
  nor (_26468_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26469_, _20790_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26470_, _26469_, _26468_);
  and (_26471_, _26470_, _26158_);
  nor (_26472_, _26471_, _26467_);
  and (_26473_, _26472_, _26463_);
  nor (_26474_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26475_, _20805_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26476_, _26475_, _26474_);
  and (_26477_, _26476_, _26210_);
  nor (_26478_, _26477_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26479_, _26478_, _26473_);
  nor (_26480_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26481_, _20372_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26482_, _26481_, _26480_);
  and (_26483_, _26482_, _26165_);
  not (_26484_, _26483_);
  nor (_26485_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26486_, _20571_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26487_, _26486_, _26485_);
  and (_26488_, _26487_, _26196_);
  nor (_26489_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26490_, _19963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26491_, _26490_, _26489_);
  and (_26492_, _26491_, _26158_);
  nor (_26493_, _26492_, _26488_);
  and (_26494_, _26493_, _26484_);
  nor (_26495_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26496_, _20165_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26497_, _26496_, _26495_);
  and (_26498_, _26497_, _26210_);
  nor (_26499_, _26498_, _16202_);
  and (_26500_, _26499_, _26494_);
  nor (_26501_, _26500_, _26479_);
  and (_26502_, _26501_, _26190_);
  nor (_26503_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26504_, _20842_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26505_, _26504_, _26503_);
  and (_26506_, _26505_, _26165_);
  not (_26507_, _26506_);
  nor (_26508_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26509_, _19770_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26510_, _26509_, _26508_);
  and (_26511_, _26510_, _26196_);
  nor (_26512_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26513_, _20836_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26514_, _26513_, _26512_);
  and (_26515_, _26514_, _26158_);
  nor (_26516_, _26515_, _26511_);
  and (_26517_, _26516_, _26507_);
  nor (_26518_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26519_, _20851_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26520_, _26519_, _26518_);
  and (_26521_, _26520_, _26210_);
  nor (_26522_, _26521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_26523_, _26522_, _26517_);
  nor (_26524_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26525_, _20382_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26526_, _26525_, _26524_);
  and (_26527_, _26526_, _26165_);
  not (_26528_, _26527_);
  nor (_26529_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26530_, _20584_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26531_, _26530_, _26529_);
  and (_26532_, _26531_, _26196_);
  nor (_26533_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26534_, _19975_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26535_, _26534_, _26533_);
  and (_26536_, _26535_, _26158_);
  nor (_26537_, _26536_, _26532_);
  and (_26538_, _26537_, _26528_);
  nor (_26539_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_26540_, _20178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_26541_, _26540_, _26539_);
  and (_26542_, _26541_, _26210_);
  nor (_26543_, _26542_, _16202_);
  and (_26544_, _26543_, _26538_);
  nor (_26545_, _26544_, _26523_);
  and (_26546_, _26545_, _26190_);
  nor (_26547_, _26546_, _26502_);
  and (_26548_, _26547_, _26458_);
  and (_26549_, _26548_, _38997_);
  and (_00008_, _26549_, _26369_);
  not (_26550_, _26236_);
  and (_26551_, _26368_, _26550_);
  and (_00007_, _26551_, _26549_);
  or (_26552_, _21983_, _15589_);
  or (_26553_, _15585_, op1_out_r[7]);
  and (_26554_, _26553_, _38997_);
  and (_00005_[7], _26554_, _26552_);
  and (_26555_, _15589_, iram_op1[7]);
  and (_26556_, _21989_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and (_26557_, _21994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_26558_, _26557_, _26556_);
  and (_26559_, _22006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_26560_, _21999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or (_26561_, _26560_, _26559_);
  or (_26562_, _26561_, _26558_);
  and (_26563_, _22013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and (_26564_, _22016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_26565_, _26564_, _26563_);
  and (_26566_, _22023_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_26567_, _22020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or (_26568_, _26567_, _26566_);
  or (_26569_, _26568_, _26565_);
  or (_26570_, _26569_, _26562_);
  and (_26571_, _22032_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_26572_, _22029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or (_26573_, _26572_, _26571_);
  and (_26574_, _22036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  and (_26575_, _22040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_26576_, _26575_, _26574_);
  or (_26577_, _26576_, _26573_);
  and (_26578_, _22048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_26579_, _22045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or (_26580_, _26579_, _26578_);
  and (_26581_, _22052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  and (_26582_, _22055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or (_26583_, _26582_, _26581_);
  or (_26584_, _26583_, _26580_);
  or (_26585_, _26584_, _26577_);
  or (_26586_, _26585_, _26570_);
  and (_26587_, _22061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_26588_, _22063_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_26589_, _26588_, _26587_);
  and (_26590_, _22068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and (_26591_, _22070_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_26592_, _26591_, _26590_);
  or (_26593_, _26592_, _26589_);
  and (_26594_, _22074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_26595_, _22076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or (_26596_, _26595_, _26594_);
  and (_26597_, _22079_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  and (_26598_, _22081_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_26599_, _26598_, _26597_);
  or (_26600_, _26599_, _26596_);
  or (_26601_, _26600_, _26593_);
  and (_26602_, _22088_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  and (_26603_, _22086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_26604_, _26603_, _26602_);
  and (_26605_, _22091_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_26606_, _22093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_26607_, _26606_, _26605_);
  or (_26608_, _26607_, _26604_);
  and (_26609_, _22097_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  and (_26610_, _22099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_26611_, _26610_, _26609_);
  and (_26612_, _22104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  and (_26613_, _22102_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_26614_, _26613_, _26612_);
  or (_26615_, _26614_, _26611_);
  or (_26616_, _26615_, _26608_);
  or (_26617_, _26616_, _26601_);
  or (_26618_, _26617_, _26586_);
  and (_26619_, _22185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_26620_, _22183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_26621_, _26620_, _26619_);
  and (_26622_, _22188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  and (_26623_, _22190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_26624_, _26623_, _26622_);
  or (_26625_, _26624_, _26621_);
  and (_26626_, _22196_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_26627_, _22194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_26628_, _26627_, _26626_);
  and (_26629_, _22204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and (_26630_, _22202_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_26631_, _26630_, _26629_);
  or (_26632_, _26631_, _26628_);
  or (_26633_, _26632_, _26625_);
  and (_26634_, _22173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and (_26635_, _22171_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_26636_, _26635_, _26634_);
  and (_26637_, _22178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and (_26638_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_26639_, _26638_, _26637_);
  or (_26640_, _26639_, _26636_);
  and (_26641_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and (_26642_, _22160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_26643_, _26642_, _26641_);
  and (_26644_, _22165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_26645_, _22167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_26646_, _26645_, _26644_);
  or (_26647_, _26646_, _26643_);
  or (_26648_, _26647_, _26640_);
  or (_26649_, _26648_, _26633_);
  and (_26650_, _22113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_26651_, _22111_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  or (_26652_, _26651_, _26650_);
  and (_26653_, _22116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and (_26654_, _22118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_26655_, _26654_, _26653_);
  or (_26656_, _26655_, _26652_);
  and (_26657_, _22122_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_26658_, _22124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  or (_26659_, _26658_, _26657_);
  and (_26660_, _22129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_26661_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_26662_, _26661_, _26660_);
  or (_26663_, _26662_, _26659_);
  or (_26664_, _26663_, _26656_);
  and (_26665_, _22149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and (_26666_, _22147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_26667_, _26666_, _26665_);
  and (_26668_, _22154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_26669_, _22152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or (_26670_, _26669_, _26668_);
  or (_26671_, _26670_, _26667_);
  and (_26672_, _22136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and (_26673_, _22134_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_26674_, _26673_, _26672_);
  and (_26675_, _22143_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_26676_, _22141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_26677_, _26676_, _26675_);
  or (_26678_, _26677_, _26674_);
  or (_26679_, _26678_, _26671_);
  or (_26680_, _26679_, _26664_);
  or (_26681_, _26680_, _26649_);
  or (_26682_, _26681_, _26618_);
  and (_26683_, _22212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  and (_26684_, _22214_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_26685_, _26684_, _26683_);
  and (_26686_, _22217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_26687_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_26688_, _26687_, _26686_);
  or (_26689_, _26688_, _26685_);
  and (_26690_, _22223_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  and (_26691_, _22225_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_26692_, _26691_, _26690_);
  and (_26693_, _22229_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_26694_, _22231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or (_26695_, _26694_, _26693_);
  or (_26696_, _26695_, _26692_);
  or (_26697_, _26696_, _26689_);
  and (_26698_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_26699_, _22236_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_26700_, _26699_, _26698_);
  and (_26701_, _22241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  and (_26702_, _22243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_26703_, _26702_, _26701_);
  or (_26704_, _26703_, _26700_);
  and (_26705_, _22247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_26706_, _22249_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_26707_, _26706_, _26705_);
  and (_26708_, _22252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  and (_26709_, _22254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_26710_, _26709_, _26708_);
  or (_26711_, _26710_, _26707_);
  or (_26712_, _26711_, _26704_);
  or (_26713_, _26712_, _26697_);
  and (_26714_, _22273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_26715_, _22271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_26716_, _26715_, _26714_);
  and (_26717_, _22276_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_26718_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or (_26719_, _26718_, _26717_);
  or (_26720_, _26719_, _26716_);
  and (_26721_, _22260_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_26722_, _22262_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_26723_, _26722_, _26721_);
  and (_26724_, _22267_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_26725_, _22265_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_26726_, _26725_, _26724_);
  or (_26727_, _26726_, _26723_);
  or (_26728_, _26727_, _26720_);
  and (_26729_, _22283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_26730_, _22285_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  or (_26731_, _26730_, _26729_);
  and (_26732_, _22290_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and (_26733_, _22288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_26734_, _26733_, _26732_);
  or (_26735_, _26734_, _26731_);
  and (_26736_, _22296_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_26737_, _22294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  or (_26738_, _26737_, _26736_);
  and (_26739_, _22302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and (_26740_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_26741_, _26740_, _26739_);
  or (_26742_, _26741_, _26738_);
  or (_26743_, _26742_, _26735_);
  or (_26744_, _26743_, _26728_);
  or (_26745_, _26744_, _26713_);
  and (_26746_, _22333_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_26747_, _22335_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or (_26748_, _26747_, _26746_);
  and (_26749_, _22338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and (_26750_, _22340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_26751_, _26750_, _26749_);
  or (_26752_, _26751_, _26748_);
  and (_26753_, _22346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_26754_, _22344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or (_26755_, _26754_, _26753_);
  and (_26756_, _22351_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_26757_, _22349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_26758_, _26757_, _26756_);
  or (_26759_, _26758_, _26755_);
  or (_26760_, _26759_, _26752_);
  and (_26761_, _22321_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and (_26762_, _22323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_26763_, _26762_, _26761_);
  and (_26764_, _22328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_26765_, _22326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or (_26766_, _26765_, _26764_);
  or (_26767_, _26766_, _26763_);
  and (_26768_, _22317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_26769_, _22314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or (_26770_, _26769_, _26768_);
  and (_26771_, _22311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and (_26772_, _22309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_26773_, _26772_, _26771_);
  or (_26774_, _26773_, _26770_);
  or (_26775_, _26774_, _26767_);
  or (_26776_, _26775_, _26760_);
  and (_26777_, _22382_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and (_26778_, _22384_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_26779_, _26778_, _26777_);
  and (_26780_, _22389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_26781_, _22387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_26782_, _26781_, _26780_);
  or (_26783_, _26782_, _26779_);
  and (_26784_, _22393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and (_26785_, _22395_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_26786_, _26785_, _26784_);
  and (_26787_, _22398_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and (_26788_, _22400_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_26789_, _26788_, _26787_);
  or (_26790_, _26789_, _26786_);
  or (_26791_, _26790_, _26783_);
  and (_26792_, _22359_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_26793_, _22357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_26794_, _26793_, _26792_);
  and (_26795_, _22366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  and (_26796_, _22362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_26797_, _26796_, _26795_);
  or (_26798_, _26797_, _26794_);
  and (_26799_, _22370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_26800_, _22372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_26801_, _26800_, _26799_);
  and (_26802_, _22375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  and (_26803_, _22377_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_26804_, _26803_, _26802_);
  or (_26805_, _26804_, _26801_);
  or (_26806_, _26805_, _26798_);
  or (_26807_, _26806_, _26791_);
  or (_26808_, _26807_, _26776_);
  or (_26809_, _26808_, _26745_);
  or (_26810_, _26809_, _26682_);
  and (_26811_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_26812_, _22444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_26813_, _26812_, _26811_);
  and (_26814_, _22451_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  and (_26815_, _22449_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_26816_, _26815_, _26814_);
  or (_26817_, _26816_, _26813_);
  and (_26818_, _22433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_26819_, _22435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or (_26820_, _26819_, _26818_);
  and (_26821_, _22438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_26822_, _22440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_26823_, _26822_, _26821_);
  or (_26824_, _26823_, _26820_);
  or (_26825_, _26824_, _26817_);
  and (_26826_, _22420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  and (_26827_, _22422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_26828_, _26827_, _26826_);
  and (_26829_, _22426_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_26830_, _22428_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or (_26831_, _26830_, _26829_);
  or (_26832_, _26831_, _26828_);
  and (_26833_, _22409_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  and (_26834_, _22411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_26835_, _26834_, _26833_);
  and (_26836_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_26837_, _22414_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_26838_, _26837_, _26836_);
  or (_26839_, _26838_, _26835_);
  or (_26840_, _26839_, _26832_);
  or (_26841_, _26840_, _26825_);
  and (_26842_, _22457_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  and (_26843_, _22459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_26844_, _26843_, _26842_);
  and (_26845_, _22464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_26846_, _22462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_26847_, _26846_, _26845_);
  or (_26848_, _26847_, _26844_);
  and (_26849_, _22468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  and (_26850_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_26851_, _26850_, _26849_);
  and (_26852_, _22475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  and (_26853_, _22473_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_26854_, _26853_, _26852_);
  or (_26855_, _26854_, _26851_);
  or (_26856_, _26855_, _26848_);
  and (_26857_, _22491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_26858_, _22493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_26859_, _26858_, _26857_);
  and (_26860_, _22499_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  and (_26861_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_26862_, _26861_, _26860_);
  or (_26863_, _26862_, _26859_);
  and (_26864_, _22482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_26865_, _22480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_26866_, _26865_, _26864_);
  and (_26867_, _22487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  and (_26868_, _22485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_26869_, _26868_, _26867_);
  or (_26870_, _26869_, _26866_);
  or (_26871_, _26870_, _26863_);
  or (_26872_, _26871_, _26856_);
  or (_26873_, _26872_, _26841_);
  and (_26874_, _22519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  and (_26875_, _22517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_26876_, _26875_, _26874_);
  and (_26877_, _22525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_26878_, _22522_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_26879_, _26878_, _26877_);
  or (_26880_, _26879_, _26876_);
  and (_26881_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  and (_26882_, _22508_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_26883_, _26882_, _26881_);
  and (_26884_, _22511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_26885_, _22513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_26886_, _26885_, _26884_);
  or (_26887_, _26886_, _26883_);
  or (_26888_, _26887_, _26880_);
  and (_26889_, _22546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_26890_, _22548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_26891_, _26890_, _26889_);
  and (_26892_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  and (_26893_, _22541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_26894_, _26893_, _26892_);
  or (_26895_, _26894_, _26891_);
  and (_26896_, _22532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_26897_, _22530_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_26898_, _26897_, _26896_);
  and (_26899_, _22537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  and (_26900_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_26901_, _26900_, _26899_);
  or (_26902_, _26901_, _26898_);
  or (_26903_, _26902_, _26895_);
  or (_26904_, _26903_, _26888_);
  and (_26905_, _22556_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_26906_, _22554_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_26907_, _26906_, _26905_);
  and (_26908_, _22563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and (_26909_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_26910_, _26909_, _26908_);
  or (_26911_, _26910_, _26907_);
  and (_26912_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_26913_, _22569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_26914_, _26913_, _26912_);
  and (_26915_, _22572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  and (_26916_, _22574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_26917_, _26916_, _26915_);
  or (_26918_, _26917_, _26914_);
  or (_26919_, _26918_, _26911_);
  and (_26920_, _22581_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and (_26921_, _22579_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_26922_, _26921_, _26920_);
  and (_26923_, _22586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_26924_, _22584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_26925_, _26924_, _26923_);
  or (_26926_, _26925_, _26922_);
  and (_26927_, _22590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and (_26928_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_26929_, _26928_, _26927_);
  and (_26930_, _22595_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_26931_, _22597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_26932_, _26931_, _26930_);
  or (_26933_, _26932_, _26929_);
  or (_26934_, _26933_, _26926_);
  or (_26935_, _26934_, _26919_);
  or (_26936_, _26935_, _26904_);
  or (_26937_, _26936_, _26873_);
  and (_26938_, _22605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_26939_, _22607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_26940_, _26939_, _26938_);
  and (_26941_, _22612_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  and (_26942_, _22610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_26943_, _26942_, _26941_);
  or (_26944_, _26943_, _26940_);
  and (_26945_, _22618_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_26946_, _22616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_26947_, _26946_, _26945_);
  and (_26948_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  and (_26949_, _22621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_26950_, _26949_, _26948_);
  or (_26951_, _26950_, _26947_);
  or (_26952_, _26951_, _26944_);
  and (_26953_, _22630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  and (_26954_, _22628_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_26955_, _26954_, _26953_);
  and (_26956_, _22635_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_26957_, _22633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_26958_, _26957_, _26956_);
  or (_26959_, _26958_, _26955_);
  and (_26960_, _22644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_26961_, _22647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_26962_, _26961_, _26960_);
  and (_26963_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  and (_26964_, _22641_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_26965_, _26964_, _26963_);
  or (_26966_, _26965_, _26962_);
  or (_26967_, _26966_, _26959_);
  or (_26968_, _26967_, _26952_);
  and (_26969_, _22664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  and (_26970_, _22666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_26971_, _26970_, _26969_);
  and (_26972_, _22669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_26973_, _22671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_26974_, _26973_, _26972_);
  or (_26975_, _26974_, _26971_);
  and (_26976_, _22655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  and (_26977_, _22653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_26978_, _26977_, _26976_);
  and (_26979_, _22660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_26980_, _22658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_26981_, _26980_, _26979_);
  or (_26982_, _26981_, _26978_);
  or (_26983_, _26982_, _26975_);
  and (_26984_, _22681_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  and (_26985_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_26986_, _26985_, _26984_);
  and (_26987_, _22676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_26988_, _22678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_26989_, _26988_, _26987_);
  or (_26990_, _26989_, _26986_);
  and (_26991_, _22689_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_26992_, _22687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_26993_, _26992_, _26991_);
  and (_26994_, _22695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  and (_26995_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_26996_, _26995_, _26994_);
  or (_26997_, _26996_, _26993_);
  or (_26998_, _26997_, _26990_);
  or (_26999_, _26998_, _26983_);
  or (_27000_, _26999_, _26968_);
  and (_27001_, _22770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  and (_27002_, _22772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_27003_, _27002_, _27001_);
  and (_27004_, _22775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_27005_, _22777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_27006_, _27005_, _27004_);
  or (_27007_, _27006_, _27003_);
  and (_27008_, _22786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  and (_27009_, _22788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_27010_, _27009_, _27008_);
  and (_27011_, _22783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_27012_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_27013_, _27012_, _27011_);
  or (_27014_, _27013_, _27010_);
  or (_27015_, _27014_, _27007_);
  and (_27016_, _22760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_27017_, _22758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_27018_, _27017_, _27016_);
  and (_27019_, _22765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_27020_, _22763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_27021_, _27020_, _27019_);
  or (_27022_, _27021_, _27018_);
  and (_27023_, _22747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_27024_, _22749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_27025_, _27024_, _27023_);
  and (_27026_, _22752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  and (_27027_, _22754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_27028_, _27027_, _27026_);
  or (_27029_, _27028_, _27025_);
  or (_27030_, _27029_, _27022_);
  or (_27031_, _27030_, _27015_);
  and (_27032_, _22708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_27033_, _22716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_27034_, _22711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_27035_, _22713_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_27036_, _27035_, _27034_);
  or (_27037_, _27036_, _27033_);
  or (_27038_, _27037_, _27032_);
  and (_27039_, _22718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_27040_, _22703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_27041_, _22705_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_27042_, _27041_, _27040_);
  or (_27043_, _27042_, _27039_);
  or (_27044_, _27043_, _27038_);
  and (_27045_, _22723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_27046_, _22725_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_27047_, _27046_, _27045_);
  and (_27048_, _22728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_27049_, _22730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_27050_, _27049_, _27048_);
  or (_27051_, _27050_, _27047_);
  and (_27052_, _22736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_27053_, _22734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_27054_, _27053_, _27052_);
  and (_27055_, _22741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_27056_, _22739_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_27057_, _27056_, _27055_);
  or (_27058_, _27057_, _27054_);
  or (_27059_, _27058_, _27051_);
  or (_27060_, _27059_, _27044_);
  or (_27061_, _27060_, _27031_);
  or (_27062_, _27061_, _27000_);
  or (_27063_, _27062_, _26937_);
  or (_27064_, _27063_, _26810_);
  and (_27065_, _23049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_27066_, _27065_, _27064_);
  and (_27067_, _27066_, _00006_);
  or (_27068_, _27067_, _26555_);
  and (_00003_[7], _27068_, _38997_);
  and (_27069_, _26196_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_27070_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_27071_, _27070_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_27072_, _27071_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_27073_, _27072_, _27069_);
  and (_27074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_27075_, _27074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_27076_, _27075_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_27077_, _27076_, _27073_);
  and (_27078_, _27077_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_27079_, _27078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_27080_, _27079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_27081_, _27079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_27082_, _27081_, _27080_);
  and (_27083_, _27082_, _21983_);
  nor (_27084_, _27078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_27085_, _27084_, _27079_);
  and (_27086_, _27085_, _21983_);
  nor (_27087_, _27077_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_27088_, _27087_, _27078_);
  and (_27089_, _27088_, _21983_);
  nor (_27090_, _27085_, _21983_);
  nor (_27091_, _27090_, _27086_);
  and (_27092_, _27075_, _27073_);
  nor (_27093_, _27092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_27094_, _27092_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_27095_, _27094_, _27093_);
  and (_27096_, _27095_, _21983_);
  nor (_27097_, _27095_, _21983_);
  and (_27098_, _27073_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_27099_, _27098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_27100_, _27099_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_27101_, _27100_, _27092_);
  and (_27102_, _27101_, _21983_);
  nor (_27103_, _27101_, _21983_);
  nor (_27104_, _27103_, _27102_);
  not (_27105_, _27104_);
  nor (_27106_, _27098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_27107_, _27106_, _27099_);
  and (_27108_, _27107_, _21983_);
  nor (_27109_, _27073_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_27110_, _27109_, _27098_);
  and (_27111_, _27110_, _21983_);
  nor (_27112_, _27107_, _21983_);
  nor (_27113_, _27112_, _27108_);
  and (_27114_, _27071_, _27069_);
  nor (_27115_, _27114_, _16218_);
  and (_27116_, _27114_, _16218_);
  nor (_27117_, _27116_, _27115_);
  not (_27118_, _27117_);
  and (_27119_, _27118_, _21983_);
  nor (_27120_, _27118_, _21983_);
  and (_27121_, _27070_, _27069_);
  nor (_27122_, _27121_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_27123_, _27122_, _27114_);
  and (_27124_, _27123_, _21690_);
  nor (_27125_, _27123_, _21690_);
  nor (_27126_, _27125_, _27124_);
  not (_27127_, _27126_);
  and (_27128_, _27069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_27129_, _27128_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_27130_, _27129_, _27121_);
  and (_27131_, _27130_, _21732_);
  nor (_27132_, _27130_, _21732_);
  nor (_27133_, _27132_, _27131_);
  not (_27134_, _27133_);
  nor (_27135_, _27069_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_27136_, _27135_, _27128_);
  and (_27137_, _27136_, _21774_);
  nor (_27138_, _26196_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_27139_, _27138_, _27069_);
  not (_27140_, _27139_);
  and (_27141_, _21816_, _27140_);
  nor (_27142_, _21816_, _27140_);
  nor (_27143_, _27142_, _27141_);
  not (_27144_, _27143_);
  nor (_27145_, _26210_, _26165_);
  not (_27146_, _27145_);
  and (_27147_, _27146_, _21857_);
  and (_27148_, _21898_, _16194_);
  and (_27149_, _21940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_27150_, _21898_, _16194_);
  nor (_27151_, _27150_, _27148_);
  and (_27152_, _27151_, _27149_);
  nor (_27153_, _27152_, _27148_);
  nor (_27154_, _27146_, _21857_);
  nor (_27155_, _27154_, _27147_);
  not (_27156_, _27155_);
  nor (_27157_, _27156_, _27153_);
  nor (_27158_, _27157_, _27147_);
  nor (_27159_, _27158_, _27144_);
  nor (_27160_, _27159_, _27141_);
  nor (_27161_, _27136_, _21774_);
  nor (_27162_, _27161_, _27137_);
  not (_27163_, _27162_);
  nor (_27164_, _27163_, _27160_);
  nor (_27165_, _27164_, _27137_);
  nor (_27166_, _27165_, _27134_);
  nor (_27167_, _27166_, _27131_);
  nor (_27168_, _27167_, _27127_);
  nor (_27169_, _27168_, _27124_);
  nor (_27170_, _27169_, _27120_);
  or (_27171_, _27170_, _27119_);
  nor (_27172_, _27110_, _21983_);
  nor (_27173_, _27172_, _27111_);
  and (_27174_, _27173_, _27171_);
  and (_27175_, _27174_, _27113_);
  or (_27176_, _27175_, _27111_);
  nor (_27177_, _27176_, _27108_);
  nor (_27178_, _27177_, _27105_);
  nor (_27179_, _27178_, _27102_);
  nor (_27180_, _27179_, _27097_);
  nor (_27181_, _27180_, _27096_);
  nor (_27182_, _27088_, _21983_);
  nor (_27183_, _27182_, _27089_);
  not (_27184_, _27183_);
  nor (_27185_, _27184_, _27181_);
  and (_27186_, _27185_, _27091_);
  or (_27187_, _27186_, _27089_);
  nor (_27188_, _27187_, _27086_);
  nor (_27189_, _27082_, _21983_);
  nor (_27190_, _27189_, _27083_);
  not (_27191_, _27190_);
  nor (_27192_, _27191_, _27188_);
  nor (_27193_, _27192_, _27083_);
  nor (_27194_, _27080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_27195_, _27080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_27196_, _27195_, _27194_);
  not (_27197_, _27196_);
  and (_27198_, _27197_, _21983_);
  nor (_27199_, _27197_, _21983_);
  nor (_27200_, _27199_, _27198_);
  and (_27201_, _27200_, _27193_);
  nor (_27202_, _27200_, _27193_);
  or (_27203_, _27202_, _27201_);
  nor (_27204_, _27203_, cy_reg);
  and (_27205_, _27196_, cy_reg);
  nor (_27206_, _27205_, _27204_);
  nand (_27207_, _27206_, _14142_);
  or (_27208_, _27206_, _14142_);
  and (_27209_, _27208_, _27207_);
  not (_27210_, cy_reg);
  nor (_27211_, _27185_, _27089_);
  and (_27212_, _27211_, _27091_);
  nor (_27213_, _27211_, _27091_);
  nor (_27214_, _27213_, _27212_);
  and (_27215_, _27214_, _27210_);
  nor (_27216_, _27085_, _27210_);
  nor (_27217_, _27216_, _27215_);
  nand (_27218_, _27217_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_27219_, _27217_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_27220_, _27219_, _27218_);
  and (_27221_, _27184_, _27181_);
  nor (_27222_, _27221_, _27185_);
  nor (_27223_, _27222_, cy_reg);
  nor (_27224_, _27088_, _27210_);
  nor (_27225_, _27224_, _27223_);
  nand (_27226_, _27225_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_27227_, _27225_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_27228_, _27227_, _27226_);
  and (_27229_, _27177_, _27105_);
  nor (_27230_, _27229_, _27178_);
  or (_27231_, _27230_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_27232_, _27230_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_27233_, _27232_, _27231_);
  nor (_27234_, _27097_, _27096_);
  nor (_27235_, _27234_, _27179_);
  and (_27236_, _27234_, _27179_);
  nor (_27237_, _27236_, _27235_);
  or (_27238_, _27237_, _14106_);
  nand (_27239_, _27237_, _14106_);
  and (_27240_, _27239_, _27238_);
  or (_27241_, _27240_, _27233_);
  or (_27242_, _27241_, cy_reg);
  nor (_27243_, _27101_, _14121_);
  and (_27244_, _27101_, _14121_);
  or (_27245_, _27244_, _27243_);
  nor (_27246_, _27095_, _14106_);
  and (_27247_, _27095_, _14106_);
  or (_27248_, _27247_, _27246_);
  or (_27249_, _27248_, _27210_);
  or (_27250_, _27249_, _27245_);
  and (_27251_, _27250_, _27242_);
  nor (_27252_, _27174_, _27111_);
  and (_27253_, _27252_, _27113_);
  nor (_27254_, _27252_, _27113_);
  nor (_27255_, _27254_, _27253_);
  nor (_27256_, _27255_, cy_reg);
  and (_27257_, _27107_, cy_reg);
  nor (_27258_, _27257_, _27256_);
  nor (_27259_, _27258_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_27260_, _27258_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_27261_, _27110_, cy_reg);
  nor (_27262_, _27173_, _27171_);
  nor (_27263_, _27262_, _27174_);
  and (_27264_, _27263_, _27210_);
  nor (_27265_, _27264_, _27261_);
  and (_27266_, _27265_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_27267_, _27265_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_27268_, _27117_, _27210_);
  nor (_27269_, _27119_, _27120_);
  nor (_27270_, _27269_, _27169_);
  and (_27271_, _27269_, _27169_);
  or (_27272_, _27271_, _27270_);
  and (_27273_, _27272_, _27210_);
  nor (_27274_, _27273_, _27268_);
  and (_27275_, _27274_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_27276_, _27274_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_27277_, _27123_, cy_reg);
  and (_27278_, _27167_, _27127_);
  nor (_27279_, _27278_, _27168_);
  and (_27280_, _27279_, _27210_);
  nor (_27281_, _27280_, _27277_);
  and (_27282_, _27281_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_27283_, _27281_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_27284_, _27165_, _27134_);
  nor (_27285_, _27284_, _27166_);
  and (_27286_, _27285_, _27210_);
  and (_27287_, _27130_, cy_reg);
  nor (_27288_, _27287_, _27286_);
  and (_27289_, _27288_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_27290_, _27288_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_27291_, _27136_, cy_reg);
  and (_27292_, _27163_, _27160_);
  nor (_27293_, _27292_, _27164_);
  and (_27294_, _27293_, _27210_);
  nor (_27295_, _27294_, _27291_);
  and (_27296_, _27295_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_27297_, _27158_, _27144_);
  nor (_27298_, _27297_, _27159_);
  and (_27299_, _27298_, _27210_);
  nor (_27300_, _27139_, _27210_);
  nor (_27301_, _27300_, _27299_);
  and (_27302_, _27301_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_27303_, _27301_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27304_, _27156_, _27153_);
  nor (_27305_, _27304_, _27157_);
  and (_27306_, _27305_, _27210_);
  nor (_27307_, _27145_, _27210_);
  nor (_27308_, _27307_, _27306_);
  and (_27309_, _27308_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27310_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_27311_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_27312_, _27311_, _27310_);
  not (_27313_, _27312_);
  and (_27314_, _21940_, _27210_);
  nand (_27315_, _27314_, _27313_);
  or (_27316_, _27314_, _27313_);
  and (_27317_, _27316_, _27315_);
  and (_27318_, cy_reg, _16194_);
  nor (_27319_, _27151_, _27149_);
  nor (_27320_, _27319_, _27152_);
  and (_27321_, _27320_, _27210_);
  nor (_27322_, _27321_, _27318_);
  nor (_27323_, _27322_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27324_, _27322_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_27325_, _27324_, _27323_);
  or (_27326_, _27325_, _27317_);
  nor (_27327_, _27308_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_27328_, _27327_, _27326_);
  or (_27329_, _27328_, _27309_);
  or (_27330_, _27329_, _27303_);
  or (_27331_, _27330_, _27302_);
  nor (_27332_, _27295_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_27333_, _27332_, _27331_);
  or (_27334_, _27333_, _27296_);
  or (_27335_, _27334_, _27290_);
  or (_27336_, _27335_, _27289_);
  or (_27337_, _27336_, _27283_);
  or (_27338_, _27337_, _27282_);
  or (_27339_, _27338_, _27276_);
  or (_27340_, _27339_, _27275_);
  or (_27341_, _27340_, _27267_);
  or (_27342_, _27341_, _27266_);
  or (_27343_, _27342_, _27260_);
  or (_27344_, _27343_, _27259_);
  or (_27345_, _27344_, _27251_);
  or (_27346_, _27345_, _27228_);
  or (_27347_, _27346_, _27220_);
  and (_27348_, _27191_, _27188_);
  nor (_27349_, _27348_, _27192_);
  nor (_27350_, _27349_, cy_reg);
  nor (_27351_, _27082_, _27210_);
  nor (_27352_, _27351_, _27350_);
  and (_27353_, _27352_, _14137_);
  nor (_27354_, _27352_, _14137_);
  or (_27355_, _27354_, _27353_);
  or (_27356_, _27355_, _27347_);
  or (_27357_, _27356_, _27209_);
  and (_27358_, _26323_, _26190_);
  nor (_27359_, _27358_, _26236_);
  and (_27360_, _26366_, _26190_);
  nor (_27361_, _27360_, _26280_);
  and (_27362_, _27361_, _27359_);
  not (_27363_, _26545_);
  and (_27364_, _27363_, _26502_);
  and (_27365_, _27364_, _27362_);
  not (_27366_, _26457_);
  and (_27367_, _27366_, _26413_);
  or (_27368_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_27369_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27370_, \oc8051_symbolic_cxrom1.regvalid [1], _27369_);
  and (_27371_, _27370_, _15852_);
  and (_27372_, _27371_, _27368_);
  or (_27373_, \oc8051_symbolic_cxrom1.regvalid [13], _27369_);
  or (_27374_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27375_, _27374_, _27373_);
  not (_27376_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27377_, _27376_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27378_, _27377_, _27375_);
  or (_27379_, _27378_, _27372_);
  not (_27380_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_27381_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_27382_, _27381_, _27376_);
  nor (_27383_, _27382_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27384_, _27382_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_27385_, _27384_, _27383_);
  and (_27386_, _27385_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_27387_, _27381_, _27376_);
  nor (_27388_, _27387_, _27382_);
  nand (_27389_, \oc8051_symbolic_cxrom1.regvalid [7], _27369_);
  nand (_27390_, _27389_, _27388_);
  or (_27391_, _27390_, _27386_);
  and (_27392_, _27391_, _27380_);
  nor (_27393_, _27385_, _18609_);
  and (_27394_, _27385_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_27395_, _27394_, _27393_);
  or (_27396_, _27388_, _27395_);
  and (_27397_, _27396_, _27392_);
  or (_27398_, _27397_, _27379_);
  and (_27399_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27400_, \oc8051_symbolic_cxrom1.regvalid [0], _27369_);
  or (_27401_, _27400_, _27399_);
  and (_27402_, _27401_, _27376_);
  and (_27403_, \oc8051_symbolic_cxrom1.regvalid [4], _27369_);
  and (_27404_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27405_, _27404_, _27403_);
  and (_27406_, _27405_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_27407_, _27406_, _27402_);
  and (_27408_, _27407_, _27380_);
  and (_27409_, _15852_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_27410_, _27409_, _27369_);
  and (_27411_, _27409_, _27369_);
  nor (_27412_, _27411_, _27410_);
  nand (_27413_, _27412_, _18508_);
  and (_27414_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_27415_, _27414_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_27416_, _27415_, _27409_);
  and (_27417_, _27416_, _27373_);
  and (_27418_, _27417_, _27413_);
  or (_27419_, _27412_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not (_27420_, _27416_);
  nand (_27421_, _27412_, _18635_);
  and (_27422_, _27421_, _27420_);
  and (_27423_, _27422_, _27419_);
  or (_27424_, _27423_, _27418_);
  and (_27425_, _27424_, _27408_);
  not (_27426_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_27427_, _27412_, _27426_);
  or (_27428_, \oc8051_symbolic_cxrom1.regvalid [15], _27369_);
  and (_27429_, _27428_, _27416_);
  and (_27430_, _27429_, _27427_);
  or (_27431_, _27412_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand (_27432_, _27412_, _18609_);
  and (_27433_, _27432_, _27420_);
  and (_27434_, _27433_, _27431_);
  or (_27435_, _27434_, _27430_);
  and (_27436_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27437_, \oc8051_symbolic_cxrom1.regvalid [6], _27369_);
  or (_27438_, _27437_, _27376_);
  or (_27439_, _27438_, _27436_);
  or (_27440_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27441_, \oc8051_symbolic_cxrom1.regvalid [10], _27369_);
  and (_27442_, _27441_, _27440_);
  or (_27443_, _27442_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27444_, _27443_, _27439_);
  and (_27445_, _27444_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27446_, _27405_, _27377_);
  or (_27447_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27448_, \oc8051_symbolic_cxrom1.regvalid [0], _27369_);
  and (_27449_, _27448_, _15852_);
  and (_27450_, _27449_, _27447_);
  or (_27451_, _27450_, _27446_);
  and (_27452_, _27451_, _27445_);
  and (_27453_, _27452_, _27435_);
  or (_27454_, _27453_, _27425_);
  not (_27455_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_27456_, _27451_, _27444_);
  and (_27457_, _27456_, _27455_);
  and (_27458_, _27457_, _27454_);
  and (_27459_, _27458_, _27398_);
  or (_27460_, \oc8051_symbolic_cxrom1.regvalid [2], _27380_);
  or (_27461_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27462_, _27461_, _27460_);
  or (_27463_, _27462_, _27385_);
  or (_27464_, \oc8051_symbolic_cxrom1.regvalid [10], _27380_);
  or (_27465_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_27466_, _27465_, _27464_);
  and (_27467_, _27466_, _27385_);
  nor (_27468_, _27467_, _27388_);
  and (_27469_, _27468_, _27463_);
  and (_27470_, _27385_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_27471_, _27403_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_27472_, _27471_, _27470_);
  and (_27473_, _27385_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_27474_, _27437_, _27380_);
  or (_27475_, _27474_, _27473_);
  and (_27476_, _27475_, _27388_);
  and (_27477_, _27476_, _27472_);
  or (_27478_, _27477_, _27469_);
  nand (_27479_, _27412_, _18543_);
  or (_27480_, \oc8051_symbolic_cxrom1.regvalid [14], _27369_);
  and (_27481_, _27480_, _27479_);
  or (_27482_, _27481_, _27420_);
  or (_27483_, _27412_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_27484_, _27412_, _18644_);
  and (_27485_, _27484_, _27483_);
  or (_27486_, _27485_, _27416_);
  and (_27487_, _27486_, _27482_);
  or (_27488_, _27487_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_27489_, _27412_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_27490_, _27412_, _18657_);
  and (_27491_, _27490_, _27420_);
  and (_27492_, _27491_, _27489_);
  nand (_27493_, _27412_, _18532_);
  or (_27494_, \oc8051_symbolic_cxrom1.regvalid [12], _27369_);
  and (_27495_, _27494_, _27416_);
  and (_27496_, _27495_, _27493_);
  or (_27497_, _27496_, _27380_);
  or (_27498_, _27497_, _27492_);
  or (_27499_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27500_, _27499_, _27428_);
  or (_27501_, _27500_, _27376_);
  or (_27502_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27503_, \oc8051_symbolic_cxrom1.regvalid [11], _27369_);
  and (_27504_, _27503_, _27502_);
  or (_27505_, _27504_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27506_, _27505_, _27501_);
  and (_27507_, _27506_, _27414_);
  and (_27508_, _27380_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_27509_, _27375_, _27376_);
  or (_27510_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27511_, \oc8051_symbolic_cxrom1.regvalid [9], _27369_);
  and (_27512_, _27511_, _27510_);
  or (_27513_, _27512_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_27514_, _27513_, _27509_);
  and (_27515_, _27514_, _27508_);
  or (_27516_, _27515_, _27507_);
  and (_27517_, _27506_, _27380_);
  or (_27518_, _27517_, _27379_);
  and (_27519_, _27518_, _27516_);
  and (_27520_, _27519_, _27498_);
  and (_27521_, _27520_, _27488_);
  and (_27522_, _27521_, _27478_);
  or (_27523_, _27522_, _27459_);
  nor (_27524_, _26178_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_27525_, _26210_, _26185_);
  nor (_27526_, _27525_, _27524_);
  nor (_27527_, _27526_, _16190_);
  not (_27528_, _27527_);
  and (_27529_, _26156_, _16194_);
  and (_27530_, _26210_, _26164_);
  nor (_27531_, _27530_, _27529_);
  nor (_27532_, _27531_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_27533_, _21603_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_27534_, _18657_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_27535_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_27536_, _27535_, _27534_);
  and (_27537_, _27536_, _27533_);
  and (_27538_, _18635_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_27539_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_27540_, _27539_, _27538_);
  and (_27541_, _27540_, _21596_);
  nor (_27542_, _27541_, _27537_);
  not (_27543_, _27542_);
  nor (_27544_, _27543_, _27532_);
  and (_27545_, _27544_, _27528_);
  not (_27546_, _27545_);
  and (_27547_, _27546_, _26190_);
  nor (_27548_, _21608_, _16198_);
  and (_27549_, _27548_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_27550_, _27548_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_27551_, _27550_, _27549_);
  nand (_27552_, _27551_, _18622_);
  and (_27553_, _21608_, _16198_);
  nor (_27554_, _27553_, _27548_);
  not (_27555_, _27554_);
  nor (_27556_, _27555_, _21670_);
  and (_27557_, _27556_, _27552_);
  and (_27558_, _27551_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_27559_, _27551_, _18609_);
  or (_27560_, _27559_, _27558_);
  and (_27561_, _27560_, _27555_);
  or (_27562_, _27561_, _27557_);
  and (_27563_, _27562_, _21608_);
  nand (_27564_, _27551_, _18630_);
  nor (_27565_, _27555_, _21679_);
  and (_27566_, _27565_, _27564_);
  and (_27567_, _27551_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_27568_, _27551_, _18635_);
  or (_27569_, _27568_, _27567_);
  and (_27570_, _27569_, _27555_);
  or (_27571_, _27570_, _27566_);
  and (_27572_, _27571_, _21603_);
  or (_27573_, _27572_, _27563_);
  nand (_27574_, _27551_, _18646_);
  or (_27575_, _27551_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_27576_, _27575_, _27555_);
  and (_27577_, _27576_, _27574_);
  or (_27578_, _27551_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_27579_, _27555_, _26149_);
  and (_27580_, _27579_, _27578_);
  or (_27581_, _27580_, _27577_);
  and (_27582_, _27581_, _21595_);
  nand (_27583_, _27551_, _18663_);
  nor (_27584_, _27555_, _21675_);
  and (_27585_, _27584_, _27583_);
  and (_27586_, _27551_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_27587_, _27551_, _18657_);
  or (_27588_, _27587_, _27586_);
  and (_27589_, _27588_, _27555_);
  or (_27590_, _27589_, _27585_);
  and (_27591_, _27590_, _21605_);
  or (_27592_, _27591_, _27582_);
  or (_27593_, _27592_, _27573_);
  and (_27594_, _27593_, _21689_);
  and (_27595_, _27594_, _27547_);
  and (_27596_, _27595_, _27523_);
  and (_27597_, _15585_, _26138_);
  and (_27598_, _27597_, _27596_);
  and (_27599_, _27598_, _27367_);
  and (_27600_, _27599_, _27365_);
  and (property_invalid_jnc, _27600_, _27357_);
  and (_27601_, _27196_, _27210_);
  nor (_27602_, _27203_, _27210_);
  nor (_27603_, _27602_, _27601_);
  and (_27604_, _27603_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_27605_, _27603_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_27606_, _27088_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_27607_, _27088_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_27608_, _27607_, _27606_);
  and (_27609_, _27085_, _14132_);
  nor (_27610_, _27085_, _14132_);
  or (_27611_, _27610_, _27609_);
  or (_27612_, _27611_, _27608_);
  or (_27613_, _27612_, cy_reg);
  or (_27614_, _27214_, _14132_);
  nand (_27615_, _27214_, _14132_);
  and (_27616_, _27615_, _27614_);
  or (_27617_, _27222_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_27618_, _27222_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_27619_, _27618_, _27617_);
  or (_27620_, _27619_, _27210_);
  or (_27621_, _27620_, _27616_);
  and (_27622_, _27621_, _27613_);
  and (_27623_, _27095_, _27210_);
  nor (_27624_, _27237_, _27210_);
  nor (_27625_, _27624_, _27623_);
  and (_27626_, _27625_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_27627_, _27625_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_27628_, _27107_, _27210_);
  nor (_27629_, _27255_, _27210_);
  nor (_27630_, _27629_, _27628_);
  and (_27631_, _27630_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_27632_, _27630_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_27633_, _27117_, cy_reg);
  and (_27634_, _27272_, cy_reg);
  nor (_27635_, _27634_, _27633_);
  and (_27636_, _27635_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_27637_, _27635_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_27638_, _27123_, _27210_);
  and (_27639_, _27279_, cy_reg);
  nor (_27640_, _27639_, _27638_);
  and (_27641_, _27640_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_27642_, _27640_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_27643_, _27285_, cy_reg);
  and (_27644_, _27130_, _27210_);
  nor (_27645_, _27644_, _27643_);
  and (_27646_, _27645_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_27647_, _27645_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_27648_, _27136_, _27210_);
  and (_27649_, _27293_, cy_reg);
  nor (_27650_, _27649_, _27648_);
  and (_27651_, _27650_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_27652_, _27139_, cy_reg);
  and (_27653_, _27298_, cy_reg);
  nor (_27654_, _27653_, _27652_);
  and (_27655_, _27654_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_27656_, _27654_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27657_, _27305_, cy_reg);
  nor (_27658_, _27145_, cy_reg);
  nor (_27659_, _27658_, _27657_);
  and (_27660_, _27659_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_27661_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_27662_, _27320_, cy_reg);
  nor (_27663_, _27662_, _27661_);
  and (_27664_, _27663_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27665_, _27312_, _21940_);
  nor (_27666_, _27312_, _21940_);
  or (_27667_, _27666_, _27665_);
  or (_27668_, _27667_, _27210_);
  nand (_27669_, _27312_, _27210_);
  and (_27670_, _27669_, _27668_);
  nor (_27671_, _27663_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_27672_, _27671_, _27670_);
  or (_27673_, _27672_, _27664_);
  nor (_27674_, _27659_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_27675_, _27674_, _27673_);
  or (_27676_, _27675_, _27660_);
  or (_27677_, _27676_, _27656_);
  or (_27678_, _27677_, _27655_);
  nor (_27679_, _27650_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_27680_, _27679_, _27678_);
  or (_27681_, _27680_, _27651_);
  or (_27682_, _27681_, _27647_);
  or (_27683_, _27682_, _27646_);
  or (_27684_, _27683_, _27642_);
  or (_27685_, _27684_, _27641_);
  or (_27686_, _27685_, _27637_);
  or (_27687_, _27686_, _27636_);
  and (_27688_, _27110_, _27210_);
  and (_27689_, _27263_, cy_reg);
  nor (_27690_, _27689_, _27688_);
  nor (_27691_, _27690_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_27692_, _27690_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_27693_, _27692_, _27691_);
  or (_27694_, _27693_, _27687_);
  or (_27695_, _27694_, _27632_);
  or (_27696_, _27695_, _27631_);
  and (_27697_, _27101_, _27210_);
  and (_27698_, _27230_, cy_reg);
  nor (_27699_, _27698_, _27697_);
  and (_27700_, _27699_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_27701_, _27699_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_27702_, _27701_, _27700_);
  or (_27703_, _27702_, _27696_);
  or (_27704_, _27703_, _27627_);
  or (_27705_, _27704_, _27626_);
  or (_27706_, _27705_, _27622_);
  nor (_27707_, _27082_, cy_reg);
  nor (_27708_, _27349_, _27210_);
  nor (_27709_, _27708_, _27707_);
  and (_27710_, _27709_, _14137_);
  nor (_27711_, _27709_, _14137_);
  or (_27712_, _27711_, _27710_);
  or (_27713_, _27712_, _27706_);
  or (_27714_, _27713_, _27605_);
  or (_27715_, _27714_, _27604_);
  and (_27716_, _27362_, _26547_);
  and (_27717_, _27716_, _27599_);
  and (property_invalid_jc, _27717_, _27715_);
  or (_27718_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_27719_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_27720_, _27719_, _27718_);
  and (_27721_, _21940_, _27455_);
  nor (_27722_, _21940_, _27455_);
  or (_27723_, _27722_, _27721_);
  or (_27724_, _27723_, _27720_);
  or (_27725_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_27726_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27727_, _27726_, _27725_);
  and (_27728_, _21857_, _27376_);
  nor (_27729_, _21857_, _27376_);
  or (_27730_, _27729_, _27728_);
  or (_27731_, _27730_, _27727_);
  or (_27732_, _27731_, _27724_);
  or (_27733_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_27734_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_27735_, _27734_, _27733_);
  not (_27736_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_27737_, _21774_, _27736_);
  and (_27738_, _21774_, _27736_);
  or (_27739_, _27738_, _27737_);
  or (_27740_, _27739_, _27735_);
  not (_27741_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_27742_, _21983_, _27741_);
  nor (_27743_, _21983_, _27741_);
  or (_27744_, _27743_, _27742_);
  not (_27745_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_27746_, _21690_, _27745_);
  nor (_27747_, _21690_, _27745_);
  or (_27748_, _27747_, _27746_);
  or (_27749_, _27748_, _27744_);
  or (_27750_, _27749_, _27740_);
  or (_27751_, _27750_, _27732_);
  nor (_27752_, _27196_, _14142_);
  and (_27753_, _27196_, _14142_);
  or (_27754_, _27753_, _27752_);
  nor (_27755_, _27082_, _14137_);
  and (_27756_, _27082_, _14137_);
  or (_27757_, _27756_, _27755_);
  or (_27758_, _27757_, _27612_);
  or (_27759_, _27758_, _27754_);
  nor (_27760_, _26546_, _14110_);
  and (_27761_, _26546_, _14110_);
  or (_27762_, _27761_, _27760_);
  nor (_27763_, _26413_, _14116_);
  and (_27764_, _26413_, _14116_);
  or (_27765_, _27764_, _27763_);
  or (_27766_, _27765_, _27762_);
  and (_27767_, _26457_, _14121_);
  nor (_27768_, _26457_, _14121_);
  or (_27769_, _27768_, _27767_);
  or (_27770_, _27769_, _27248_);
  or (_27771_, _27770_, _27766_);
  or (_27772_, _27771_, _27759_);
  or (_27773_, _27772_, _27751_);
  nor (_27774_, _26323_, _26550_);
  and (_27775_, _27361_, _27774_);
  and (_27776_, _27775_, _27598_);
  and (property_invalid_ajmp, _27776_, _27773_);
  and (_27777_, _26210_, _26193_);
  and (_27778_, _26199_, _26165_);
  and (_27779_, _26203_, _26196_);
  or (_27780_, _27779_, _27778_);
  or (_27781_, _27780_, _27777_);
  and (_27782_, _26209_, _26158_);
  or (_27783_, _27782_, _27140_);
  or (_27784_, _27783_, _27781_);
  and (_27785_, _26216_, _26210_);
  or (_27786_, _27785_, _27139_);
  and (_27787_, _26225_, _26196_);
  and (_27788_, _26231_, _26158_);
  and (_27789_, _26221_, _26165_);
  or (_27790_, _27789_, _27788_);
  or (_27791_, _27790_, _27787_);
  or (_27792_, _27791_, _27786_);
  nand (_27793_, _27792_, _27784_);
  nor (_27794_, _27793_, _27545_);
  nand (_27795_, _27794_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_27796_, _27794_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_27797_, _27796_, _27795_);
  and (_27798_, _26461_, _26210_);
  and (_27799_, _26466_, _26165_);
  and (_27800_, _26470_, _26196_);
  or (_27801_, _27800_, _27799_);
  or (_27802_, _27801_, _27798_);
  and (_27803_, _26476_, _26158_);
  or (_27804_, _27803_, _27140_);
  or (_27805_, _27804_, _27802_);
  and (_27806_, _26482_, _26210_);
  or (_27807_, _27806_, _27139_);
  and (_27808_, _26491_, _26196_);
  and (_27809_, _26497_, _26158_);
  and (_27810_, _26487_, _26165_);
  or (_27811_, _27810_, _27809_);
  or (_27812_, _27811_, _27808_);
  or (_27813_, _27812_, _27807_);
  nand (_27814_, _27813_, _27805_);
  nor (_27815_, _27814_, _27545_);
  nand (_27816_, _27815_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_27817_, _27815_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_27818_, _27817_, _27816_);
  or (_27819_, _27818_, _27797_);
  and (_27820_, _26326_, _26210_);
  and (_27821_, _26331_, _26165_);
  and (_27822_, _26335_, _26196_);
  or (_27823_, _27822_, _27821_);
  or (_27824_, _27823_, _27820_);
  and (_27825_, _26341_, _26158_);
  or (_27826_, _27825_, _27140_);
  or (_27827_, _27826_, _27824_);
  and (_27828_, _26352_, _26165_);
  or (_27829_, _27828_, _27139_);
  and (_27830_, _26356_, _26196_);
  and (_27831_, _26362_, _26158_);
  and (_27832_, _26347_, _26210_);
  or (_27833_, _27832_, _27831_);
  or (_27834_, _27833_, _27830_);
  or (_27835_, _27834_, _27829_);
  nand (_27836_, _27835_, _27827_);
  nor (_27837_, _27836_, _27545_);
  nand (_27838_, _27837_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_27839_, _27837_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_27840_, _27839_, _27838_);
  and (_27841_, _26510_, _26165_);
  and (_27842_, _26505_, _26210_);
  and (_27843_, _26514_, _26196_);
  or (_27844_, _27843_, _27842_);
  or (_27845_, _27844_, _27841_);
  and (_27846_, _26520_, _26158_);
  or (_27847_, _27846_, _27140_);
  or (_27848_, _27847_, _27845_);
  and (_27849_, _26526_, _26210_);
  or (_27850_, _27849_, _27139_);
  and (_27851_, _26535_, _26196_);
  and (_27852_, _26541_, _26158_);
  and (_27853_, _26531_, _26165_);
  or (_27854_, _27853_, _27852_);
  or (_27855_, _27854_, _27851_);
  or (_27856_, _27855_, _27850_);
  nand (_27857_, _27856_, _27848_);
  nor (_27858_, _27857_, _27545_);
  nand (_27859_, _27858_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_27860_, _27858_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_27861_, _27860_, _27859_);
  or (_27862_, _27861_, _27840_);
  or (_27863_, _27862_, _27819_);
  and (_27864_, _26288_, _26165_);
  and (_27865_, _26283_, _26210_);
  and (_27866_, _26292_, _26196_);
  or (_27867_, _27866_, _27865_);
  or (_27868_, _27867_, _27864_);
  and (_27869_, _26298_, _26158_);
  or (_27870_, _27869_, _27140_);
  or (_27871_, _27870_, _27868_);
  and (_27872_, _26304_, _26210_);
  or (_27873_, _27872_, _27139_);
  and (_27874_, _26313_, _26196_);
  and (_27875_, _26319_, _26158_);
  and (_27876_, _26309_, _26165_);
  or (_27877_, _27876_, _27875_);
  or (_27878_, _27877_, _27874_);
  or (_27879_, _27878_, _27873_);
  nand (_27880_, _27879_, _27871_);
  nor (_27881_, _27880_, _27545_);
  nor (_27882_, _27881_, _27380_);
  and (_27883_, _27881_, _27380_);
  or (_27884_, _27883_, _27882_);
  and (_27885_, _26372_, _26210_);
  and (_27886_, _26377_, _26165_);
  and (_27887_, _26381_, _26196_);
  or (_27888_, _27887_, _27886_);
  or (_27889_, _27888_, _27885_);
  and (_27890_, _26387_, _26158_);
  or (_27891_, _27890_, _27140_);
  or (_27892_, _27891_, _27889_);
  and (_27893_, _26393_, _26210_);
  or (_27894_, _27893_, _27139_);
  and (_27895_, _26402_, _26196_);
  and (_27896_, _26408_, _26158_);
  and (_27897_, _26398_, _26165_);
  or (_27898_, _27897_, _27896_);
  or (_27899_, _27898_, _27895_);
  or (_27900_, _27899_, _27894_);
  nand (_27901_, _27900_, _27892_);
  nor (_27902_, _27901_, _27545_);
  and (_27903_, _27902_, _27745_);
  nor (_27904_, _27902_, _27745_);
  or (_27905_, _27904_, _27903_);
  or (_27906_, _27905_, _27884_);
  and (_27907_, _26260_, _26210_);
  and (_27908_, _26269_, _26196_);
  nor (_27909_, _27908_, _27907_);
  and (_27910_, _26275_, _26158_);
  and (_27911_, _26265_, _26165_);
  nor (_27912_, _27911_, _27910_);
  and (_27913_, _27912_, _27909_);
  nor (_27914_, _27913_, _27139_);
  and (_27915_, _26239_, _26210_);
  and (_27916_, _26248_, _26196_);
  nor (_27917_, _27916_, _27915_);
  and (_27918_, _26254_, _26158_);
  and (_27919_, _26244_, _26165_);
  nor (_27920_, _27919_, _27918_);
  and (_27921_, _27920_, _27917_);
  nor (_27922_, _27921_, _27140_);
  nor (_27923_, _27922_, _27914_);
  nor (_27924_, _27923_, _27545_);
  nor (_27925_, _27924_, _27376_);
  and (_27926_, _27924_, _27376_);
  or (_27927_, _27926_, _27925_);
  and (_27928_, _26416_, _26210_);
  and (_27929_, _26421_, _26165_);
  and (_27930_, _26425_, _26196_);
  or (_27931_, _27930_, _27929_);
  or (_27932_, _27931_, _27928_);
  and (_27933_, _26431_, _26158_);
  or (_27934_, _27933_, _27140_);
  or (_27935_, _27934_, _27932_);
  and (_27936_, _26437_, _26210_);
  or (_27937_, _27936_, _27139_);
  and (_27938_, _26446_, _26196_);
  and (_27939_, _26452_, _26158_);
  and (_27940_, _26442_, _26165_);
  or (_27941_, _27940_, _27939_);
  or (_27942_, _27941_, _27938_);
  or (_27943_, _27942_, _27937_);
  nand (_27944_, _27943_, _27935_);
  nor (_27945_, _27944_, _27545_);
  nor (_27946_, _27945_, _27741_);
  and (_27947_, _27945_, _27741_);
  or (_27948_, _27947_, _27946_);
  or (_27949_, _27948_, _27927_);
  or (_27950_, _27949_, _27906_);
  or (_27951_, _27950_, _27863_);
  or (_27952_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_27953_, _21898_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_27954_, _27953_, _27952_);
  nor (_27955_, _21940_, _14110_);
  and (_27956_, _21940_, _14110_);
  or (_27957_, _27956_, _27955_);
  or (_27958_, _27957_, _27954_);
  or (_27959_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_27960_, _21816_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_27961_, _27960_, _27959_);
  and (_27962_, _21857_, _14121_);
  nor (_27963_, _21857_, _14121_);
  or (_27964_, _27963_, _27962_);
  or (_27965_, _27964_, _27961_);
  or (_27966_, _27965_, _27958_);
  or (_27967_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_27968_, _21732_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_27969_, _27968_, _27967_);
  and (_27970_, _21774_, _14127_);
  nor (_27971_, _21774_, _14127_);
  or (_27972_, _27971_, _27970_);
  or (_27973_, _27972_, _27969_);
  and (_27974_, _21983_, _14142_);
  nor (_27975_, _21983_, _14142_);
  or (_27976_, _27975_, _27974_);
  nor (_27977_, _21690_, _14137_);
  and (_27978_, _21690_, _14137_);
  or (_27979_, _27978_, _27977_);
  or (_27980_, _27979_, _27976_);
  or (_27981_, _27980_, _27973_);
  or (_27982_, _27981_, _27966_);
  or (_27983_, _27982_, _27951_);
  not (_27984_, _26546_);
  and (_27985_, _27984_, _26458_);
  and (_27986_, _27361_, _26550_);
  and (_27987_, _27986_, _27358_);
  and (_27988_, _27987_, _27985_);
  and (_27989_, _27988_, _27598_);
  and (property_invalid_ljmp, _27989_, _27983_);
  and (_27990_, _27203_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_27991_, _27203_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_27992_, _27255_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_27993_, _27255_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_27994_, _27263_, _14110_);
  nor (_27995_, _27263_, _14110_);
  and (_27996_, _27272_, _27741_);
  nor (_27997_, _27272_, _27741_);
  and (_27998_, _27279_, _27745_);
  nor (_27999_, _27279_, _27745_);
  not (_28000_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_28001_, _27285_, _28000_);
  nor (_28002_, _27285_, _28000_);
  and (_28003_, _27293_, _27736_);
  and (_28004_, _27298_, _27369_);
  nor (_28005_, _27298_, _27369_);
  and (_28006_, _27305_, _27376_);
  or (_28007_, _27320_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_28008_, _27320_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_28009_, _28008_, _28007_);
  or (_28010_, _28009_, _27667_);
  nor (_28011_, _27305_, _27376_);
  or (_28012_, _28011_, _28010_);
  or (_28013_, _28012_, _28006_);
  or (_28014_, _28013_, _28005_);
  or (_28015_, _28014_, _28004_);
  nor (_28016_, _27293_, _27736_);
  or (_28017_, _28016_, _28015_);
  or (_28018_, _28017_, _28003_);
  or (_28019_, _28018_, _28002_);
  or (_28020_, _28019_, _28001_);
  or (_28021_, _28020_, _27999_);
  or (_28022_, _28021_, _27998_);
  or (_28023_, _28022_, _27997_);
  or (_28024_, _28023_, _27996_);
  or (_28025_, _28024_, _27995_);
  or (_28026_, _28025_, _27994_);
  or (_28027_, _28026_, _27993_);
  or (_28028_, _28027_, _27992_);
  or (_28029_, _28028_, _27241_);
  or (_28030_, _28029_, _27619_);
  or (_28031_, _28030_, _27616_);
  nor (_28032_, _27349_, _14137_);
  and (_28033_, _27349_, _14137_);
  or (_28034_, _28033_, _28032_);
  or (_28035_, _28034_, _28031_);
  or (_28036_, _28035_, _27991_);
  or (_28037_, _28036_, _27990_);
  not (_28038_, _26413_);
  and (_28039_, _26457_, _28038_);
  and (_28040_, _28039_, _26547_);
  and (_28041_, _28040_, _27362_);
  and (_28042_, _28041_, _27598_);
  and (property_invalid_sjmp, _28042_, _28037_);
  and (_28043_, _27549_, _27072_);
  and (_28044_, _28043_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_28045_, _28044_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_28046_, _28045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_28047_, _28046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_28048_, _28047_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_28049_, _28048_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_28050_, _28049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_28051_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_28052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_28053_, _28052_, _28051_);
  nor (_28054_, _28049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_28055_, _28054_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_28056_, _28055_, _28053_);
  nor (_28057_, _28056_, _28050_);
  or (_28058_, _28054_, _28050_);
  and (_28059_, _28058_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_28060_, _28043_, _27075_);
  nor (_28061_, _28045_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_28062_, _28061_, _28060_);
  and (_28063_, _28062_, _14121_);
  and (_28064_, _27549_, _27071_);
  nor (_28065_, _28064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_28066_, _28065_, _28043_);
  and (_28067_, _28066_, _27741_);
  nor (_28068_, _28066_, _27741_);
  or (_28069_, _28068_, _28067_);
  or (_28070_, _28069_, _28063_);
  and (_28071_, _27549_, _27070_);
  and (_28072_, _27549_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_28073_, _28072_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_28074_, _28073_, _28071_);
  nor (_28075_, _28074_, _28000_);
  or (_28076_, _27551_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_28077_, _27551_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_28078_, _28077_, _28076_);
  and (_28079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_28080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_28081_, _28080_, _28079_);
  nand (_28082_, _28081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_28083_, _28081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_28084_, _28083_, _28082_);
  nand (_28085_, _28084_, _27313_);
  or (_28086_, _27554_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_28087_, _27554_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_28088_, _28087_, _28086_);
  or (_28089_, _28088_, _28085_);
  or (_28090_, _28089_, _28078_);
  or (_28091_, _28090_, _28075_);
  nor (_28092_, _28043_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_28093_, _28092_, _28044_);
  nor (_28094_, _28093_, _14110_);
  and (_28095_, _28093_, _14110_);
  or (_28096_, _28095_, _28094_);
  or (_28097_, _28096_, _28091_);
  nor (_28098_, _28071_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_28099_, _28098_, _28064_);
  nor (_28100_, _28099_, _27745_);
  and (_28101_, _28099_, _27745_);
  or (_28102_, _28101_, _28100_);
  or (_28103_, _28102_, _28097_);
  nor (_28104_, _28062_, _14121_);
  nor (_28105_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_28106_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_28107_, _28106_, _28105_);
  or (_28108_, _28107_, _28044_);
  nand (_28109_, _28107_, _28044_);
  and (_28110_, _28109_, _28108_);
  nor (_28111_, _27549_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_28112_, _28111_, _28072_);
  nand (_28113_, _28112_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_28114_, _28112_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_28115_, _28114_, _28113_);
  and (_28116_, _28074_, _28000_);
  or (_28117_, _28116_, _28115_);
  or (_28118_, _28117_, _28110_);
  or (_28119_, _28118_, _28104_);
  or (_28120_, _28119_, _28103_);
  or (_28121_, _28120_, _28070_);
  and (_28122_, _28060_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_28123_, _28122_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_28124_, _28123_, _28048_);
  and (_28125_, _28124_, _14127_);
  nor (_28126_, _28124_, _14127_);
  or (_28127_, _28126_, _28125_);
  or (_28128_, _28127_, _28121_);
  not (_28129_, _28053_);
  and (_28130_, _28129_, _28050_);
  nor (_28131_, _28046_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_28132_, _28131_, _28047_);
  nor (_28133_, _28132_, _14106_);
  and (_28134_, _28132_, _14106_);
  or (_28135_, _28134_, _28133_);
  nor (_28136_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_28137_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_28138_, _28137_, _28136_);
  not (_28139_, _28138_);
  and (_28140_, _28139_, _28048_);
  nor (_28141_, _28139_, _28048_);
  or (_28142_, _28141_, _28140_);
  or (_28143_, _28142_, _28135_);
  or (_28144_, _28143_, _28130_);
  or (_28145_, _28144_, _28128_);
  or (_28146_, _28145_, _28059_);
  or (_28147_, _28146_, _28057_);
  not (_28148_, _26502_);
  and (_28149_, _28148_, _26369_);
  and (_28150_, _28149_, _27984_);
  or (_28151_, _28150_, _27365_);
  and (_28152_, _28151_, _28039_);
  and (_28153_, _26545_, _26413_);
  and (_28154_, _28153_, _26369_);
  and (_28155_, _26502_, _27366_);
  and (_28156_, _28155_, _28154_);
  and (_28157_, _26545_, _26502_);
  and (_28158_, _27358_, _26236_);
  and (_28159_, _28158_, _27361_);
  nand (_28160_, _28159_, _27367_);
  nor (_28161_, _28160_, _28157_);
  or (_28162_, _28161_, _28156_);
  or (_28163_, _28162_, _28152_);
  and (_28164_, _28163_, _27598_);
  and (property_invalid_pcp3, _28164_, _28147_);
  and (_28165_, _28148_, _27360_);
  and (_28166_, _27364_, _26368_);
  or (_28167_, _28166_, _28165_);
  and (_28168_, _28167_, _28038_);
  or (_28169_, _26413_, _27358_);
  and (_28170_, _28169_, _27984_);
  and (_28171_, _28170_, _27986_);
  or (_28172_, _28154_, _27366_);
  or (_28173_, _28172_, _28171_);
  or (_28174_, _28173_, _28168_);
  and (_28175_, _27984_, _26369_);
  and (_28176_, _28153_, _27360_);
  and (_28177_, _28176_, _26502_);
  or (_28178_, _28177_, _26457_);
  or (_28179_, _28178_, _28175_);
  and (_28180_, _28179_, _28174_);
  or (_28181_, _27987_, _26551_);
  and (_28182_, _28181_, _27366_);
  or (_28183_, _28182_, _28149_);
  and (_28184_, _28183_, _26413_);
  and (_28185_, _27358_, _26280_);
  and (_28186_, _28185_, _28148_);
  and (_28187_, _27986_, _26545_);
  or (_28188_, _28187_, _28186_);
  and (_28189_, _28188_, _28039_);
  and (_28190_, _28157_, _27367_);
  and (_28191_, _28190_, _28185_);
  and (_28192_, _26546_, _26368_);
  and (_28193_, _28192_, _26458_);
  or (_28194_, _28193_, _28191_);
  or (_28195_, _28194_, _28189_);
  or (_28196_, _28195_, _28184_);
  or (_28197_, _28196_, _28180_);
  nor (_28198_, _27123_, _27745_);
  nor (_28199_, _27110_, _14110_);
  or (_28200_, _28199_, _28198_);
  and (_28201_, _27123_, _27745_);
  and (_28202_, _27110_, _14110_);
  or (_28203_, _28202_, _28201_);
  or (_28204_, _28203_, _28200_);
  and (_28205_, _27117_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_28206_, _27130_, _28000_);
  or (_28207_, _28206_, _28205_);
  and (_28208_, _27130_, _28000_);
  not (_28209_, _27098_);
  nor (_28210_, _28107_, _28209_);
  or (_28211_, _28210_, _28208_);
  or (_28212_, _28211_, _28207_);
  and (_28213_, _27139_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_28214_, _27139_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_28215_, _28214_, _28213_);
  and (_28216_, _27145_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_28217_, _28081_, _27312_);
  nor (_28218_, _27145_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_28219_, _28218_, _28217_);
  or (_28220_, _28219_, _28216_);
  or (_28221_, _28220_, _28215_);
  nor (_28222_, _27136_, _27736_);
  and (_28223_, _27136_, _27736_);
  or (_28224_, _28223_, _28222_);
  or (_28225_, _28224_, _28221_);
  and (_28226_, _28107_, _28209_);
  nor (_28227_, _27117_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_28228_, _28227_, _28226_);
  or (_28229_, _28228_, _28225_);
  or (_28230_, _28229_, _28212_);
  or (_28231_, _28230_, _28204_);
  or (_28232_, _28231_, _27248_);
  or (_28233_, _28232_, _27245_);
  or (_28234_, _28233_, _27759_);
  and (_28235_, _28234_, _27598_);
  and (property_invalid_pcp2, _28235_, _28197_);
  not (_28236_, _26235_);
  and (_28237_, _26280_, _28236_);
  or (_28238_, _28237_, _28158_);
  nor (_28239_, _27366_, _26366_);
  and (_28240_, _28239_, _28238_);
  and (_28241_, _26545_, _28236_);
  and (_28242_, _28241_, _26457_);
  or (_28243_, _28165_, _28038_);
  or (_28244_, _28243_, _28242_);
  or (_28245_, _28244_, _28186_);
  or (_28246_, _28245_, _28240_);
  and (_28247_, _26551_, _26547_);
  and (_28248_, _27363_, _27360_);
  and (_28249_, _28248_, _26502_);
  or (_28250_, _28159_, _26413_);
  or (_28251_, _28250_, _28249_);
  or (_28252_, _28251_, _28247_);
  and (_28253_, _28252_, _28246_);
  and (_28254_, _28176_, _26457_);
  and (_28255_, _27359_, _26548_);
  nor (_28256_, _27363_, _26502_);
  and (_28257_, _28256_, _26368_);
  and (_28258_, _28257_, _28039_);
  or (_28259_, _28258_, _28255_);
  or (_28260_, _28259_, _28254_);
  or (_28261_, _28185_, _27360_);
  nand (_28262_, _27984_, _26501_);
  nor (_28263_, _28262_, _27360_);
  or (_28264_, _28263_, _26458_);
  and (_28265_, _28264_, _28261_);
  and (_28266_, _28248_, _27366_);
  and (_28267_, _28237_, _27985_);
  or (_28268_, _28267_, _28266_);
  or (_28269_, _28268_, _28265_);
  or (_28270_, _28269_, _28260_);
  or (_28271_, _28270_, _28253_);
  nor (_28272_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_28273_, _27072_, _21597_);
  and (_28274_, _28273_, _27075_);
  or (_28275_, _28274_, _28272_);
  nor (_28276_, _28275_, _27100_);
  nor (_28277_, _28276_, _14121_);
  and (_28278_, _28273_, _27076_);
  and (_28279_, _28278_, _16238_);
  nor (_28280_, _28278_, _16238_);
  or (_28281_, _28280_, _28279_);
  nand (_28282_, _28281_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_28283_, _28281_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_28284_, _28283_, _28282_);
  or (_28285_, _28284_, _28277_);
  and (_28286_, _27078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_28287_, _28286_, _28138_);
  or (_28288_, _28286_, _28138_);
  and (_28289_, _28288_, _28287_);
  and (_28290_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], _16190_);
  and (_28291_, _27130_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_28292_, _28291_, _28290_);
  or (_28293_, _28292_, _28000_);
  nand (_28294_, _28292_, _28000_);
  and (_28295_, _28294_, _28293_);
  or (_28296_, _28295_, _28289_);
  or (_28297_, _28296_, _28285_);
  and (_28298_, _27114_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_28299_, _27070_, _21597_);
  nor (_28300_, _28299_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_28301_, _28300_, _28298_);
  and (_28302_, _28301_, _27745_);
  nor (_28303_, _28301_, _27745_);
  and (_28304_, _21602_, _27376_);
  nor (_28305_, _21602_, _27376_);
  or (_28306_, _28305_, _28084_);
  or (_28307_, _28306_, _28304_);
  or (_28308_, _28307_, _28303_);
  or (_28309_, _28308_, _28302_);
  nor (_28310_, _28298_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_28311_, _28310_, _28273_);
  nor (_28312_, _28311_, _27741_);
  and (_28313_, _21599_, _27369_);
  nor (_28314_, _21599_, _27369_);
  nor (_28315_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_28316_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_28317_, _28316_, _28315_);
  not (_28318_, _28317_);
  nor (_28319_, _28318_, _21597_);
  and (_28320_, _28318_, _21597_);
  or (_28321_, _28320_, _27312_);
  or (_28322_, _28321_, _28319_);
  or (_28323_, _28322_, _28314_);
  or (_28324_, _28323_, _28313_);
  or (_28325_, _28324_, _28312_);
  nor (_28326_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_28327_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28328_, _28327_, _28326_);
  or (_28329_, _28328_, _28274_);
  nand (_28330_, _28328_, _28274_);
  and (_28331_, _28330_, _28329_);
  and (_28332_, _28311_, _27741_);
  or (_28333_, _28332_, _28331_);
  or (_28334_, _28333_, _28325_);
  or (_28335_, _28334_, _28309_);
  and (_28336_, _28276_, _14121_);
  nand (_28337_, _28273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_28338_, _28337_, _28107_);
  and (_28339_, _28210_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_28340_, _28339_, _28338_);
  or (_28341_, _28273_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_28342_, _28341_, _28337_);
  and (_28343_, _28342_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_28344_, _28342_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_28345_, _28344_, _28343_);
  or (_28346_, _28345_, _28340_);
  or (_28347_, _28346_, _28336_);
  or (_28348_, _28347_, _28335_);
  or (_28349_, _28348_, _28297_);
  and (_28350_, _27080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_28351_, _28350_, _28053_);
  nand (_28352_, _28350_, _28053_);
  and (_28353_, _28352_, _28351_);
  nand (_28354_, _27079_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_28355_, _28354_, _16246_);
  nor (_28356_, _28355_, _28350_);
  and (_28357_, _28356_, _14137_);
  nor (_28358_, _28356_, _14137_);
  or (_28359_, _28358_, _28357_);
  or (_28360_, _28359_, _28353_);
  or (_28361_, _28360_, _28349_);
  and (_28362_, _28361_, _27598_);
  and (property_invalid_pcp1, _28362_, _28271_);
  and (_28363_, _26138_, pc_change_r);
  and (_28364_, _28363_, _27596_);
  and (_28365_, acc_reg[0], acc_reg[1]);
  and (_28366_, _28365_, acc_reg[2]);
  and (_28367_, _28366_, acc_reg[3]);
  and (_28368_, _28367_, acc_reg[4]);
  and (_28369_, _28368_, acc_reg[5]);
  and (_28370_, _28369_, acc_reg[6]);
  nor (_28371_, acc_reg[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_28372_, acc_reg[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_28373_, _28372_, _28371_);
  nor (_28374_, _28369_, acc_reg[6]);
  nor (_28375_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_28376_, _28375_, _28373_);
  nor (_28377_, _28376_, _28370_);
  not (_28378_, _28373_);
  and (_28379_, _28378_, _28370_);
  nor (_28380_, _28368_, acc_reg[5]);
  nor (_28381_, _28380_, _28369_);
  nor (_28382_, _28381_, _33948_);
  and (_28383_, _28381_, _33948_);
  or (_28384_, _28383_, _28382_);
  or (_28385_, _28384_, _28379_);
  or (_28386_, _28374_, _28370_);
  and (_28387_, _28386_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_28388_, _28366_, acc_reg[3]);
  nor (_28389_, _28388_, _28367_);
  and (_28390_, _28389_, _34032_);
  nor (_28391_, _28389_, _34032_);
  or (_28392_, _28391_, _28390_);
  and (_28393_, acc_reg[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_28394_, acc_reg[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_28395_, _28394_, _28393_);
  not (_28396_, acc_reg[0]);
  and (_28397_, _28396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand (_28398_, _28397_, _28395_);
  or (_28399_, _28396_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_28400_, _28399_, _28395_);
  and (_28401_, _28400_, _28398_);
  nor (_28402_, _28365_, acc_reg[2]);
  nor (_28403_, _28402_, _28366_);
  nor (_28404_, _28403_, _34059_);
  and (_28405_, _28403_, _34059_);
  or (_28406_, _28405_, _28404_);
  or (_28407_, _28406_, _28401_);
  or (_28408_, _28407_, _28392_);
  nor (_28409_, _28367_, acc_reg[4]);
  nor (_28410_, _28409_, _28368_);
  nor (_28411_, _28410_, _33984_);
  and (_28412_, _28410_, _33984_);
  or (_28413_, _28412_, _28411_);
  or (_28414_, _28413_, _28408_);
  or (_28415_, _28414_, _28387_);
  or (_28416_, _28415_, _28385_);
  or (_28417_, _28416_, _28377_);
  and (_28418_, _28417_, pc_inc_acc_r);
  and (property_invalid_inc_acc, _28418_, _28364_);
  not (_28419_, op1_out_r[0]);
  and (_28420_, _28419_, op1_out_r[1]);
  and (_28421_, op1_out_r[2], op1_out_r[3]);
  and (_28422_, _28421_, _28420_);
  not (_28423_, op1_out_r[5]);
  and (_28424_, op1_out_r[4], _28423_);
  and (_28425_, op1_out_r[7], op1_out_r[6]);
  and (_28426_, _28425_, _28424_);
  and (_28427_, _28426_, _28422_);
  nor (_28428_, _28419_, op1_out_r[1]);
  not (_28429_, op1_out_r[3]);
  and (_28430_, op1_out_r[2], _28429_);
  and (_28431_, _28430_, _28428_);
  and (_28432_, _28431_, _28426_);
  nor (_28433_, _28432_, _28427_);
  and (_28434_, _28428_, _28421_);
  and (_28435_, _28434_, _28426_);
  nor (_28436_, op1_out_r[2], op1_out_r[3]);
  and (_28437_, _28436_, _28428_);
  nor (_28438_, op1_out_r[4], op1_out_r[5]);
  not (_28439_, op1_out_r[7]);
  and (_28440_, _28439_, op1_out_r[6]);
  and (_28441_, _28440_, _28438_);
  and (_28442_, _28441_, _28437_);
  nor (_28443_, _28442_, _28435_);
  and (_28444_, _28443_, _28433_);
  and (_28445_, op1_out_r[0], op1_out_r[1]);
  and (_28446_, _28445_, _28421_);
  and (_28447_, _28438_, _28425_);
  and (_28448_, _28447_, _28446_);
  and (_28449_, _28436_, _28420_);
  and (_28450_, _28449_, _28426_);
  nor (_28451_, _28450_, _28448_);
  and (_28452_, _28440_, _28424_);
  and (_28453_, _28452_, _28446_);
  nor (_28454_, op1_out_r[4], _28423_);
  and (_28455_, _28454_, _28440_);
  and (_28456_, _28455_, _28449_);
  nor (_28457_, _28456_, _28453_);
  and (_28458_, _28457_, _28451_);
  and (_28459_, _28458_, _28444_);
  nor (_28460_, _28439_, op1_out_r[6]);
  and (_28461_, _28460_, _28454_);
  and (_28462_, _28461_, _28431_);
  and (_28463_, _28430_, _28420_);
  and (_28464_, _28463_, _28461_);
  nor (_28465_, _28464_, _28462_);
  and (_28466_, op1_out_r[4], op1_out_r[5]);
  and (_28467_, _28466_, _28460_);
  and (_28468_, _28467_, _28434_);
  nor (_28469_, op1_out_r[2], _28429_);
  and (_28470_, _28469_, _28445_);
  and (_28471_, _28470_, _28467_);
  nor (_28472_, _28471_, _28468_);
  and (_28473_, _28472_, _28465_);
  and (_28474_, _28467_, _28463_);
  nor (_28475_, op1_out_r[0], op1_out_r[1]);
  and (_28476_, _28475_, _28469_);
  and (_28477_, _28476_, _28467_);
  nor (_28478_, _28477_, _28474_);
  and (_28479_, _28445_, _28436_);
  and (_28480_, _28479_, _28426_);
  and (_28481_, _28463_, _28426_);
  nor (_28482_, _28481_, _28480_);
  and (_28483_, _28482_, _28478_);
  and (_28484_, _28483_, _28473_);
  and (_28485_, _28484_, _28459_);
  and (_28486_, _28467_, _28437_);
  and (_28487_, _28445_, _28430_);
  and (_28488_, _28487_, _28467_);
  nor (_28489_, _28488_, _28486_);
  and (_28490_, _28475_, _28436_);
  and (_28491_, _28490_, _28467_);
  and (_28492_, _28469_, _28420_);
  and (_28493_, _28492_, _28467_);
  nor (_28494_, _28493_, _28491_);
  and (_28495_, _28494_, _28489_);
  and (_28496_, _28467_, _28449_);
  and (_28497_, _28461_, _28446_);
  nor (_28498_, _28497_, _28496_);
  and (_28499_, _28454_, _28425_);
  and (_28500_, _28499_, _28479_);
  and (_28501_, _28446_, _28426_);
  nor (_28502_, _28501_, _28500_);
  and (_28503_, _28502_, _28498_);
  and (_28504_, _28503_, _28495_);
  and (_28505_, _28466_, _28440_);
  and (_28506_, _28505_, _28463_);
  and (_28507_, _28505_, _28431_);
  nor (_28508_, _28507_, _28506_);
  and (_28509_, _28475_, _28430_);
  and (_28510_, _28509_, _28467_);
  and (_28511_, _28509_, _28505_);
  nor (_28512_, _28511_, _28510_);
  and (_28513_, _28512_, _28508_);
  and (_28514_, _28475_, _28421_);
  and (_28515_, _28514_, _28426_);
  and (_28516_, _28470_, _28426_);
  nor (_28517_, _28516_, _28515_);
  and (_28518_, _28467_, _28431_);
  and (_28519_, _28467_, _28422_);
  nor (_28520_, _28519_, _28518_);
  and (_28521_, _28520_, _28517_);
  and (_28522_, _28521_, _28513_);
  and (_28523_, _28522_, _28504_);
  and (_28524_, _28523_, _28485_);
  and (_28525_, _28460_, _28438_);
  and (_28526_, _28525_, _28437_);
  nor (_28527_, op1_out_r[7], op1_out_r[6]);
  and (_28528_, _28527_, _28454_);
  and (_28529_, _28528_, _28431_);
  nor (_28530_, _28529_, _28526_);
  and (_28531_, _28525_, _28470_);
  and (_28532_, _28525_, _28490_);
  nor (_28533_, _28532_, _28531_);
  and (_28534_, _28533_, _28530_);
  and (_28535_, _28455_, _28431_);
  and (_28536_, _28509_, _28455_);
  nor (_28537_, _28536_, _28535_);
  and (_28538_, _28527_, _28438_);
  and (_28539_, _28538_, _28431_);
  and (_28540_, _28538_, _28509_);
  nor (_28541_, _28540_, _28539_);
  and (_28542_, _28541_, _28537_);
  and (_28543_, _28542_, _28534_);
  and (_28544_, _28466_, _28425_);
  and (_28545_, _28544_, _28509_);
  and (_28546_, _28544_, _28479_);
  nor (_28547_, _28546_, _28545_);
  and (_28548_, _28525_, _28422_);
  and (_28549_, _28460_, _28424_);
  and (_28550_, _28549_, _28490_);
  nor (_28551_, _28550_, _28548_);
  and (_28552_, _28551_, _28547_);
  and (_28553_, _28525_, _28514_);
  and (_28554_, _28469_, _28428_);
  and (_28555_, _28554_, _28528_);
  nor (_28556_, _28555_, _28553_);
  and (_28557_, _28549_, _28437_);
  and (_28558_, _28525_, _28449_);
  nor (_28559_, _28558_, _28557_);
  and (_28560_, _28559_, _28556_);
  and (_28561_, _28560_, _28552_);
  and (_28562_, _28561_, _28543_);
  and (_28563_, _28499_, _28434_);
  and (_28564_, _28499_, _28422_);
  nor (_28565_, _28564_, _28563_);
  and (_28566_, _28514_, _28499_);
  and (_28567_, _28525_, _28463_);
  nor (_28568_, _28567_, _28566_);
  and (_28569_, _28568_, _28565_);
  and (_28570_, _28479_, _28461_);
  and (_28571_, _28525_, _28509_);
  nor (_28572_, _28571_, _28570_);
  and (_28573_, _28554_, _28549_);
  and (_28574_, _28505_, _28446_);
  nor (_28575_, _28574_, _28573_);
  and (_28576_, _28575_, _28572_);
  and (_28577_, _28576_, _28569_);
  and (_28578_, _28490_, _28461_);
  and (_28579_, _28527_, _28424_);
  and (_28580_, _28579_, _28446_);
  nor (_28581_, _28580_, _28578_);
  and (_28582_, _28538_, _28463_);
  and (_28583_, _28479_, _28455_);
  nor (_28584_, _28583_, _28582_);
  and (_28585_, _28584_, _28581_);
  and (_28586_, _28525_, _28479_);
  and (_28587_, _28525_, _28431_);
  nor (_28588_, _28587_, _28586_);
  and (_28589_, _28461_, _28437_);
  and (_28590_, _28487_, _28461_);
  nor (_28591_, _28590_, _28589_);
  and (_28592_, _28591_, _28588_);
  and (_28593_, _28592_, _28585_);
  and (_28594_, _28593_, _28577_);
  and (_28595_, _28594_, _28562_);
  and (_28596_, _28595_, _28524_);
  and (_28597_, _28528_, _28487_);
  and (_28598_, _28527_, _28466_);
  and (_28599_, _28598_, _28554_);
  nor (_28600_, _28599_, _28597_);
  and (_28601_, _28505_, _28476_);
  and (_28602_, _28505_, _28422_);
  nor (_28603_, _28602_, _28601_);
  and (_28604_, _28603_, _28600_);
  and (_28605_, _28598_, _28476_);
  and (_28606_, _28598_, _28422_);
  nor (_28607_, _28606_, _28605_);
  and (_28608_, _28528_, _28492_);
  and (_28609_, _28528_, _28476_);
  nor (_28610_, _28609_, _28608_);
  and (_28611_, _28610_, _28607_);
  and (_28612_, _28611_, _28604_);
  and (_28613_, _28554_, _28467_);
  and (_28614_, _28455_, _28422_);
  nor (_28615_, _28614_, _28613_);
  and (_28616_, _28499_, _28431_);
  and (_28617_, _28455_, _28434_);
  nor (_28618_, _28617_, _28616_);
  and (_28619_, _28618_, _28615_);
  and (_28620_, _28505_, _28492_);
  and (_28621_, _28598_, _28492_);
  nor (_28622_, _28621_, _28620_);
  and (_28623_, _28505_, _28487_);
  and (_28624_, _28598_, _28487_);
  nor (_28625_, _28624_, _28623_);
  and (_28626_, _28625_, _28622_);
  and (_28627_, _28626_, _28619_);
  and (_28628_, _28627_, _28612_);
  and (_28629_, _28549_, _28422_);
  and (_28630_, _28549_, _28434_);
  nor (_28631_, _28630_, _28629_);
  and (_28632_, _28549_, _28470_);
  and (_28633_, _28549_, _28514_);
  nor (_28634_, _28633_, _28632_);
  and (_28635_, _28634_, _28631_);
  and (_28636_, _28461_, _28422_);
  and (_28637_, _28461_, _28434_);
  nor (_28638_, _28637_, _28636_);
  and (_28639_, _28470_, _28461_);
  and (_28640_, _28514_, _28461_);
  nor (_28641_, _28640_, _28639_);
  and (_28642_, _28641_, _28638_);
  and (_28643_, _28642_, _28635_);
  and (_28644_, _28544_, _28487_);
  and (_28645_, _28544_, _28476_);
  nor (_28646_, _28645_, _28644_);
  and (_28647_, _28452_, _28431_);
  and (_28648_, _28479_, _28452_);
  nor (_28649_, _28648_, _28647_);
  and (_28650_, _28649_, _28646_);
  and (_28651_, _28549_, _28487_);
  and (_28652_, _28549_, _28476_);
  nor (_28653_, _28652_, _28651_);
  and (_28654_, _28487_, _28441_);
  and (_28655_, _28549_, _28492_);
  nor (_28656_, _28655_, _28654_);
  and (_28657_, _28656_, _28653_);
  and (_28658_, _28657_, _28650_);
  and (_28659_, _28658_, _28643_);
  and (_28660_, _28659_, _28628_);
  and (_28661_, _28452_, _28449_);
  and (_28662_, _28505_, _28449_);
  nor (_28663_, _28662_, _28661_);
  and (_28664_, _28441_, _28422_);
  and (_28665_, _28455_, _28446_);
  nor (_28666_, _28665_, _28664_);
  and (_28667_, _28666_, _28663_);
  and (_28668_, _28452_, _28437_);
  and (_28669_, _28505_, _28479_);
  nor (_28670_, _28669_, _28668_);
  and (_28671_, _28509_, _28452_);
  and (_28672_, _28490_, _28452_);
  nor (_28673_, _28672_, _28671_);
  and (_28674_, _28673_, _28670_);
  and (_28675_, _28674_, _28667_);
  and (_28676_, _28598_, _28437_);
  and (_28677_, _28554_, _28447_);
  nor (_28678_, _28677_, _28676_);
  and (_28679_, _28554_, _28499_);
  and (_28680_, _28447_, _28434_);
  nor (_28681_, _28680_, _28679_);
  and (_28682_, _28681_, _28678_);
  and (_28683_, _28490_, _28455_);
  and (_28684_, _28455_, _28437_);
  nor (_28685_, _28684_, _28683_);
  and (_28686_, _28598_, _28449_);
  and (_28687_, _28598_, _28490_);
  nor (_28688_, _28687_, _28686_);
  and (_28689_, _28688_, _28685_);
  and (_28690_, _28689_, _28682_);
  and (_28691_, _28690_, _28675_);
  and (_28692_, _28499_, _28449_);
  and (_28693_, _28499_, _28437_);
  nor (_28694_, _28693_, _28692_);
  and (_28695_, _28449_, _28447_);
  and (_28696_, _28509_, _28447_);
  nor (_28697_, _28696_, _28695_);
  and (_28698_, _28697_, _28694_);
  and (_28699_, _28499_, _28490_);
  and (_28700_, _28499_, _28492_);
  nor (_28701_, _28700_, _28699_);
  and (_28702_, _28463_, _28447_);
  and (_28703_, _28499_, _28476_);
  nor (_28704_, _28703_, _28702_);
  and (_28705_, _28704_, _28701_);
  and (_28706_, _28705_, _28698_);
  and (_28707_, _28579_, _28449_);
  and (_28708_, _28492_, _28447_);
  nor (_28709_, _28708_, _28707_);
  and (_28710_, _28579_, _28463_);
  and (_28711_, _28579_, _28509_);
  nor (_28712_, _28711_, _28710_);
  and (_28713_, _28712_, _28709_);
  and (_28714_, _28487_, _28447_);
  and (_28715_, _28470_, _28447_);
  nor (_28716_, _28715_, _28714_);
  and (_28717_, _28447_, _28437_);
  and (_28718_, _28476_, _28447_);
  nor (_28719_, _28718_, _28717_);
  and (_28720_, _28719_, _28716_);
  and (_28721_, _28720_, _28713_);
  and (_28722_, _28721_, _28706_);
  and (_28723_, _28722_, _28691_);
  and (_28724_, _28723_, _28660_);
  and (_28725_, _28724_, _28596_);
  and (_28726_, _28538_, _28476_);
  and (_28727_, _28538_, _28492_);
  nor (_28728_, _28727_, _28726_);
  and (_28729_, _28579_, _28554_);
  and (_28730_, _28538_, _28487_);
  nor (_28731_, _28730_, _28729_);
  and (_28732_, _28731_, _28728_);
  and (_28733_, _28598_, _28446_);
  and (_28734_, _28509_, _28441_);
  nor (_28735_, _28734_, _28733_);
  and (_28736_, _28449_, _28441_);
  and (_28737_, _28490_, _28441_);
  nor (_28738_, _28737_, _28736_);
  and (_28739_, _28738_, _28735_);
  and (_28740_, _28739_, _28732_);
  and (_28741_, _28528_, _28446_);
  and (_28742_, _28528_, _28437_);
  nor (_28743_, _28742_, _28741_);
  and (_28744_, _28598_, _28431_);
  and (_28745_, _28598_, _28479_);
  nor (_28746_, _28745_, _28744_);
  and (_28747_, _28746_, _28743_);
  and (_28748_, _28487_, _28452_);
  and (_28749_, _28441_, _28431_);
  nor (_28750_, _28749_, _28748_);
  and (_28751_, _28479_, _28441_);
  and (_28752_, _28463_, _28441_);
  nor (_28753_, _28752_, _28751_);
  and (_28754_, _28753_, _28750_);
  and (_28755_, _28754_, _28747_);
  and (_28756_, _28755_, _28740_);
  and (_28757_, _28470_, _28452_);
  and (_28758_, _28514_, _28452_);
  nor (_28759_, _28758_, _28757_);
  and (_28760_, _28549_, _28509_);
  and (_28761_, _28554_, _28538_);
  nor (_28762_, _28761_, _28760_);
  and (_28763_, _28762_, _28759_);
  and (_28764_, _28525_, _28434_);
  and (_28765_, _28549_, _28463_);
  nor (_28766_, _28765_, _28764_);
  and (_28767_, _28549_, _28479_);
  and (_28768_, _28549_, _28431_);
  nor (_28769_, _28768_, _28767_);
  and (_28770_, _28769_, _28766_);
  and (_28771_, _28770_, _28763_);
  and (_28772_, _28538_, _28422_);
  and (_28773_, _28476_, _28452_);
  nor (_28774_, _28773_, _28772_);
  and (_28775_, _28538_, _28434_);
  and (_28776_, _28538_, _28470_);
  nor (_28777_, _28776_, _28775_);
  and (_28778_, _28777_, _28774_);
  and (_28779_, _28554_, _28452_);
  and (_28780_, _28492_, _28452_);
  nor (_28781_, _28780_, _28779_);
  and (_28782_, _28452_, _28422_);
  and (_28783_, _28452_, _28434_);
  nor (_28784_, _28783_, _28782_);
  and (_28785_, _28784_, _28781_);
  and (_28786_, _28785_, _28778_);
  and (_28787_, _28786_, _28771_);
  and (_28788_, _28787_, _28756_);
  and (_28789_, _28492_, _28455_);
  and (_28790_, _28598_, _28470_);
  nor (_28791_, _28790_, _28789_);
  and (_28792_, _28554_, _28505_);
  and (_28793_, _28487_, _28455_);
  nor (_28794_, _28793_, _28792_);
  and (_28795_, _28794_, _28791_);
  and (_28796_, _28554_, _28426_);
  and (_28797_, _28514_, _28467_);
  nor (_28798_, _28797_, _28796_);
  and (_28799_, _28479_, _28467_);
  and (_28800_, _28476_, _28455_);
  nor (_28801_, _28800_, _28799_);
  and (_28802_, _28801_, _28798_);
  and (_28803_, _28437_, _28426_);
  and (_28804_, _28490_, _28426_);
  nor (_28805_, _28804_, _28803_);
  and (_28806_, _28492_, _28426_);
  and (_28807_, _28476_, _28426_);
  nor (_28808_, _28807_, _28806_);
  and (_28809_, _28808_, _28805_);
  and (_28810_, _28809_, _28802_);
  and (_28811_, _28810_, _28795_);
  and (_28812_, _28505_, _28437_);
  and (_28813_, _28505_, _28490_);
  nor (_28814_, _28813_, _28812_);
  and (_28815_, _28441_, _28434_);
  and (_28816_, _28538_, _28436_);
  nor (_28817_, _28816_, _28815_);
  and (_28818_, _28817_, _28814_);
  and (_28819_, _28598_, _28509_);
  and (_28820_, _28528_, _28449_);
  nor (_28821_, _28820_, _28819_);
  and (_28822_, _28579_, _28479_);
  and (_28823_, _28463_, _28455_);
  nor (_28824_, _28823_, _28822_);
  and (_28825_, _28824_, _28821_);
  and (_28826_, _28825_, _28818_);
  and (_28827_, _28598_, _28463_);
  and (_28828_, _28528_, _28490_);
  nor (_28829_, _28828_, _28827_);
  and (_28830_, _28487_, _28426_);
  and (_28831_, _28509_, _28426_);
  nor (_28832_, _28831_, _28830_);
  and (_28833_, _28832_, _28829_);
  and (_28834_, _28579_, _28437_);
  and (_28835_, _28579_, _28490_);
  nor (_28836_, _28835_, _28834_);
  and (_28837_, _28538_, _28446_);
  and (_28838_, _28579_, _28431_);
  nor (_28839_, _28838_, _28837_);
  and (_28840_, _28839_, _28836_);
  and (_28841_, _28840_, _28833_);
  and (_28842_, _28841_, _28826_);
  and (_28843_, _28842_, _28811_);
  and (_28844_, _28843_, _28788_);
  and (_28845_, _28544_, _28422_);
  and (_28846_, _28544_, _28449_);
  nor (_28847_, _28846_, _28845_);
  and (_28848_, _28544_, _28434_);
  and (_28849_, _28528_, _28422_);
  nor (_28850_, _28849_, _28848_);
  and (_28851_, _28850_, _28847_);
  and (_28852_, _28544_, _28514_);
  and (_28853_, _28499_, _28446_);
  nor (_28854_, _28853_, _28852_);
  and (_28855_, _28544_, _28470_);
  and (_28856_, _28544_, _28490_);
  nor (_28857_, _28856_, _28855_);
  and (_28858_, _28857_, _28854_);
  and (_28859_, _28858_, _28851_);
  and (_28860_, _28492_, _28461_);
  and (_28861_, _28554_, _28461_);
  nor (_28862_, _28861_, _28860_);
  and (_28863_, _28598_, _28434_);
  and (_28864_, _28598_, _28514_);
  nor (_28865_, _28864_, _28863_);
  and (_28866_, _28865_, _28862_);
  and (_28867_, _28528_, _28434_);
  and (_28868_, _28528_, _28470_);
  nor (_28869_, _28868_, _28867_);
  and (_28870_, _28528_, _28514_);
  and (_28871_, _28554_, _28455_);
  nor (_28872_, _28871_, _28870_);
  and (_28873_, _28872_, _28869_);
  and (_28874_, _28873_, _28866_);
  and (_28875_, _28874_, _28859_);
  and (_28876_, _28514_, _28447_);
  and (_28877_, _28514_, _28455_);
  nor (_28878_, _28877_, _28876_);
  and (_28879_, _28479_, _28447_);
  and (_28880_, _28447_, _28422_);
  nor (_28881_, _28880_, _28879_);
  and (_28882_, _28881_, _28878_);
  and (_28883_, _28514_, _28505_);
  and (_28884_, _28470_, _28455_);
  nor (_28885_, _28884_, _28883_);
  and (_28886_, _28505_, _28434_);
  and (_28887_, _28505_, _28470_);
  nor (_28888_, _28887_, _28886_);
  and (_28889_, _28888_, _28885_);
  and (_28890_, _28889_, _28882_);
  and (_28891_, _28499_, _28463_);
  and (_28892_, _28499_, _28470_);
  nor (_28893_, _28892_, _28891_);
  and (_28894_, _28544_, _28437_);
  and (_28895_, _28499_, _28487_);
  nor (_28896_, _28895_, _28894_);
  and (_28897_, _28896_, _28893_);
  and (_28898_, _28467_, _28446_);
  and (_28899_, _28447_, _28431_);
  nor (_28900_, _28899_, _28898_);
  and (_28901_, _28509_, _28499_);
  and (_28902_, _28490_, _28447_);
  nor (_28903_, _28902_, _28901_);
  and (_28904_, _28903_, _28900_);
  and (_28905_, _28904_, _28897_);
  and (_28906_, _28905_, _28890_);
  and (_28907_, _28906_, _28875_);
  and (_28908_, _28525_, _28487_);
  and (_28909_, _28525_, _28476_);
  nor (_28910_, _28909_, _28908_);
  and (_28911_, _28525_, _28492_);
  and (_28912_, _28554_, _28525_);
  nor (_28913_, _28912_, _28911_);
  and (_28914_, _28913_, _28910_);
  and (_28915_, _28544_, _28463_);
  and (_28916_, _28544_, _28431_);
  nor (_28917_, _28916_, _28915_);
  and (_28918_, _28525_, _28446_);
  and (_28919_, _28549_, _28449_);
  nor (_28920_, _28919_, _28918_);
  and (_28921_, _28920_, _28917_);
  and (_28922_, _28921_, _28914_);
  and (_28923_, _28579_, _28422_);
  and (_28924_, _28579_, _28434_);
  nor (_28925_, _28924_, _28923_);
  and (_28926_, _28538_, _28514_);
  and (_28927_, _28579_, _28470_);
  nor (_28928_, _28927_, _28926_);
  and (_28929_, _28928_, _28925_);
  and (_28930_, _28579_, _28487_);
  and (_28931_, _28579_, _28492_);
  nor (_28932_, _28931_, _28930_);
  and (_28933_, _28579_, _28476_);
  and (_28934_, _28579_, _28514_);
  nor (_28935_, _28934_, _28933_);
  and (_28936_, _28935_, _28932_);
  and (_28937_, _28936_, _28929_);
  and (_28938_, _28937_, _28922_);
  and (_28939_, _28528_, _28479_);
  and (_28940_, _28528_, _28509_);
  nor (_28941_, _28940_, _28939_);
  and (_28942_, _28476_, _28441_);
  and (_28943_, _28528_, _28463_);
  nor (_28944_, _28943_, _28942_);
  and (_28945_, _28944_, _28941_);
  and (_28946_, _28461_, _28449_);
  and (_28947_, _28476_, _28461_);
  nor (_28948_, _28947_, _28946_);
  and (_28949_, _28549_, _28446_);
  and (_28950_, _28509_, _28461_);
  nor (_28951_, _28950_, _28949_);
  and (_28952_, _28951_, _28948_);
  and (_28953_, _28952_, _28945_);
  and (_28954_, _28544_, _28492_);
  and (_28955_, _28470_, _28441_);
  nor (_28956_, _28955_, _28954_);
  and (_28957_, _28554_, _28544_);
  and (_28958_, _28446_, _28441_);
  nor (_28959_, _28958_, _28957_);
  and (_28960_, _28959_, _28956_);
  and (_28961_, _28463_, _28452_);
  and (_28962_, _28492_, _28441_);
  nor (_28963_, _28962_, _28961_);
  and (_28964_, _28514_, _28441_);
  and (_28965_, _28554_, _28441_);
  nor (_28966_, _28965_, _28964_);
  and (_28967_, _28966_, _28963_);
  and (_28968_, _28967_, _28960_);
  and (_28969_, _28968_, _28953_);
  and (_28970_, _28969_, _28938_);
  and (_28971_, _28970_, _28907_);
  and (_28972_, _28971_, _28844_);
  and (_28973_, _28972_, _28725_);
  and (_28974_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  not (_28975_, _28974_);
  and (_28976_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_28977_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor (_28978_, _28977_, _28976_);
  and (_28979_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  and (_28980_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor (_28981_, _28980_, _28979_);
  and (_28982_, _28981_, _28978_);
  and (_28983_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_28984_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor (_28985_, _28984_, _28983_);
  and (_28986_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  and (_28987_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nor (_28988_, _28987_, _28986_);
  and (_28989_, _28988_, _28985_);
  and (_28990_, _28989_, _28982_);
  and (_28991_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  and (_28992_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nor (_28993_, _28992_, _28991_);
  and (_28994_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_28995_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nor (_28996_, _28995_, _28994_);
  and (_28997_, _28996_, _28993_);
  and (_28998_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  and (_28999_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nor (_29000_, _28999_, _28998_);
  and (_29001_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_29002_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor (_29003_, _29002_, _29001_);
  and (_29004_, _29003_, _29000_);
  and (_29005_, _29004_, _28997_);
  and (_29006_, _29005_, _28990_);
  and (_29007_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_29008_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor (_29009_, _29008_, _29007_);
  and (_29010_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  and (_29011_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nor (_29012_, _29011_, _29010_);
  and (_29013_, _29012_, _29009_);
  and (_29014_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  and (_29015_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nor (_29016_, _29015_, _29014_);
  and (_29017_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_29018_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nor (_29019_, _29018_, _29017_);
  and (_29020_, _29019_, _29016_);
  and (_29021_, _29020_, _29013_);
  and (_29022_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_29023_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nor (_29024_, _29023_, _29022_);
  and (_29025_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  and (_29026_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nor (_29027_, _29026_, _29025_);
  and (_29028_, _29027_, _29024_);
  and (_29029_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_29030_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nor (_29031_, _29030_, _29029_);
  and (_29032_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  and (_29033_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor (_29034_, _29033_, _29032_);
  and (_29035_, _29034_, _29031_);
  and (_29036_, _29035_, _29028_);
  and (_29037_, _29036_, _29021_);
  and (_29038_, _29037_, _29006_);
  and (_29039_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_29040_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nor (_29041_, _29040_, _29039_);
  and (_29042_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and (_29043_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor (_29044_, _29043_, _29042_);
  and (_29045_, _29044_, _29041_);
  and (_29046_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_29047_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor (_29048_, _29047_, _29046_);
  and (_29049_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and (_29050_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nor (_29051_, _29050_, _29049_);
  and (_29052_, _29051_, _29048_);
  and (_29053_, _29052_, _29045_);
  and (_29054_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and (_29055_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nor (_29056_, _29055_, _29054_);
  and (_29057_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_29058_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nor (_29059_, _29058_, _29057_);
  and (_29060_, _29059_, _29056_);
  and (_29061_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and (_29062_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nor (_29063_, _29062_, _29061_);
  and (_29064_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_29065_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor (_29066_, _29065_, _29064_);
  and (_29067_, _29066_, _29063_);
  and (_29068_, _29067_, _29060_);
  and (_29069_, _29068_, _29053_);
  and (_29070_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  and (_29071_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor (_29072_, _29071_, _29070_);
  and (_29073_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  and (_29074_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor (_29075_, _29074_, _29073_);
  and (_29076_, _29075_, _29072_);
  and (_29077_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  and (_29078_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor (_29079_, _29078_, _29077_);
  and (_29080_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_29081_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nor (_29082_, _29081_, _29080_);
  and (_29083_, _29082_, _29079_);
  and (_29084_, _29083_, _29076_);
  and (_29085_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_29086_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nor (_29087_, _29086_, _29085_);
  and (_29088_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  and (_29089_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nor (_29090_, _29089_, _29088_);
  and (_29091_, _29090_, _29087_);
  and (_29092_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_29093_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nor (_29094_, _29093_, _29092_);
  and (_29095_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  and (_29096_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nor (_29097_, _29096_, _29095_);
  and (_29098_, _29097_, _29094_);
  and (_29099_, _29098_, _29091_);
  and (_29100_, _29099_, _29084_);
  and (_29101_, _29100_, _29069_);
  and (_29102_, _29101_, _29038_);
  and (_29103_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  and (_29104_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nor (_29105_, _29104_, _29103_);
  and (_29106_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_29107_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nor (_29108_, _29107_, _29106_);
  and (_29109_, _29108_, _29105_);
  and (_29110_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  and (_29111_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nor (_29112_, _29111_, _29110_);
  and (_29113_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_29114_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nor (_29115_, _29114_, _29113_);
  and (_29116_, _29115_, _29112_);
  and (_29117_, _29116_, _29109_);
  and (_29118_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_29119_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor (_29120_, _29119_, _29118_);
  and (_29121_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  and (_29122_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nor (_29123_, _29122_, _29121_);
  and (_29124_, _29123_, _29120_);
  and (_29125_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_29126_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor (_29127_, _29126_, _29125_);
  and (_29128_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  and (_29129_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nor (_29130_, _29129_, _29128_);
  and (_29131_, _29130_, _29127_);
  and (_29132_, _29131_, _29124_);
  and (_29133_, _29132_, _29117_);
  and (_29134_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and (_29135_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nor (_29136_, _29135_, _29134_);
  and (_29137_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_29138_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nor (_29139_, _29138_, _29137_);
  and (_29140_, _29139_, _29136_);
  and (_29141_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_29142_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nor (_29143_, _29142_, _29141_);
  and (_29144_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and (_29145_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nor (_29146_, _29145_, _29144_);
  and (_29147_, _29146_, _29143_);
  and (_29148_, _29147_, _29140_);
  and (_29149_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_29150_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nor (_29151_, _29150_, _29149_);
  and (_29152_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_29153_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nor (_29154_, _29153_, _29152_);
  and (_29155_, _29154_, _29151_);
  and (_29156_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_29157_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nor (_29158_, _29157_, _29156_);
  and (_29159_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  and (_29160_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nor (_29161_, _29160_, _29159_);
  and (_29162_, _29161_, _29158_);
  and (_29163_, _29162_, _29155_);
  and (_29164_, _29163_, _29148_);
  and (_29165_, _29164_, _29133_);
  and (_29166_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_29167_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nor (_29168_, _29167_, _29166_);
  and (_29169_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  and (_29170_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nor (_29171_, _29170_, _29169_);
  and (_29172_, _29171_, _29168_);
  and (_29173_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_29174_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nor (_29175_, _29174_, _29173_);
  and (_29176_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  and (_29177_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nor (_29178_, _29177_, _29176_);
  and (_29179_, _29178_, _29175_);
  and (_29180_, _29179_, _29172_);
  and (_29181_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  and (_29182_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nor (_29183_, _29182_, _29181_);
  and (_29184_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  and (_29185_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nor (_29186_, _29185_, _29184_);
  and (_29187_, _29186_, _29183_);
  and (_29188_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  and (_29189_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nor (_29190_, _29189_, _29188_);
  and (_29191_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_29192_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor (_29193_, _29192_, _29191_);
  and (_29194_, _29193_, _29190_);
  and (_29195_, _29194_, _29187_);
  and (_29196_, _29195_, _29180_);
  and (_29197_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_29198_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor (_29199_, _29198_, _29197_);
  and (_29200_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  and (_29201_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor (_29202_, _29201_, _29200_);
  and (_29203_, _29202_, _29199_);
  and (_29204_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_29205_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor (_29206_, _29205_, _29204_);
  and (_29207_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_29208_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor (_29209_, _29208_, _29207_);
  and (_29210_, _29209_, _29206_);
  and (_29211_, _29210_, _29203_);
  and (_29212_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  and (_29213_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nor (_29214_, _29213_, _29212_);
  and (_29215_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_29216_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nor (_29217_, _29216_, _29215_);
  and (_29218_, _29217_, _29214_);
  and (_29219_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  and (_29220_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nor (_29221_, _29220_, _29219_);
  and (_29222_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_29223_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor (_29224_, _29223_, _29222_);
  and (_29225_, _29224_, _29221_);
  and (_29226_, _29225_, _29218_);
  and (_29227_, _29226_, _29211_);
  and (_29228_, _29227_, _29196_);
  and (_29229_, _29228_, _29165_);
  and (_29230_, _29229_, _29102_);
  and (_29231_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  and (_29232_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor (_29233_, _29232_, _29231_);
  and (_29234_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_29235_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nor (_29236_, _29235_, _29234_);
  and (_29237_, _29236_, _29233_);
  and (_29238_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  and (_29239_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nor (_29240_, _29239_, _29238_);
  and (_29241_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_29242_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nor (_29243_, _29242_, _29241_);
  and (_29244_, _29243_, _29240_);
  and (_29245_, _29244_, _29237_);
  and (_29246_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_29247_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nor (_29248_, _29247_, _29246_);
  and (_29249_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  and (_29250_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nor (_29251_, _29250_, _29249_);
  and (_29252_, _29251_, _29248_);
  and (_29253_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_29254_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nor (_29255_, _29254_, _29253_);
  and (_29256_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  and (_29257_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nor (_29258_, _29257_, _29256_);
  and (_29259_, _29258_, _29255_);
  and (_29260_, _29259_, _29252_);
  and (_29261_, _29260_, _29245_);
  and (_29262_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_29263_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor (_29264_, _29263_, _29262_);
  and (_29265_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  and (_29266_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor (_29267_, _29266_, _29265_);
  and (_29268_, _29267_, _29264_);
  and (_29269_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_29270_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor (_29271_, _29270_, _29269_);
  and (_29272_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  and (_29273_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nor (_29274_, _29273_, _29272_);
  and (_29275_, _29274_, _29271_);
  and (_29276_, _29275_, _29268_);
  and (_29277_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  and (_29278_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nor (_29279_, _29278_, _29277_);
  and (_29280_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_29281_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nor (_29282_, _29281_, _29280_);
  and (_29283_, _29282_, _29279_);
  and (_29284_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_29285_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nor (_29286_, _29285_, _29284_);
  and (_29287_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  and (_29288_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nor (_29289_, _29288_, _29287_);
  and (_29290_, _29289_, _29286_);
  and (_29291_, _29290_, _29283_);
  and (_29292_, _29291_, _29276_);
  and (_29293_, _29292_, _29261_);
  and (_29294_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and (_29295_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nor (_29296_, _29295_, _29294_);
  and (_29297_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  and (_29298_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor (_29299_, _29298_, _29297_);
  and (_29300_, _29299_, _29296_);
  and (_29301_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and (_29302_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor (_29303_, _29302_, _29301_);
  and (_29304_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  and (_29305_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nor (_29306_, _29305_, _29304_);
  and (_29307_, _29306_, _29303_);
  and (_29308_, _29307_, _29300_);
  and (_29309_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and (_29310_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nor (_29311_, _29310_, _29309_);
  and (_29312_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  and (_29313_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nor (_29314_, _29313_, _29312_);
  and (_29315_, _29314_, _29311_);
  and (_29316_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  and (_29317_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nor (_29318_, _29317_, _29316_);
  and (_29319_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and (_29320_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor (_29321_, _29320_, _29319_);
  and (_29322_, _29321_, _29318_);
  and (_29323_, _29322_, _29315_);
  and (_29324_, _29323_, _29308_);
  and (_29325_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_29326_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor (_29327_, _29326_, _29325_);
  and (_29328_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  and (_29329_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor (_29330_, _29329_, _29328_);
  and (_29331_, _29330_, _29327_);
  and (_29332_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_29333_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor (_29334_, _29333_, _29332_);
  and (_29335_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_29336_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor (_29337_, _29336_, _29335_);
  and (_29338_, _29337_, _29334_);
  and (_29339_, _29338_, _29331_);
  and (_29340_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  and (_29341_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nor (_29342_, _29341_, _29340_);
  and (_29343_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_29344_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nor (_29345_, _29344_, _29343_);
  and (_29346_, _29345_, _29342_);
  and (_29347_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  and (_29348_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nor (_29349_, _29348_, _29347_);
  and (_29350_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  and (_29351_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nor (_29352_, _29351_, _29350_);
  and (_29353_, _29352_, _29349_);
  and (_29354_, _29353_, _29346_);
  and (_29355_, _29354_, _29339_);
  and (_29356_, _29355_, _29324_);
  and (_29357_, _29356_, _29293_);
  and (_29358_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  and (_29359_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nor (_29360_, _29359_, _29358_);
  and (_29361_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_29362_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nor (_29363_, _29362_, _29361_);
  and (_29364_, _29363_, _29360_);
  and (_29365_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  and (_29366_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nor (_29367_, _29366_, _29365_);
  and (_29368_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_29369_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nor (_29370_, _29369_, _29368_);
  and (_29371_, _29370_, _29367_);
  and (_29372_, _29371_, _29364_);
  and (_29373_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_29374_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nor (_29375_, _29374_, _29373_);
  and (_29376_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_29377_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nor (_29378_, _29377_, _29376_);
  and (_29379_, _29378_, _29375_);
  and (_29380_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_29381_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor (_29382_, _29381_, _29380_);
  and (_29383_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  and (_29384_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor (_29385_, _29384_, _29383_);
  and (_29386_, _29385_, _29382_);
  and (_29387_, _29386_, _29379_);
  and (_29388_, _29387_, _29372_);
  and (_29389_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_29390_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nor (_29391_, _29390_, _29389_);
  and (_29392_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  and (_29393_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nor (_29394_, _29393_, _29392_);
  and (_29395_, _29394_, _29391_);
  and (_29396_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_29397_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nor (_29398_, _29397_, _29396_);
  and (_29399_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  and (_29400_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor (_29401_, _29400_, _29399_);
  and (_29402_, _29401_, _29398_);
  and (_29403_, _29402_, _29395_);
  and (_29404_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  and (_29405_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nor (_29406_, _29405_, _29404_);
  and (_29407_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  and (_29408_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor (_29409_, _29408_, _29407_);
  and (_29410_, _29409_, _29406_);
  and (_29411_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  and (_29412_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nor (_29413_, _29412_, _29411_);
  and (_29414_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_29415_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor (_29416_, _29415_, _29414_);
  and (_29417_, _29416_, _29413_);
  and (_29418_, _29417_, _29410_);
  and (_29419_, _29418_, _29403_);
  and (_29420_, _29419_, _29388_);
  and (_29421_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  and (_29422_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nor (_29423_, _29422_, _29421_);
  and (_29424_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_29425_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nor (_29426_, _29425_, _29424_);
  and (_29427_, _29426_, _29423_);
  and (_29428_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  and (_29429_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nor (_29430_, _29429_, _29428_);
  and (_29431_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_29432_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nor (_29433_, _29432_, _29431_);
  and (_29434_, _29433_, _29430_);
  and (_29435_, _29434_, _29427_);
  and (_29436_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_29437_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nor (_29438_, _29437_, _29436_);
  and (_29439_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  and (_29440_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor (_29441_, _29440_, _29439_);
  and (_29442_, _29441_, _29438_);
  and (_29443_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_29444_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nor (_29445_, _29444_, _29443_);
  and (_29446_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_29447_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor (_29448_, _29447_, _29446_);
  and (_29449_, _29448_, _29445_);
  and (_29450_, _29449_, _29442_);
  and (_29451_, _29450_, _29435_);
  and (_29452_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_29453_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_29454_, _29453_, _29452_);
  and (_29455_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_29456_, _28538_, _28479_);
  and (_29457_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_29458_, _29457_, _29455_);
  and (_29459_, _29458_, _29454_);
  and (_29460_, _28538_, _28490_);
  and (_29461_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_29462_, _28538_, _28449_);
  and (_29463_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_29464_, _28538_, _28437_);
  and (_29465_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_29466_, _29465_, _29463_);
  nor (_29467_, _29466_, _29461_);
  and (_29468_, _29467_, _29459_);
  and (_29469_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_29470_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_29471_, _29470_, _29469_);
  and (_29472_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_29473_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_29474_, _29473_, _29472_);
  and (_29475_, _29474_, _29471_);
  and (_29476_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_29477_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_29478_, _29477_, _29476_);
  and (_29479_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_29480_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_29481_, _29480_, _29479_);
  and (_29482_, _29481_, _29478_);
  and (_29483_, _29482_, _29475_);
  and (_29484_, _29483_, _29468_);
  and (_29485_, _29484_, _29451_);
  and (_29486_, _29485_, _29420_);
  and (_29487_, _29486_, _29357_);
  and (_29488_, _29487_, _29230_);
  and (_29489_, _29488_, _28975_);
  and (_29490_, iram_op1_reg[0], iram_op1_reg[1]);
  and (_29491_, _29490_, iram_op1_reg[2]);
  nor (_29492_, _29490_, iram_op1_reg[2]);
  nor (_29493_, _29492_, _29491_);
  nor (_29494_, _29493_, _29489_);
  and (_29495_, _29493_, _29489_);
  or (_29496_, _29495_, _29494_);
  and (_29497_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  not (_29498_, _29497_);
  and (_29499_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  and (_29500_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor (_29501_, _29500_, _29499_);
  and (_29502_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_29503_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nor (_29504_, _29503_, _29502_);
  and (_29505_, _29504_, _29501_);
  and (_29506_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_29507_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor (_29508_, _29507_, _29506_);
  and (_29509_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_29510_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor (_29511_, _29510_, _29509_);
  and (_29512_, _29511_, _29508_);
  and (_29513_, _29512_, _29505_);
  and (_29514_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_29515_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nor (_29516_, _29515_, _29514_);
  and (_29517_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  and (_29518_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nor (_29519_, _29518_, _29517_);
  and (_29520_, _29519_, _29516_);
  and (_29521_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  and (_29522_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nor (_29523_, _29522_, _29521_);
  and (_29524_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_29525_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor (_29526_, _29525_, _29524_);
  and (_29527_, _29526_, _29523_);
  and (_29528_, _29527_, _29520_);
  and (_29529_, _29528_, _29513_);
  and (_29530_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_29531_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nor (_29532_, _29531_, _29530_);
  and (_29533_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  and (_29534_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nor (_29535_, _29534_, _29533_);
  and (_29536_, _29535_, _29532_);
  and (_29537_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_29538_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nor (_29539_, _29538_, _29537_);
  and (_29540_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and (_29541_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nor (_29542_, _29541_, _29540_);
  and (_29543_, _29542_, _29539_);
  and (_29544_, _29543_, _29536_);
  and (_29545_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  and (_29546_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nor (_29547_, _29546_, _29545_);
  and (_29548_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  and (_29549_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nor (_29550_, _29549_, _29548_);
  and (_29551_, _29550_, _29547_);
  and (_29552_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  and (_29553_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nor (_29554_, _29553_, _29552_);
  and (_29555_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_29556_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nor (_29557_, _29556_, _29555_);
  and (_29558_, _29557_, _29554_);
  and (_29559_, _29558_, _29551_);
  and (_29560_, _29559_, _29544_);
  and (_29561_, _29560_, _29529_);
  and (_29562_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_29563_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor (_29564_, _29563_, _29562_);
  and (_29565_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and (_29566_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor (_29567_, _29566_, _29565_);
  and (_29568_, _29567_, _29564_);
  and (_29569_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_29570_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor (_29571_, _29570_, _29569_);
  and (_29572_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_29573_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nor (_29574_, _29573_, _29572_);
  and (_29575_, _29574_, _29571_);
  and (_29576_, _29575_, _29568_);
  and (_29577_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and (_29578_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nor (_29579_, _29578_, _29577_);
  and (_29580_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_29581_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nor (_29582_, _29581_, _29580_);
  and (_29583_, _29582_, _29579_);
  and (_29584_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and (_29585_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nor (_29586_, _29585_, _29584_);
  and (_29587_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_29588_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor (_29589_, _29588_, _29587_);
  and (_29590_, _29589_, _29586_);
  and (_29591_, _29590_, _29583_);
  and (_29592_, _29591_, _29576_);
  and (_29593_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  and (_29594_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nor (_29595_, _29594_, _29593_);
  and (_29596_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_29597_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor (_29598_, _29597_, _29596_);
  and (_29599_, _29598_, _29595_);
  and (_29600_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  and (_29601_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nor (_29602_, _29601_, _29600_);
  and (_29603_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  and (_29604_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor (_29605_, _29604_, _29603_);
  and (_29606_, _29605_, _29602_);
  and (_29607_, _29606_, _29599_);
  and (_29608_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_29609_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nor (_29610_, _29609_, _29608_);
  and (_29611_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  and (_29612_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nor (_29613_, _29612_, _29611_);
  and (_29614_, _29613_, _29610_);
  and (_29615_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_29616_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nor (_29617_, _29616_, _29615_);
  and (_29618_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  and (_29619_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor (_29620_, _29619_, _29618_);
  and (_29621_, _29620_, _29617_);
  and (_29622_, _29621_, _29614_);
  and (_29623_, _29622_, _29607_);
  and (_29624_, _29623_, _29592_);
  and (_29625_, _29624_, _29561_);
  and (_29626_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and (_29627_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor (_29628_, _29627_, _29626_);
  and (_29629_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_29630_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor (_29631_, _29630_, _29629_);
  and (_29632_, _29631_, _29628_);
  and (_29633_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_29634_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nor (_29635_, _29634_, _29633_);
  and (_29636_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_29637_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nor (_29638_, _29637_, _29636_);
  and (_29639_, _29638_, _29635_);
  and (_29640_, _29639_, _29632_);
  and (_29641_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_29642_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nor (_29643_, _29642_, _29641_);
  and (_29644_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_29645_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor (_29646_, _29645_, _29644_);
  and (_29647_, _29646_, _29643_);
  and (_29648_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_29649_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nor (_29650_, _29649_, _29648_);
  and (_29651_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and (_29652_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nor (_29653_, _29652_, _29651_);
  and (_29654_, _29653_, _29650_);
  and (_29655_, _29654_, _29647_);
  and (_29656_, _29655_, _29640_);
  and (_29657_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  and (_29658_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor (_29659_, _29658_, _29657_);
  and (_29660_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_29661_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor (_29662_, _29661_, _29660_);
  and (_29663_, _29662_, _29659_);
  and (_29664_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_29665_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor (_29666_, _29665_, _29664_);
  and (_29667_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_29668_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nor (_29669_, _29668_, _29667_);
  and (_29670_, _29669_, _29666_);
  and (_29671_, _29670_, _29663_);
  and (_29672_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  and (_29673_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nor (_29674_, _29673_, _29672_);
  and (_29675_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_29676_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nor (_29677_, _29676_, _29675_);
  and (_29678_, _29677_, _29674_);
  and (_29679_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_29680_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor (_29681_, _29680_, _29679_);
  and (_29682_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  and (_29683_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nor (_29684_, _29683_, _29682_);
  and (_29685_, _29684_, _29681_);
  and (_29686_, _29685_, _29678_);
  and (_29687_, _29686_, _29671_);
  and (_29688_, _29687_, _29656_);
  and (_29689_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_29690_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor (_29691_, _29690_, _29689_);
  and (_29692_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  and (_29693_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor (_29694_, _29693_, _29692_);
  and (_29695_, _29694_, _29691_);
  and (_29696_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_29697_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor (_29698_, _29697_, _29696_);
  and (_29699_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  and (_29700_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nor (_29701_, _29700_, _29699_);
  and (_29702_, _29701_, _29698_);
  and (_29703_, _29702_, _29695_);
  and (_29704_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  and (_29705_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nor (_29706_, _29705_, _29704_);
  and (_29707_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_29708_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nor (_29709_, _29708_, _29707_);
  and (_29710_, _29709_, _29706_);
  and (_29711_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  and (_29712_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nor (_29713_, _29712_, _29711_);
  and (_29714_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_29715_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nor (_29716_, _29715_, _29714_);
  and (_29717_, _29716_, _29713_);
  and (_29718_, _29717_, _29710_);
  and (_29719_, _29718_, _29703_);
  and (_29720_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  and (_29721_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nor (_29722_, _29721_, _29720_);
  and (_29723_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_29724_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nor (_29725_, _29724_, _29723_);
  and (_29726_, _29725_, _29722_);
  and (_29727_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_29728_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nor (_29729_, _29728_, _29727_);
  and (_29730_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  and (_29731_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nor (_29732_, _29731_, _29730_);
  and (_29733_, _29732_, _29729_);
  and (_29734_, _29733_, _29726_);
  and (_29735_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  and (_29736_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor (_29737_, _29736_, _29735_);
  and (_29738_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  and (_29739_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nor (_29740_, _29739_, _29738_);
  and (_29741_, _29740_, _29737_);
  and (_29742_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  and (_29743_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor (_29744_, _29743_, _29742_);
  and (_29745_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_29746_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nor (_29747_, _29746_, _29745_);
  and (_29748_, _29747_, _29744_);
  and (_29749_, _29748_, _29741_);
  and (_29750_, _29749_, _29734_);
  and (_29751_, _29750_, _29719_);
  and (_29752_, _29751_, _29688_);
  and (_29753_, _29752_, _29625_);
  and (_29754_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  and (_29755_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor (_29756_, _29755_, _29754_);
  and (_29757_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_29758_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nor (_29759_, _29758_, _29757_);
  and (_29760_, _29759_, _29756_);
  and (_29761_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  and (_29762_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nor (_29763_, _29762_, _29761_);
  and (_29764_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_29765_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nor (_29766_, _29765_, _29764_);
  and (_29767_, _29766_, _29763_);
  and (_29768_, _29767_, _29760_);
  and (_29769_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_29770_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nor (_29771_, _29770_, _29769_);
  and (_29772_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  and (_29773_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor (_29774_, _29773_, _29772_);
  and (_29775_, _29774_, _29771_);
  and (_29776_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_29777_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nor (_29778_, _29777_, _29776_);
  and (_29779_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  and (_29780_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nor (_29781_, _29780_, _29779_);
  and (_29782_, _29781_, _29778_);
  and (_29783_, _29782_, _29775_);
  and (_29784_, _29783_, _29768_);
  and (_29785_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  and (_29786_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor (_29787_, _29786_, _29785_);
  and (_29788_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_29789_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor (_29790_, _29789_, _29788_);
  and (_29791_, _29790_, _29787_);
  and (_29792_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_29793_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor (_29794_, _29793_, _29792_);
  and (_29795_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_29796_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor (_29797_, _29796_, _29795_);
  and (_29798_, _29797_, _29794_);
  and (_29799_, _29798_, _29791_);
  and (_29800_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  and (_29801_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nor (_29802_, _29801_, _29800_);
  and (_29803_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_29804_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nor (_29805_, _29804_, _29803_);
  and (_29806_, _29805_, _29802_);
  and (_29807_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  and (_29808_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nor (_29809_, _29808_, _29807_);
  and (_29810_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_29811_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nor (_29812_, _29811_, _29810_);
  and (_29813_, _29812_, _29809_);
  and (_29814_, _29813_, _29806_);
  and (_29815_, _29814_, _29799_);
  and (_29816_, _29815_, _29784_);
  and (_29817_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_29818_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor (_29819_, _29818_, _29817_);
  and (_29820_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  and (_29821_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor (_29822_, _29821_, _29820_);
  and (_29823_, _29822_, _29819_);
  and (_29824_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_29825_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor (_29826_, _29825_, _29824_);
  and (_29827_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_29828_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor (_29829_, _29828_, _29827_);
  and (_29830_, _29829_, _29826_);
  and (_29831_, _29830_, _29823_);
  and (_29832_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  and (_29833_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nor (_29834_, _29833_, _29832_);
  and (_29835_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_29836_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nor (_29837_, _29836_, _29835_);
  and (_29838_, _29837_, _29834_);
  and (_29839_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  and (_29840_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nor (_29841_, _29840_, _29839_);
  and (_29842_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_29843_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nor (_29844_, _29843_, _29842_);
  and (_29845_, _29844_, _29841_);
  and (_29846_, _29845_, _29838_);
  and (_29847_, _29846_, _29831_);
  and (_29848_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  and (_29849_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor (_29850_, _29849_, _29848_);
  and (_29851_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_29852_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nor (_29853_, _29852_, _29851_);
  and (_29854_, _29853_, _29850_);
  and (_29855_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  and (_29856_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nor (_29857_, _29856_, _29855_);
  and (_29858_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  and (_29859_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nor (_29860_, _29859_, _29858_);
  and (_29861_, _29860_, _29857_);
  and (_29862_, _29861_, _29854_);
  and (_29863_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_29864_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nor (_29865_, _29864_, _29863_);
  and (_29866_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  and (_29867_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nor (_29868_, _29867_, _29866_);
  and (_29869_, _29868_, _29865_);
  and (_29870_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_29871_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nor (_29872_, _29871_, _29870_);
  and (_29873_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  and (_29874_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nor (_29875_, _29874_, _29873_);
  and (_29876_, _29875_, _29872_);
  and (_29877_, _29876_, _29869_);
  and (_29878_, _29877_, _29862_);
  and (_29879_, _29878_, _29847_);
  and (_29880_, _29879_, _29816_);
  and (_29881_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_29882_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nor (_29883_, _29882_, _29881_);
  and (_29884_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  and (_29885_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor (_29886_, _29885_, _29884_);
  and (_29887_, _29886_, _29883_);
  and (_29888_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_29889_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor (_29890_, _29889_, _29888_);
  and (_29891_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  and (_29892_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nor (_29893_, _29892_, _29891_);
  and (_29894_, _29893_, _29890_);
  and (_29895_, _29894_, _29887_);
  and (_29896_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  and (_29897_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nor (_29898_, _29897_, _29896_);
  and (_29899_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_29900_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor (_29901_, _29900_, _29899_);
  and (_29902_, _29901_, _29898_);
  and (_29903_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  and (_29904_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nor (_29905_, _29904_, _29903_);
  and (_29906_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_29907_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nor (_29908_, _29907_, _29906_);
  and (_29909_, _29908_, _29905_);
  and (_29910_, _29909_, _29902_);
  and (_29911_, _29910_, _29895_);
  and (_29912_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_29913_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nor (_29914_, _29913_, _29912_);
  and (_29915_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  and (_29916_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nor (_29917_, _29916_, _29915_);
  and (_29918_, _29917_, _29914_);
  and (_29919_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_29920_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nor (_29921_, _29920_, _29919_);
  and (_29922_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  and (_29923_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor (_29924_, _29923_, _29922_);
  and (_29925_, _29924_, _29921_);
  and (_29926_, _29925_, _29918_);
  and (_29927_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  and (_29928_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nor (_29929_, _29928_, _29927_);
  and (_29930_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  and (_29931_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nor (_29932_, _29931_, _29930_);
  and (_29933_, _29932_, _29929_);
  and (_29934_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  and (_29935_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor (_29936_, _29935_, _29934_);
  and (_29937_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_29938_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nor (_29939_, _29938_, _29937_);
  and (_29940_, _29939_, _29936_);
  and (_29941_, _29940_, _29933_);
  and (_29942_, _29941_, _29926_);
  and (_29943_, _29942_, _29911_);
  and (_29944_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_29945_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor (_29946_, _29945_, _29944_);
  and (_29947_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  and (_29948_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor (_29949_, _29948_, _29947_);
  and (_29950_, _29949_, _29946_);
  and (_29951_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_29952_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor (_29953_, _29952_, _29951_);
  and (_29954_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  and (_29955_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nor (_29956_, _29955_, _29954_);
  and (_29957_, _29956_, _29953_);
  and (_29958_, _29957_, _29950_);
  and (_29959_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  and (_29960_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nor (_29961_, _29960_, _29959_);
  and (_29962_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_29963_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nor (_29964_, _29963_, _29962_);
  and (_29965_, _29964_, _29961_);
  and (_29966_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  and (_29967_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nor (_29968_, _29967_, _29966_);
  and (_29969_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_29970_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nor (_29971_, _29970_, _29969_);
  and (_29972_, _29971_, _29968_);
  and (_29973_, _29972_, _29965_);
  and (_29974_, _29973_, _29958_);
  and (_29975_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_29976_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_29977_, _29976_, _29975_);
  and (_29978_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_29979_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_29980_, _29979_, _29978_);
  and (_29981_, _29980_, _29977_);
  and (_29982_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_29983_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_29984_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_29985_, _29984_, _29983_);
  nor (_29986_, _29985_, _29982_);
  and (_29987_, _29986_, _29981_);
  and (_29988_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_29989_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_29990_, _29989_, _29988_);
  and (_29991_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_29992_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_29993_, _29992_, _29991_);
  and (_29994_, _29993_, _29990_);
  and (_29995_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_29996_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_29997_, _29996_, _29995_);
  and (_29998_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_29999_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_30000_, _29999_, _29998_);
  and (_30001_, _30000_, _29997_);
  and (_30002_, _30001_, _29994_);
  and (_30003_, _30002_, _29987_);
  and (_30004_, _30003_, _29974_);
  and (_30005_, _30004_, _29943_);
  and (_30006_, _30005_, _29880_);
  and (_30007_, _30006_, _29753_);
  and (_30008_, _30007_, _29498_);
  and (_30009_, _29491_, iram_op1_reg[3]);
  and (_30010_, _30009_, iram_op1_reg[4]);
  nor (_30011_, _30009_, iram_op1_reg[4]);
  nor (_30012_, _30011_, _30010_);
  and (_30013_, _30012_, _30008_);
  nor (_30014_, _30012_, _30008_);
  or (_30015_, _30014_, _30013_);
  and (_30016_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  not (_30017_, _30016_);
  and (_30018_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_30019_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor (_30020_, _30019_, _30018_);
  and (_30021_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  and (_30022_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor (_30023_, _30022_, _30021_);
  and (_30024_, _30023_, _30020_);
  and (_30025_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_30026_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor (_30027_, _30026_, _30025_);
  and (_30028_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  and (_30029_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nor (_30030_, _30029_, _30028_);
  and (_30031_, _30030_, _30027_);
  and (_30032_, _30031_, _30024_);
  and (_30033_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  and (_30034_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nor (_30035_, _30034_, _30033_);
  and (_30036_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_30037_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nor (_30038_, _30037_, _30036_);
  and (_30039_, _30038_, _30035_);
  and (_30040_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  and (_30041_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nor (_30042_, _30041_, _30040_);
  and (_30043_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_30044_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nor (_30045_, _30044_, _30043_);
  and (_30046_, _30045_, _30042_);
  and (_30047_, _30046_, _30039_);
  and (_30048_, _30047_, _30032_);
  and (_30049_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_30050_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nor (_30051_, _30050_, _30049_);
  and (_30052_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  and (_30053_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nor (_30054_, _30053_, _30052_);
  and (_30055_, _30054_, _30051_);
  and (_30056_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_30057_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nor (_30058_, _30057_, _30056_);
  and (_30059_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and (_30060_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nor (_30061_, _30060_, _30059_);
  and (_30062_, _30061_, _30058_);
  and (_30063_, _30062_, _30055_);
  and (_30064_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  and (_30065_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor (_30066_, _30065_, _30064_);
  and (_30067_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  and (_30068_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nor (_30069_, _30068_, _30067_);
  and (_30070_, _30069_, _30066_);
  and (_30071_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  and (_30072_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor (_30073_, _30072_, _30071_);
  and (_30074_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_30075_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor (_30076_, _30075_, _30074_);
  and (_30077_, _30076_, _30073_);
  and (_30078_, _30077_, _30070_);
  and (_30079_, _30078_, _30063_);
  and (_30080_, _30079_, _30048_);
  and (_30081_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_30082_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nor (_30083_, _30082_, _30081_);
  and (_30084_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and (_30085_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor (_30086_, _30085_, _30084_);
  and (_30087_, _30086_, _30083_);
  and (_30088_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_30089_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nor (_30090_, _30089_, _30088_);
  and (_30091_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_30092_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor (_30093_, _30092_, _30091_);
  and (_30094_, _30093_, _30090_);
  and (_30095_, _30094_, _30087_);
  and (_30096_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and (_30097_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nor (_30098_, _30097_, _30096_);
  and (_30099_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_30100_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nor (_30101_, _30100_, _30099_);
  and (_30102_, _30101_, _30098_);
  and (_30103_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and (_30104_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nor (_30105_, _30104_, _30103_);
  and (_30106_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_30107_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nor (_30108_, _30107_, _30106_);
  and (_30109_, _30108_, _30105_);
  and (_30110_, _30109_, _30102_);
  and (_30111_, _30110_, _30095_);
  and (_30112_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_30113_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nor (_30114_, _30113_, _30112_);
  and (_30115_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  and (_30116_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nor (_30117_, _30116_, _30115_);
  and (_30118_, _30117_, _30114_);
  and (_30119_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_30120_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nor (_30121_, _30120_, _30119_);
  and (_30122_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  and (_30123_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nor (_30124_, _30123_, _30122_);
  and (_30125_, _30124_, _30121_);
  and (_30126_, _30125_, _30118_);
  and (_30127_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  and (_30128_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nor (_30129_, _30128_, _30127_);
  and (_30130_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_30131_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nor (_30132_, _30131_, _30130_);
  and (_30133_, _30132_, _30129_);
  and (_30134_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  and (_30135_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor (_30136_, _30135_, _30134_);
  and (_30137_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  and (_30138_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nor (_30139_, _30138_, _30137_);
  and (_30140_, _30139_, _30136_);
  and (_30141_, _30140_, _30133_);
  and (_30142_, _30141_, _30126_);
  and (_30143_, _30142_, _30111_);
  and (_30144_, _30143_, _30080_);
  and (_30145_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  and (_30146_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor (_30147_, _30146_, _30145_);
  and (_30148_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_30149_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor (_30150_, _30149_, _30148_);
  and (_30151_, _30150_, _30147_);
  and (_30152_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_30153_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nor (_30154_, _30153_, _30152_);
  and (_30155_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_30156_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor (_30157_, _30156_, _30155_);
  and (_30158_, _30157_, _30154_);
  and (_30159_, _30158_, _30151_);
  and (_30160_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  and (_30161_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nor (_30162_, _30161_, _30160_);
  and (_30163_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_30164_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nor (_30165_, _30164_, _30163_);
  and (_30166_, _30165_, _30162_);
  and (_30167_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  and (_30168_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nor (_30169_, _30168_, _30167_);
  and (_30170_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_30171_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nor (_30172_, _30171_, _30170_);
  and (_30173_, _30172_, _30169_);
  and (_30174_, _30173_, _30166_);
  and (_30175_, _30174_, _30159_);
  and (_30176_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_30177_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nor (_30178_, _30177_, _30176_);
  and (_30179_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and (_30180_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor (_30181_, _30180_, _30179_);
  and (_30182_, _30181_, _30178_);
  and (_30183_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_30184_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nor (_30185_, _30184_, _30183_);
  and (_30186_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and (_30187_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nor (_30188_, _30187_, _30186_);
  and (_30189_, _30188_, _30185_);
  and (_30190_, _30189_, _30182_);
  and (_30191_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and (_30192_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nor (_30193_, _30192_, _30191_);
  and (_30194_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_30195_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nor (_30196_, _30195_, _30194_);
  and (_30197_, _30196_, _30193_);
  and (_30198_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and (_30199_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor (_30200_, _30199_, _30198_);
  and (_30201_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_30202_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nor (_30203_, _30202_, _30201_);
  and (_30204_, _30203_, _30200_);
  and (_30205_, _30204_, _30197_);
  and (_30206_, _30205_, _30190_);
  and (_30207_, _30206_, _30175_);
  and (_30208_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_30209_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor (_30210_, _30209_, _30208_);
  and (_30211_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  and (_30212_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor (_30213_, _30212_, _30211_);
  and (_30214_, _30213_, _30210_);
  and (_30215_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_30216_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor (_30217_, _30216_, _30215_);
  and (_30218_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  and (_30219_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nor (_30220_, _30219_, _30218_);
  and (_30221_, _30220_, _30217_);
  and (_30222_, _30221_, _30214_);
  and (_30223_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  and (_30224_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nor (_30225_, _30224_, _30223_);
  and (_30226_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_30227_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nor (_30228_, _30227_, _30226_);
  and (_30229_, _30228_, _30225_);
  and (_30230_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  and (_30231_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nor (_30232_, _30231_, _30230_);
  and (_30233_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_30234_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nor (_30235_, _30234_, _30233_);
  and (_30236_, _30235_, _30232_);
  and (_30237_, _30236_, _30229_);
  and (_30238_, _30237_, _30222_);
  and (_30239_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_30240_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nor (_30241_, _30240_, _30239_);
  and (_30242_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  and (_30243_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nor (_30244_, _30243_, _30242_);
  and (_30245_, _30244_, _30241_);
  and (_30246_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  and (_30247_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nor (_30248_, _30247_, _30246_);
  and (_30249_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_30250_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nor (_30251_, _30250_, _30249_);
  and (_30252_, _30251_, _30248_);
  and (_30253_, _30252_, _30245_);
  and (_30254_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  and (_30255_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nor (_30256_, _30255_, _30254_);
  and (_30257_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  and (_30258_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nor (_30259_, _30258_, _30257_);
  and (_30260_, _30259_, _30256_);
  and (_30261_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  and (_30262_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nor (_30263_, _30262_, _30261_);
  and (_30264_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_30265_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nor (_30266_, _30265_, _30264_);
  and (_30267_, _30266_, _30263_);
  and (_30268_, _30267_, _30260_);
  and (_30269_, _30268_, _30253_);
  and (_30270_, _30269_, _30238_);
  and (_30271_, _30270_, _30207_);
  and (_30272_, _30271_, _30144_);
  and (_30273_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_30274_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor (_30275_, _30274_, _30273_);
  and (_30276_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_30277_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor (_30278_, _30277_, _30276_);
  and (_30279_, _30278_, _30275_);
  and (_30280_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_30281_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor (_30282_, _30281_, _30280_);
  and (_30283_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  and (_30284_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor (_30285_, _30284_, _30283_);
  and (_30286_, _30285_, _30282_);
  and (_30287_, _30286_, _30279_);
  and (_30288_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  and (_30289_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nor (_30290_, _30289_, _30288_);
  and (_30291_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_30292_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nor (_30293_, _30292_, _30291_);
  and (_30294_, _30293_, _30290_);
  and (_30295_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  and (_30296_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nor (_30297_, _30296_, _30295_);
  and (_30298_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_30299_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor (_30300_, _30299_, _30298_);
  and (_30301_, _30300_, _30297_);
  and (_30302_, _30301_, _30294_);
  and (_30303_, _30302_, _30287_);
  and (_30304_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_30305_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nor (_30306_, _30305_, _30304_);
  and (_30307_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  and (_30308_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor (_30309_, _30308_, _30307_);
  and (_30310_, _30309_, _30306_);
  and (_30311_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_30312_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nor (_30313_, _30312_, _30311_);
  and (_30314_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  and (_30315_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nor (_30316_, _30315_, _30314_);
  and (_30317_, _30316_, _30313_);
  and (_30318_, _30317_, _30310_);
  and (_30319_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  and (_30320_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nor (_30321_, _30320_, _30319_);
  and (_30322_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_30323_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor (_30324_, _30323_, _30322_);
  and (_30325_, _30324_, _30321_);
  and (_30326_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  and (_30327_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nor (_30328_, _30327_, _30326_);
  and (_30329_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_30330_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nor (_30331_, _30330_, _30329_);
  and (_30332_, _30331_, _30328_);
  and (_30333_, _30332_, _30325_);
  and (_30334_, _30333_, _30318_);
  and (_30335_, _30334_, _30303_);
  and (_30336_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_30337_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor (_30338_, _30337_, _30336_);
  and (_30339_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  and (_30340_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor (_30341_, _30340_, _30339_);
  and (_30342_, _30341_, _30338_);
  and (_30343_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_30344_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor (_30345_, _30344_, _30343_);
  and (_30346_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_30347_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor (_30348_, _30347_, _30346_);
  and (_30349_, _30348_, _30345_);
  and (_30350_, _30349_, _30342_);
  and (_30351_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  and (_30352_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nor (_30353_, _30352_, _30351_);
  and (_30354_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_30355_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nor (_30356_, _30355_, _30354_);
  and (_30357_, _30356_, _30353_);
  and (_30358_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  and (_30359_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nor (_30360_, _30359_, _30358_);
  and (_30361_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_30362_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor (_30363_, _30362_, _30361_);
  and (_30364_, _30363_, _30360_);
  and (_30365_, _30364_, _30357_);
  and (_30366_, _30365_, _30350_);
  and (_30367_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and (_30368_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nor (_30369_, _30368_, _30367_);
  and (_30370_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  and (_30371_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nor (_30372_, _30371_, _30370_);
  and (_30373_, _30372_, _30369_);
  and (_30374_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and (_30375_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nor (_30376_, _30375_, _30374_);
  and (_30377_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and (_30378_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nor (_30379_, _30378_, _30377_);
  and (_30380_, _30379_, _30376_);
  and (_30381_, _30380_, _30373_);
  and (_30382_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  and (_30383_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nor (_30384_, _30383_, _30382_);
  and (_30385_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and (_30386_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nor (_30387_, _30386_, _30385_);
  and (_30388_, _30387_, _30384_);
  and (_30389_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  and (_30390_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nor (_30391_, _30390_, _30389_);
  and (_30392_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  and (_30393_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  nor (_30394_, _30393_, _30392_);
  and (_30395_, _30394_, _30391_);
  and (_30396_, _30395_, _30388_);
  and (_30397_, _30396_, _30381_);
  and (_30398_, _30397_, _30366_);
  and (_30399_, _30398_, _30335_);
  and (_30400_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  and (_30401_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nor (_30402_, _30401_, _30400_);
  and (_30403_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_30404_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nor (_30405_, _30404_, _30403_);
  and (_30406_, _30405_, _30402_);
  and (_30407_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  and (_30408_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nor (_30409_, _30408_, _30407_);
  and (_30410_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_30411_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor (_30412_, _30411_, _30410_);
  and (_30413_, _30412_, _30409_);
  and (_30414_, _30413_, _30406_);
  and (_30415_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_30416_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor (_30417_, _30416_, _30415_);
  and (_30418_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  and (_30419_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nor (_30420_, _30419_, _30418_);
  and (_30421_, _30420_, _30417_);
  and (_30422_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_30423_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor (_30424_, _30423_, _30422_);
  and (_30425_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  and (_30426_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor (_30427_, _30426_, _30425_);
  and (_30428_, _30427_, _30424_);
  and (_30429_, _30428_, _30421_);
  and (_30430_, _30429_, _30414_);
  and (_30431_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_30432_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nor (_30433_, _30432_, _30431_);
  and (_30434_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  and (_30435_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nor (_30436_, _30435_, _30434_);
  and (_30437_, _30436_, _30433_);
  and (_30438_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  and (_30439_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nor (_30440_, _30439_, _30438_);
  and (_30441_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_30442_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nor (_30443_, _30442_, _30441_);
  and (_30444_, _30443_, _30440_);
  and (_30445_, _30444_, _30437_);
  and (_30446_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  and (_30447_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor (_30448_, _30447_, _30446_);
  and (_30449_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_30450_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nor (_30451_, _30450_, _30449_);
  and (_30452_, _30451_, _30448_);
  and (_30453_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  and (_30454_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor (_30455_, _30454_, _30453_);
  and (_30456_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_30457_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nor (_30458_, _30457_, _30456_);
  and (_30459_, _30458_, _30455_);
  and (_30460_, _30459_, _30452_);
  and (_30461_, _30460_, _30445_);
  and (_30462_, _30461_, _30430_);
  and (_30463_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_30464_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor (_30465_, _30464_, _30463_);
  and (_30466_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  and (_30467_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor (_30468_, _30467_, _30466_);
  and (_30469_, _30468_, _30465_);
  and (_30470_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_30471_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor (_30472_, _30471_, _30470_);
  and (_30473_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  and (_30474_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nor (_30475_, _30474_, _30473_);
  and (_30476_, _30475_, _30472_);
  and (_30477_, _30476_, _30469_);
  and (_30478_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  and (_30479_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nor (_30480_, _30479_, _30478_);
  and (_30481_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_30482_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nor (_30483_, _30482_, _30481_);
  and (_30484_, _30483_, _30480_);
  and (_30485_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  and (_30486_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nor (_30487_, _30486_, _30485_);
  and (_30488_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_30489_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_30490_, _30489_, _30488_);
  and (_30491_, _30490_, _30487_);
  and (_30492_, _30491_, _30484_);
  and (_30493_, _30492_, _30477_);
  and (_30494_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_30495_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_30496_, _30495_, _30494_);
  and (_30497_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_30498_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_30499_, _30498_, _30497_);
  and (_30500_, _30499_, _30496_);
  and (_30501_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_30502_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_30503_, _30502_, _30501_);
  and (_30504_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_30505_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_30506_, _30505_, _30504_);
  and (_30507_, _30506_, _30503_);
  and (_30508_, _30507_, _30500_);
  and (_30509_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_30510_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_30511_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_30512_, _30511_, _30510_);
  nor (_30513_, _30512_, _30509_);
  and (_30514_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_30515_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_30516_, _30515_, _30514_);
  and (_30517_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_30518_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_30519_, _30518_, _30517_);
  and (_30520_, _30519_, _30516_);
  and (_30521_, _30520_, _30513_);
  and (_30522_, _30521_, _30508_);
  and (_30523_, _30522_, _30493_);
  and (_30524_, _30523_, _30462_);
  and (_30525_, _30524_, _30399_);
  and (_30526_, _30525_, _30272_);
  and (_30527_, _30526_, _30017_);
  nor (_30528_, _29491_, iram_op1_reg[3]);
  nor (_30529_, _30528_, _30009_);
  and (_30530_, _30529_, _30527_);
  and (_30531_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  not (_30532_, _30531_);
  and (_30533_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_30534_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_30535_, _30534_, _30533_);
  and (_30536_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  and (_30537_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_30538_, _30537_, _30536_);
  or (_30539_, _30538_, _30535_);
  and (_30540_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  and (_30541_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_30542_, _30541_, _30540_);
  and (_30543_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_30544_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or (_30545_, _30544_, _30543_);
  or (_30546_, _30545_, _30542_);
  or (_30547_, _30546_, _30539_);
  and (_30548_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_30549_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_30550_, _30549_, _30548_);
  and (_30551_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  and (_30552_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_30553_, _30552_, _30551_);
  or (_30554_, _30553_, _30550_);
  and (_30555_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_30556_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_30557_, _30556_, _30555_);
  and (_30558_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_30559_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_30560_, _30559_, _30558_);
  or (_30561_, _30560_, _30557_);
  or (_30562_, _30561_, _30554_);
  or (_30563_, _30562_, _30547_);
  and (_30564_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_30565_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_30566_, _30565_, _30564_);
  and (_30567_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  and (_30568_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or (_30569_, _30568_, _30567_);
  or (_30570_, _30569_, _30566_);
  and (_30571_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_30572_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_30573_, _30572_, _30571_);
  and (_30574_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  and (_30575_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_30576_, _30575_, _30574_);
  or (_30577_, _30576_, _30573_);
  or (_30578_, _30577_, _30570_);
  and (_30579_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  and (_30580_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_30581_, _30580_, _30579_);
  and (_30582_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  and (_30583_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_30584_, _30583_, _30582_);
  or (_30585_, _30584_, _30581_);
  and (_30586_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_30587_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_30588_, _30587_, _30586_);
  and (_30589_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  and (_30590_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_30591_, _30590_, _30589_);
  or (_30592_, _30591_, _30588_);
  or (_30593_, _30592_, _30585_);
  or (_30594_, _30593_, _30578_);
  or (_30595_, _30594_, _30563_);
  and (_30596_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_30597_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or (_30598_, _30597_, _30596_);
  and (_30599_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_30600_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_30601_, _30600_, _30599_);
  or (_30602_, _30601_, _30598_);
  and (_30603_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_30604_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_30605_, _30604_, _30603_);
  and (_30606_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_30607_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nor (_30608_, _30607_, _30606_);
  nand (_30609_, _30608_, _30605_);
  or (_30610_, _30609_, _30602_);
  and (_30611_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  and (_30612_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_30613_, _30612_, _30611_);
  and (_30614_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  and (_30615_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_30616_, _30615_, _30614_);
  or (_30617_, _30616_, _30613_);
  and (_30618_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  and (_30619_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_30620_, _30619_, _30618_);
  and (_30621_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_30622_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_30623_, _30622_, _30621_);
  or (_30624_, _30623_, _30620_);
  or (_30625_, _30624_, _30617_);
  or (_30626_, _30625_, _30610_);
  and (_30627_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  and (_30628_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_30629_, _30628_, _30627_);
  and (_30630_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_30631_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_30632_, _30631_, _30630_);
  or (_30633_, _30632_, _30629_);
  and (_30634_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  and (_30635_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nor (_30636_, _30635_, _30634_);
  and (_30637_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_30638_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nor (_30639_, _30638_, _30637_);
  nand (_30640_, _30639_, _30636_);
  or (_30641_, _30640_, _30633_);
  and (_30642_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_30643_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_30644_, _30643_, _30642_);
  and (_30645_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_30646_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_30647_, _30646_, _30645_);
  or (_30648_, _30647_, _30644_);
  and (_30649_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_30650_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_30651_, _30650_, _30649_);
  and (_30652_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  and (_30653_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_30654_, _30653_, _30652_);
  or (_30655_, _30654_, _30651_);
  or (_30656_, _30655_, _30648_);
  or (_30657_, _30656_, _30641_);
  or (_30658_, _30657_, _30626_);
  or (_30659_, _30658_, _30595_);
  and (_30660_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_30661_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  or (_30662_, _30661_, _30660_);
  and (_30663_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_30664_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_30665_, _30664_, _30663_);
  or (_30666_, _30665_, _30662_);
  and (_30667_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  and (_30668_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_30669_, _30668_, _30667_);
  and (_30670_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_30671_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_30672_, _30671_, _30670_);
  or (_30673_, _30672_, _30669_);
  or (_30674_, _30673_, _30666_);
  and (_30675_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_30676_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_30677_, _30676_, _30675_);
  and (_30678_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_30679_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or (_30680_, _30679_, _30678_);
  or (_30681_, _30680_, _30677_);
  and (_30682_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_30683_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor (_30684_, _30683_, _30682_);
  and (_30685_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and (_30686_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor (_30687_, _30686_, _30685_);
  nand (_30688_, _30687_, _30684_);
  or (_30689_, _30688_, _30681_);
  or (_30690_, _30689_, _30674_);
  and (_30691_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_30692_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_30693_, _30692_, _30691_);
  and (_30694_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_30695_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_30696_, _30695_, _30694_);
  or (_30697_, _30696_, _30693_);
  and (_30698_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  and (_30699_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor (_30700_, _30699_, _30698_);
  and (_30701_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_30702_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor (_30703_, _30702_, _30701_);
  nand (_30704_, _30703_, _30700_);
  or (_30705_, _30704_, _30697_);
  and (_30706_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_30707_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_30708_, _30707_, _30706_);
  and (_30709_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  and (_30710_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_30711_, _30710_, _30709_);
  or (_30712_, _30711_, _30708_);
  and (_30713_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  and (_30714_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_30715_, _30714_, _30713_);
  and (_30716_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  and (_30717_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_30718_, _30717_, _30716_);
  or (_30719_, _30718_, _30715_);
  or (_30720_, _30719_, _30712_);
  or (_30721_, _30720_, _30705_);
  or (_30722_, _30721_, _30690_);
  and (_30723_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_30724_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_30725_, _30724_, _30723_);
  and (_30726_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  and (_30727_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nor (_30728_, _30727_, _30726_);
  nand (_30729_, _30728_, _30725_);
  and (_30730_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_30731_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nor (_30732_, _30731_, _30730_);
  and (_30733_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  and (_30734_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nor (_30735_, _30734_, _30733_);
  nand (_30736_, _30735_, _30732_);
  or (_30737_, _30736_, _30729_);
  and (_30738_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  and (_30739_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_30740_, _30739_, _30738_);
  and (_30741_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  and (_30742_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_30743_, _30742_, _30741_);
  or (_30744_, _30743_, _30740_);
  and (_30745_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  and (_30746_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_30747_, _30746_, _30745_);
  and (_30748_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_30749_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_30750_, _30749_, _30748_);
  or (_30751_, _30750_, _30747_);
  or (_30752_, _30751_, _30744_);
  or (_30753_, _30752_, _30737_);
  and (_30754_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_30755_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_30756_, _30755_, _30754_);
  and (_30757_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_30758_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_30759_, _30758_, _30757_);
  or (_30760_, _30759_, _30756_);
  and (_30761_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_30762_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_30763_, _30762_, _30761_);
  and (_30764_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_30765_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_30766_, _30765_, _30764_);
  or (_30767_, _30766_, _30763_);
  or (_30768_, _30767_, _30760_);
  and (_30769_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  and (_30770_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  or (_30771_, _30770_, _30769_);
  and (_30772_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_30773_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_30774_, _30773_, _30772_);
  or (_30775_, _30774_, _30771_);
  and (_30776_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_30777_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_30778_, _30777_, _30776_);
  and (_30779_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  and (_30780_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_30781_, _30780_, _30779_);
  or (_30782_, _30781_, _30778_);
  or (_30783_, _30782_, _30775_);
  or (_30784_, _30783_, _30768_);
  or (_30785_, _30784_, _30753_);
  or (_30786_, _30785_, _30722_);
  or (_30787_, _30786_, _30659_);
  and (_30788_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_30789_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_30790_, _30789_, _30788_);
  and (_30791_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  and (_30792_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_30793_, _30792_, _30791_);
  or (_30794_, _30793_, _30790_);
  and (_30795_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  and (_30796_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_30797_, _30796_, _30795_);
  and (_30798_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_30799_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_30800_, _30799_, _30798_);
  or (_30801_, _30800_, _30797_);
  or (_30802_, _30801_, _30794_);
  and (_30803_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  and (_30804_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or (_30805_, _30804_, _30803_);
  and (_30806_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_30807_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or (_30808_, _30807_, _30806_);
  or (_30809_, _30808_, _30805_);
  and (_30810_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_30811_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  or (_30812_, _30811_, _30810_);
  and (_30813_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  and (_30814_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_30815_, _30814_, _30813_);
  or (_30816_, _30815_, _30812_);
  or (_30817_, _30816_, _30809_);
  or (_30818_, _30817_, _30802_);
  and (_30819_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  and (_30820_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or (_30821_, _30820_, _30819_);
  and (_30822_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_30823_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_30824_, _30823_, _30822_);
  or (_30825_, _30824_, _30821_);
  and (_30826_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  and (_30827_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or (_30828_, _30827_, _30826_);
  and (_30829_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  and (_30830_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_30831_, _30830_, _30829_);
  or (_30832_, _30831_, _30828_);
  or (_30833_, _30832_, _30825_);
  and (_30834_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_30835_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_30836_, _30835_, _30834_);
  and (_30837_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_30838_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_30839_, _30838_, _30837_);
  or (_30840_, _30839_, _30836_);
  and (_30841_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  and (_30842_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor (_30843_, _30842_, _30841_);
  and (_30844_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_30845_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_30846_, _30845_, _30844_);
  nand (_30847_, _30846_, _30843_);
  or (_30848_, _30847_, _30840_);
  or (_30849_, _30848_, _30833_);
  or (_30850_, _30849_, _30818_);
  and (_30851_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_30852_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor (_30853_, _30852_, _30851_);
  and (_30854_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  and (_30855_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nor (_30856_, _30855_, _30854_);
  nand (_30857_, _30856_, _30853_);
  and (_30858_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and (_30859_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  or (_30860_, _30859_, _30858_);
  and (_30861_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_30862_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or (_30863_, _30862_, _30861_);
  or (_30864_, _30863_, _30860_);
  or (_30865_, _30864_, _30857_);
  and (_30866_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  and (_30867_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  and (_30868_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_30869_, _30868_, _30867_);
  or (_30870_, _30869_, _30866_);
  and (_30871_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_30872_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor (_30873_, _30872_, _30871_);
  and (_30874_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  and (_30875_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nor (_30876_, _30875_, _30874_);
  nand (_30877_, _30876_, _30873_);
  or (_30878_, _30877_, _30870_);
  or (_30879_, _30878_, _30865_);
  and (_30880_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_30881_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_30882_, _30881_, _30880_);
  and (_30883_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  and (_30884_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_30885_, _30884_, _30883_);
  or (_30886_, _30885_, _30882_);
  and (_30887_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  and (_30888_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_30889_, _30888_, _30887_);
  and (_30890_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_30891_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  or (_30892_, _30891_, _30890_);
  or (_30893_, _30892_, _30889_);
  or (_30894_, _30893_, _30886_);
  and (_30895_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  and (_30896_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_30897_, _30896_, _30895_);
  and (_30898_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and (_30899_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_30900_, _30899_, _30898_);
  or (_30901_, _30900_, _30897_);
  and (_30902_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_30903_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_30904_, _30903_, _30902_);
  and (_30905_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_30906_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_30907_, _30906_, _30905_);
  or (_30908_, _30907_, _30904_);
  or (_30909_, _30908_, _30901_);
  or (_30910_, _30909_, _30894_);
  or (_30911_, _30910_, _30879_);
  or (_30912_, _30911_, _30850_);
  and (_30913_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  and (_30914_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_30915_, _30914_, _30913_);
  and (_30916_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_30917_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_30918_, _30917_, _30916_);
  or (_30919_, _30918_, _30915_);
  and (_30920_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_30921_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_30922_, _30921_, _30920_);
  and (_30923_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  and (_30924_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or (_30925_, _30924_, _30923_);
  or (_30926_, _30925_, _30922_);
  or (_30927_, _30926_, _30919_);
  and (_30928_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_30929_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_30930_, _30929_, _30928_);
  and (_30931_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  and (_30932_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_30933_, _30932_, _30931_);
  or (_30934_, _30933_, _30930_);
  and (_30935_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_30936_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_30937_, _30936_, _30935_);
  and (_30938_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_30939_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_30940_, _30939_, _30938_);
  or (_30941_, _30940_, _30937_);
  or (_30942_, _30941_, _30934_);
  or (_30943_, _30942_, _30927_);
  and (_30944_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_30945_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_30946_, _30945_, _30944_);
  and (_30947_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  and (_30948_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_30949_, _30948_, _30947_);
  or (_30950_, _30949_, _30946_);
  and (_30951_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_30952_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_30953_, _30952_, _30951_);
  and (_30954_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_30955_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_30956_, _30955_, _30954_);
  or (_30957_, _30956_, _30953_);
  or (_30958_, _30957_, _30950_);
  and (_30959_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  and (_30960_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_30961_, _30960_, _30959_);
  and (_30962_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and (_30963_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_30964_, _30963_, _30962_);
  or (_30965_, _30964_, _30961_);
  and (_30966_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  and (_30967_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_30968_, _30967_, _30966_);
  and (_30969_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_30970_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_30971_, _30970_, _30969_);
  or (_30972_, _30971_, _30968_);
  or (_30973_, _30972_, _30965_);
  or (_30974_, _30973_, _30958_);
  or (_30975_, _30974_, _30943_);
  and (_30976_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_30977_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_30978_, _30977_, _30976_);
  and (_30979_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  and (_30980_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_30981_, _30980_, _30979_);
  or (_30982_, _30981_, _30978_);
  and (_30983_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_30984_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_30985_, _30984_, _30983_);
  and (_30986_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and (_30987_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_30988_, _30987_, _30986_);
  or (_30989_, _30988_, _30985_);
  or (_30990_, _30989_, _30982_);
  and (_30991_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_30992_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  or (_30993_, _30992_, _30991_);
  and (_30994_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_30995_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_30996_, _30995_, _30994_);
  or (_30997_, _30996_, _30993_);
  and (_30998_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  and (_30999_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_31000_, _30999_, _30998_);
  and (_31001_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_31002_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_31003_, _31002_, _31001_);
  or (_31004_, _31003_, _31000_);
  or (_31005_, _31004_, _30997_);
  or (_31006_, _31005_, _30990_);
  and (_31007_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_31008_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_31009_, _31008_, _31007_);
  and (_31010_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  and (_31011_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_31012_, _31011_, _31010_);
  or (_31013_, _31012_, _31009_);
  and (_31014_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  and (_31015_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nor (_31016_, _31015_, _31014_);
  and (_31017_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_31018_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nor (_31019_, _31018_, _31017_);
  nand (_31020_, _31019_, _31016_);
  or (_31021_, _31020_, _31013_);
  and (_31022_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_31023_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or (_31024_, _31023_, _31022_);
  and (_31025_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_31026_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_31027_, _31026_, _31025_);
  or (_31028_, _31027_, _31024_);
  and (_31029_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_31030_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_31031_, _31030_, _31029_);
  and (_31032_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_31033_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_31034_, _31033_, _31032_);
  or (_31035_, _31034_, _31031_);
  or (_31036_, _31035_, _31028_);
  or (_31037_, _31036_, _31021_);
  or (_31038_, _31037_, _31006_);
  or (_31039_, _31038_, _30975_);
  or (_31040_, _31039_, _30912_);
  nor (_31041_, _31040_, _30787_);
  and (_31042_, _31041_, _30532_);
  and (_31043_, _30010_, iram_op1_reg[5]);
  and (_31044_, _31043_, iram_op1_reg[6]);
  nor (_31045_, _31044_, iram_op1_reg[7]);
  and (_31046_, _31044_, iram_op1_reg[7]);
  nor (_31047_, _31046_, _31045_);
  nor (_31048_, _31047_, _31042_);
  or (_31049_, _31048_, _30530_);
  or (_31050_, _31049_, _30015_);
  or (_31051_, _31050_, _29496_);
  and (_31052_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  not (_31053_, _31052_);
  and (_31054_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  and (_31055_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nor (_31056_, _31055_, _31054_);
  and (_31057_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_31058_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nor (_31059_, _31058_, _31057_);
  and (_31060_, _31059_, _31056_);
  and (_31061_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  and (_31062_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nor (_31063_, _31062_, _31061_);
  and (_31064_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_31065_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nor (_31066_, _31065_, _31064_);
  and (_31067_, _31066_, _31063_);
  and (_31068_, _31067_, _31060_);
  and (_31069_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_31070_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor (_31071_, _31070_, _31069_);
  and (_31072_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  and (_31073_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor (_31074_, _31073_, _31072_);
  and (_31075_, _31074_, _31071_);
  and (_31076_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_31077_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor (_31078_, _31077_, _31076_);
  and (_31079_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  and (_31080_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nor (_31081_, _31080_, _31079_);
  and (_31082_, _31081_, _31078_);
  and (_31083_, _31082_, _31075_);
  and (_31084_, _31083_, _31068_);
  and (_31085_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  and (_31086_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nor (_31087_, _31086_, _31085_);
  and (_31088_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_31089_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nor (_31090_, _31089_, _31088_);
  and (_31091_, _31090_, _31087_);
  and (_31092_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  and (_31093_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nor (_31094_, _31093_, _31092_);
  and (_31095_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_31096_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nor (_31097_, _31096_, _31095_);
  and (_31098_, _31097_, _31094_);
  and (_31099_, _31098_, _31091_);
  and (_31100_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_31101_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nor (_31102_, _31101_, _31100_);
  and (_31103_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  and (_31104_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nor (_31105_, _31104_, _31103_);
  and (_31106_, _31105_, _31102_);
  and (_31107_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_31108_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nor (_31109_, _31108_, _31107_);
  and (_31110_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and (_31111_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nor (_31112_, _31111_, _31110_);
  and (_31113_, _31112_, _31109_);
  and (_31114_, _31113_, _31106_);
  and (_31115_, _31114_, _31099_);
  and (_31116_, _31115_, _31084_);
  and (_31117_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_31118_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor (_31119_, _31118_, _31117_);
  and (_31120_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and (_31121_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor (_31122_, _31121_, _31120_);
  and (_31123_, _31122_, _31119_);
  and (_31124_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_31125_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor (_31126_, _31125_, _31124_);
  and (_31127_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and (_31128_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nor (_31129_, _31128_, _31127_);
  and (_31130_, _31129_, _31126_);
  and (_31131_, _31130_, _31123_);
  and (_31132_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and (_31133_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nor (_31134_, _31133_, _31132_);
  and (_31135_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_31136_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nor (_31137_, _31136_, _31135_);
  and (_31138_, _31137_, _31134_);
  and (_31139_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and (_31140_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nor (_31141_, _31140_, _31139_);
  and (_31142_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_31143_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nor (_31144_, _31143_, _31142_);
  and (_31145_, _31144_, _31141_);
  and (_31146_, _31145_, _31138_);
  and (_31147_, _31146_, _31131_);
  and (_31148_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_31149_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor (_31150_, _31149_, _31148_);
  and (_31151_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  and (_31152_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nor (_31153_, _31152_, _31151_);
  and (_31154_, _31153_, _31150_);
  and (_31155_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  and (_31156_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor (_31157_, _31156_, _31155_);
  and (_31158_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  and (_31159_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nor (_31160_, _31159_, _31158_);
  and (_31161_, _31160_, _31157_);
  and (_31162_, _31161_, _31154_);
  and (_31163_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_31164_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nor (_31165_, _31164_, _31163_);
  and (_31166_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  and (_31167_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor (_31168_, _31167_, _31166_);
  and (_31169_, _31168_, _31165_);
  and (_31170_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_31171_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nor (_31172_, _31171_, _31170_);
  and (_31173_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  and (_31174_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nor (_31175_, _31174_, _31173_);
  and (_31176_, _31175_, _31172_);
  and (_31177_, _31176_, _31169_);
  and (_31178_, _31177_, _31162_);
  and (_31179_, _31178_, _31147_);
  and (_31180_, _31179_, _31116_);
  and (_31181_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_31182_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nor (_31183_, _31182_, _31181_);
  and (_31184_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  and (_31185_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor (_31186_, _31185_, _31184_);
  and (_31187_, _31186_, _31183_);
  and (_31188_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_31189_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor (_31190_, _31189_, _31188_);
  and (_31191_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  and (_31192_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nor (_31193_, _31192_, _31191_);
  and (_31194_, _31193_, _31190_);
  and (_31195_, _31194_, _31187_);
  and (_31196_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  and (_31197_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nor (_31198_, _31197_, _31196_);
  and (_31199_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_31200_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor (_31201_, _31200_, _31199_);
  and (_31202_, _31201_, _31198_);
  and (_31203_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  and (_31204_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nor (_31205_, _31204_, _31203_);
  and (_31206_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_31207_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nor (_31208_, _31207_, _31206_);
  and (_31209_, _31208_, _31205_);
  and (_31210_, _31209_, _31202_);
  and (_31211_, _31210_, _31195_);
  and (_31212_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and (_31213_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor (_31214_, _31213_, _31212_);
  and (_31215_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_31216_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nor (_31217_, _31216_, _31215_);
  and (_31218_, _31217_, _31214_);
  and (_31219_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_31220_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nor (_31221_, _31220_, _31219_);
  and (_31222_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_31223_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nor (_31224_, _31223_, _31222_);
  and (_31225_, _31224_, _31221_);
  and (_31226_, _31225_, _31218_);
  and (_31227_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_31228_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nor (_31229_, _31228_, _31227_);
  and (_31230_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_31231_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nor (_31232_, _31231_, _31230_);
  and (_31233_, _31232_, _31229_);
  and (_31234_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_31235_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nor (_31236_, _31235_, _31234_);
  and (_31237_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  and (_31238_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nor (_31239_, _31238_, _31237_);
  and (_31240_, _31239_, _31236_);
  and (_31241_, _31240_, _31233_);
  and (_31242_, _31241_, _31226_);
  and (_31243_, _31242_, _31211_);
  and (_31244_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_31245_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor (_31246_, _31245_, _31244_);
  and (_31247_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  and (_31248_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nor (_31249_, _31248_, _31247_);
  and (_31250_, _31249_, _31246_);
  and (_31251_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  and (_31252_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nor (_31253_, _31252_, _31251_);
  and (_31254_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_31255_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nor (_31256_, _31255_, _31254_);
  and (_31257_, _31256_, _31253_);
  and (_31258_, _31257_, _31250_);
  and (_31259_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_31260_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor (_31261_, _31260_, _31259_);
  and (_31262_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  and (_31263_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor (_31264_, _31263_, _31262_);
  and (_31265_, _31264_, _31261_);
  and (_31266_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_31267_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor (_31268_, _31267_, _31266_);
  and (_31269_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  and (_31270_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nor (_31271_, _31270_, _31269_);
  and (_31272_, _31271_, _31268_);
  and (_31273_, _31272_, _31265_);
  and (_31274_, _31273_, _31258_);
  and (_31275_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_31276_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nor (_31277_, _31276_, _31275_);
  and (_31278_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  and (_31279_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor (_31280_, _31279_, _31278_);
  and (_31281_, _31280_, _31277_);
  and (_31282_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_31283_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nor (_31284_, _31283_, _31282_);
  and (_31285_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  and (_31286_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nor (_31287_, _31286_, _31285_);
  and (_31288_, _31287_, _31284_);
  and (_31289_, _31288_, _31281_);
  and (_31290_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  and (_31291_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nor (_31292_, _31291_, _31290_);
  and (_31293_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_31294_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor (_31295_, _31294_, _31293_);
  and (_31296_, _31295_, _31292_);
  and (_31297_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  and (_31298_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nor (_31299_, _31298_, _31297_);
  and (_31300_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  and (_31301_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nor (_31302_, _31301_, _31300_);
  and (_31303_, _31302_, _31299_);
  and (_31304_, _31303_, _31296_);
  and (_31305_, _31304_, _31289_);
  and (_31306_, _31305_, _31274_);
  and (_31307_, _31306_, _31243_);
  and (_31308_, _31307_, _31180_);
  and (_31309_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_31310_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor (_31311_, _31310_, _31309_);
  and (_31312_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  and (_31313_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor (_31314_, _31313_, _31312_);
  and (_31315_, _31314_, _31311_);
  and (_31316_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_31317_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor (_31318_, _31317_, _31316_);
  and (_31319_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  and (_31320_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nor (_31321_, _31320_, _31319_);
  and (_31322_, _31321_, _31318_);
  and (_31323_, _31322_, _31315_);
  and (_31324_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  and (_31325_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nor (_31326_, _31325_, _31324_);
  and (_31327_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_31328_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor (_31329_, _31328_, _31327_);
  and (_31330_, _31329_, _31326_);
  and (_31331_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  and (_31332_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nor (_31333_, _31332_, _31331_);
  and (_31334_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_31335_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nor (_31336_, _31335_, _31334_);
  and (_31337_, _31336_, _31333_);
  and (_31338_, _31337_, _31330_);
  and (_31339_, _31338_, _31323_);
  and (_31340_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  and (_31341_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nor (_31342_, _31341_, _31340_);
  and (_31343_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_31344_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nor (_31345_, _31344_, _31343_);
  and (_31346_, _31345_, _31342_);
  and (_31347_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  and (_31348_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor (_31349_, _31348_, _31347_);
  and (_31350_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  and (_31351_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nor (_31352_, _31351_, _31350_);
  and (_31353_, _31352_, _31349_);
  and (_31354_, _31353_, _31346_);
  and (_31355_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_31356_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nor (_31357_, _31356_, _31355_);
  and (_31358_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  and (_31359_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nor (_31360_, _31359_, _31358_);
  and (_31361_, _31360_, _31357_);
  and (_31362_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_31363_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nor (_31364_, _31363_, _31362_);
  and (_31365_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  and (_31366_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nor (_31367_, _31366_, _31365_);
  and (_31368_, _31367_, _31364_);
  and (_31369_, _31368_, _31361_);
  and (_31370_, _31369_, _31354_);
  and (_31371_, _31370_, _31339_);
  and (_31372_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_31373_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor (_31374_, _31373_, _31372_);
  and (_31375_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  and (_31376_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nor (_31377_, _31376_, _31375_);
  and (_31378_, _31377_, _31374_);
  and (_31379_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  and (_31380_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nor (_31381_, _31380_, _31379_);
  and (_31382_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_31383_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nor (_31384_, _31383_, _31382_);
  and (_31385_, _31384_, _31381_);
  and (_31386_, _31385_, _31378_);
  and (_31387_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_31388_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor (_31389_, _31388_, _31387_);
  and (_31390_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  and (_31391_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor (_31392_, _31391_, _31390_);
  and (_31393_, _31392_, _31389_);
  and (_31394_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_31395_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor (_31396_, _31395_, _31394_);
  and (_31397_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  and (_31398_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nor (_31399_, _31398_, _31397_);
  and (_31400_, _31399_, _31396_);
  and (_31401_, _31400_, _31393_);
  and (_31402_, _31401_, _31386_);
  and (_31403_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_31404_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nor (_31405_, _31404_, _31403_);
  and (_31406_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  and (_31407_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nor (_31408_, _31407_, _31406_);
  and (_31409_, _31408_, _31405_);
  and (_31410_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and (_31411_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nor (_31412_, _31411_, _31410_);
  and (_31413_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  and (_31414_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nor (_31415_, _31414_, _31413_);
  and (_31416_, _31415_, _31412_);
  and (_31417_, _31416_, _31409_);
  and (_31418_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  and (_31419_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nor (_31420_, _31419_, _31418_);
  and (_31421_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_31422_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor (_31423_, _31422_, _31421_);
  and (_31424_, _31423_, _31420_);
  and (_31425_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  and (_31426_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor (_31427_, _31426_, _31425_);
  and (_31428_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  and (_31429_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor (_31430_, _31429_, _31428_);
  and (_31431_, _31430_, _31427_);
  and (_31432_, _31431_, _31424_);
  and (_31433_, _31432_, _31417_);
  and (_31434_, _31433_, _31402_);
  and (_31435_, _31434_, _31371_);
  and (_31436_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_31437_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor (_31438_, _31437_, _31436_);
  and (_31439_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  and (_31440_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nor (_31441_, _31440_, _31439_);
  and (_31442_, _31441_, _31438_);
  and (_31443_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_31444_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor (_31445_, _31444_, _31443_);
  and (_31446_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  and (_31447_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor (_31448_, _31447_, _31446_);
  and (_31449_, _31448_, _31445_);
  and (_31450_, _31449_, _31442_);
  and (_31451_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  and (_31452_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nor (_31453_, _31452_, _31451_);
  and (_31454_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_31455_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nor (_31456_, _31455_, _31454_);
  and (_31457_, _31456_, _31453_);
  and (_31458_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  and (_31459_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nor (_31460_, _31459_, _31458_);
  and (_31461_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_31462_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor (_31463_, _31462_, _31461_);
  and (_31464_, _31463_, _31460_);
  and (_31465_, _31464_, _31457_);
  and (_31466_, _31465_, _31450_);
  and (_31467_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  and (_31468_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nor (_31469_, _31468_, _31467_);
  and (_31470_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_31471_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nor (_31472_, _31471_, _31470_);
  and (_31473_, _31472_, _31469_);
  and (_31474_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  and (_31475_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nor (_31476_, _31475_, _31474_);
  and (_31477_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_31478_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor (_31479_, _31478_, _31477_);
  and (_31480_, _31479_, _31476_);
  and (_31481_, _31480_, _31473_);
  and (_31482_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_31483_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nor (_31484_, _31483_, _31482_);
  and (_31485_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  and (_31486_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nor (_31487_, _31486_, _31485_);
  and (_31488_, _31487_, _31484_);
  and (_31489_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_31490_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nor (_31491_, _31490_, _31489_);
  and (_31492_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  and (_31493_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor (_31494_, _31493_, _31492_);
  and (_31495_, _31494_, _31491_);
  and (_31496_, _31495_, _31488_);
  and (_31497_, _31496_, _31481_);
  and (_31498_, _31497_, _31466_);
  and (_31499_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  and (_31500_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor (_31501_, _31500_, _31499_);
  and (_31502_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_31503_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor (_31504_, _31503_, _31502_);
  and (_31505_, _31504_, _31501_);
  and (_31506_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_31507_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nor (_31508_, _31507_, _31506_);
  and (_31509_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_31510_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor (_31511_, _31510_, _31509_);
  and (_31512_, _31511_, _31508_);
  and (_31513_, _31512_, _31505_);
  and (_31514_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  and (_31515_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nor (_31516_, _31515_, _31514_);
  and (_31517_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_31518_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nor (_31519_, _31518_, _31517_);
  and (_31520_, _31519_, _31516_);
  and (_31521_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  and (_31522_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nor (_31523_, _31522_, _31521_);
  and (_31524_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_31525_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nor (_31526_, _31525_, _31524_);
  and (_31527_, _31526_, _31523_);
  and (_31528_, _31527_, _31520_);
  and (_31529_, _31528_, _31513_);
  and (_31530_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_31531_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_31532_, _31531_, _31530_);
  and (_31533_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_31534_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_31535_, _31534_, _31533_);
  and (_31536_, _31535_, _31532_);
  and (_31537_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_31538_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_31539_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_31540_, _31539_, _31538_);
  nor (_31541_, _31540_, _31537_);
  and (_31542_, _31541_, _31536_);
  and (_31543_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_31544_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_31545_, _31544_, _31543_);
  and (_31546_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_31547_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_31548_, _31547_, _31546_);
  and (_31549_, _31548_, _31545_);
  and (_31550_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_31551_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_31552_, _31551_, _31550_);
  and (_31553_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_31554_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_31555_, _31554_, _31553_);
  and (_31556_, _31555_, _31552_);
  and (_31557_, _31556_, _31549_);
  and (_31558_, _31557_, _31542_);
  and (_31559_, _31558_, _31529_);
  and (_31560_, _31559_, _31498_);
  and (_31561_, _31560_, _31435_);
  and (_31562_, _31561_, _31308_);
  and (_31563_, _31562_, _31053_);
  nor (_31564_, _31563_, _21566_);
  and (_31565_, _31563_, _21566_);
  or (_31566_, _31565_, _31564_);
  and (_31567_, _31566_, iram_op1_reg[0]);
  and (_31568_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  not (_31569_, _31568_);
  and (_31570_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  and (_31571_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor (_31572_, _31571_, _31570_);
  and (_31573_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_31574_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor (_31575_, _31574_, _31573_);
  and (_31576_, _31575_, _31572_);
  and (_31577_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_31578_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor (_31579_, _31578_, _31577_);
  and (_31580_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_31581_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor (_31582_, _31581_, _31580_);
  and (_31583_, _31582_, _31579_);
  and (_31584_, _31583_, _31576_);
  and (_31585_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_31586_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nor (_31587_, _31586_, _31585_);
  and (_31588_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  and (_31589_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nor (_31590_, _31589_, _31588_);
  and (_31591_, _31590_, _31587_);
  and (_31592_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  and (_31593_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nor (_31594_, _31593_, _31592_);
  and (_31595_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_31596_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nor (_31597_, _31596_, _31595_);
  and (_31598_, _31597_, _31594_);
  and (_31599_, _31598_, _31591_);
  and (_31600_, _31599_, _31584_);
  and (_31601_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  and (_31602_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nor (_31603_, _31602_, _31601_);
  and (_31604_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_31605_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nor (_31606_, _31605_, _31604_);
  and (_31607_, _31606_, _31603_);
  and (_31608_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_31609_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nor (_31610_, _31609_, _31608_);
  and (_31611_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and (_31612_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nor (_31613_, _31612_, _31611_);
  and (_31614_, _31613_, _31610_);
  and (_31615_, _31614_, _31607_);
  and (_31616_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  and (_31617_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor (_31618_, _31617_, _31616_);
  and (_31619_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  and (_31620_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nor (_31621_, _31620_, _31619_);
  and (_31622_, _31621_, _31618_);
  and (_31623_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  and (_31624_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor (_31625_, _31624_, _31623_);
  and (_31626_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_31627_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor (_31628_, _31627_, _31626_);
  and (_31629_, _31628_, _31625_);
  and (_31630_, _31629_, _31622_);
  and (_31631_, _31630_, _31615_);
  and (_31632_, _31631_, _31600_);
  and (_31633_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_31634_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  nor (_31635_, _31634_, _31633_);
  and (_31636_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and (_31637_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  nor (_31638_, _31637_, _31636_);
  and (_31639_, _31638_, _31635_);
  and (_31640_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_31641_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  nor (_31642_, _31641_, _31640_);
  and (_31643_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and (_31644_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  nor (_31645_, _31644_, _31643_);
  and (_31646_, _31645_, _31642_);
  and (_31647_, _31646_, _31639_);
  and (_31648_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and (_31649_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  nor (_31650_, _31649_, _31648_);
  and (_31651_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_31652_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  nor (_31653_, _31652_, _31651_);
  and (_31654_, _31653_, _31650_);
  and (_31655_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and (_31656_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  nor (_31657_, _31656_, _31655_);
  and (_31658_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_31659_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor (_31660_, _31659_, _31658_);
  and (_31661_, _31660_, _31657_);
  and (_31662_, _31661_, _31654_);
  and (_31663_, _31662_, _31647_);
  and (_31664_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_31665_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nor (_31666_, _31665_, _31664_);
  and (_31667_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  and (_31668_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nor (_31669_, _31668_, _31667_);
  and (_31670_, _31669_, _31666_);
  and (_31671_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_31672_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nor (_31673_, _31672_, _31671_);
  and (_31674_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  and (_31675_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nor (_31676_, _31675_, _31674_);
  and (_31677_, _31676_, _31673_);
  and (_31678_, _31677_, _31670_);
  and (_31679_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  and (_31680_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nor (_31681_, _31680_, _31679_);
  and (_31682_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_31683_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nor (_31684_, _31683_, _31682_);
  and (_31685_, _31684_, _31681_);
  and (_31686_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  and (_31687_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nor (_31688_, _31687_, _31686_);
  and (_31689_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_31690_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nor (_31691_, _31690_, _31689_);
  and (_31692_, _31691_, _31688_);
  and (_31693_, _31692_, _31685_);
  and (_31694_, _31693_, _31678_);
  and (_31695_, _31694_, _31663_);
  and (_31696_, _31695_, _31632_);
  and (_31697_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  and (_31698_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nor (_31699_, _31698_, _31697_);
  and (_31700_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_31701_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nor (_31702_, _31701_, _31700_);
  and (_31703_, _31702_, _31699_);
  and (_31704_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_31705_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nor (_31706_, _31705_, _31704_);
  and (_31707_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  and (_31708_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nor (_31709_, _31708_, _31707_);
  and (_31710_, _31709_, _31706_);
  and (_31711_, _31710_, _31703_);
  and (_31712_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_31713_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor (_31714_, _31713_, _31712_);
  and (_31715_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  and (_31716_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor (_31717_, _31716_, _31715_);
  and (_31718_, _31717_, _31714_);
  and (_31719_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_31720_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor (_31721_, _31720_, _31719_);
  and (_31722_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_31723_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor (_31724_, _31723_, _31722_);
  and (_31725_, _31724_, _31721_);
  and (_31726_, _31725_, _31718_);
  and (_31727_, _31726_, _31711_);
  and (_31728_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_31729_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  nor (_31730_, _31729_, _31728_);
  and (_31731_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  and (_31732_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  nor (_31733_, _31732_, _31731_);
  and (_31734_, _31733_, _31730_);
  and (_31735_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_31736_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  nor (_31737_, _31736_, _31735_);
  and (_31738_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_31739_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  nor (_31740_, _31739_, _31738_);
  and (_31741_, _31740_, _31737_);
  and (_31742_, _31741_, _31734_);
  and (_31743_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_31744_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  nor (_31745_, _31744_, _31743_);
  and (_31746_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_31747_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  nor (_31748_, _31747_, _31746_);
  and (_31749_, _31748_, _31745_);
  and (_31750_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_31751_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  nor (_31752_, _31751_, _31750_);
  and (_31753_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_31754_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  nor (_31755_, _31754_, _31753_);
  and (_31756_, _31755_, _31752_);
  and (_31757_, _31756_, _31749_);
  and (_31758_, _31757_, _31742_);
  and (_31759_, _31758_, _31727_);
  and (_31760_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_31761_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor (_31762_, _31761_, _31760_);
  and (_31763_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  and (_31764_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor (_31765_, _31764_, _31763_);
  and (_31766_, _31765_, _31762_);
  and (_31767_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_31768_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor (_31769_, _31768_, _31767_);
  and (_31770_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  and (_31771_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nor (_31772_, _31771_, _31770_);
  and (_31773_, _31772_, _31769_);
  and (_31774_, _31773_, _31766_);
  and (_31775_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  and (_31776_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nor (_31777_, _31776_, _31775_);
  and (_31778_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_31779_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nor (_31780_, _31779_, _31778_);
  and (_31781_, _31780_, _31777_);
  and (_31782_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  and (_31783_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nor (_31784_, _31783_, _31782_);
  and (_31785_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_31786_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor (_31787_, _31786_, _31785_);
  and (_31788_, _31787_, _31784_);
  and (_31789_, _31788_, _31781_);
  and (_31790_, _31789_, _31774_);
  and (_31791_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  and (_31792_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nor (_31793_, _31792_, _31791_);
  and (_31794_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_31795_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nor (_31796_, _31795_, _31794_);
  and (_31797_, _31796_, _31793_);
  and (_31798_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  and (_31799_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nor (_31800_, _31799_, _31798_);
  and (_31801_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  and (_31802_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nor (_31803_, _31802_, _31801_);
  and (_31804_, _31803_, _31800_);
  and (_31805_, _31804_, _31797_);
  and (_31806_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_31807_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nor (_31808_, _31807_, _31806_);
  and (_31809_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  and (_31810_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nor (_31811_, _31810_, _31809_);
  and (_31812_, _31811_, _31808_);
  and (_31813_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  and (_31814_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nor (_31815_, _31814_, _31813_);
  and (_31816_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_31817_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nor (_31818_, _31817_, _31816_);
  and (_31819_, _31818_, _31815_);
  and (_31820_, _31819_, _31812_);
  and (_31821_, _31820_, _31805_);
  and (_31822_, _31821_, _31790_);
  and (_31823_, _31822_, _31759_);
  and (_31824_, _31823_, _31696_);
  and (_31825_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_31826_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor (_31827_, _31826_, _31825_);
  and (_31828_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_31829_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor (_31830_, _31829_, _31828_);
  and (_31831_, _31830_, _31827_);
  and (_31832_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_31833_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor (_31834_, _31833_, _31832_);
  and (_31835_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  and (_31836_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor (_31837_, _31836_, _31835_);
  and (_31838_, _31837_, _31834_);
  and (_31839_, _31838_, _31831_);
  and (_31840_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  and (_31841_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nor (_31842_, _31841_, _31840_);
  and (_31843_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_31844_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nor (_31845_, _31844_, _31843_);
  and (_31846_, _31845_, _31842_);
  and (_31847_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_31848_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor (_31849_, _31848_, _31847_);
  and (_31850_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  and (_31851_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nor (_31852_, _31851_, _31850_);
  and (_31853_, _31852_, _31849_);
  and (_31854_, _31853_, _31846_);
  and (_31855_, _31854_, _31839_);
  and (_31856_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  and (_31857_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nor (_31858_, _31857_, _31856_);
  and (_31859_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_31860_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nor (_31861_, _31860_, _31859_);
  and (_31862_, _31861_, _31858_);
  and (_31863_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_31864_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nor (_31865_, _31864_, _31863_);
  and (_31866_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  and (_31867_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nor (_31868_, _31867_, _31866_);
  and (_31869_, _31868_, _31865_);
  and (_31870_, _31869_, _31862_);
  and (_31871_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  and (_31872_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor (_31873_, _31872_, _31871_);
  and (_31874_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_31875_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nor (_31876_, _31875_, _31874_);
  and (_31877_, _31876_, _31873_);
  and (_31878_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_31879_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nor (_31880_, _31879_, _31878_);
  and (_31881_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  and (_31882_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nor (_31883_, _31882_, _31881_);
  and (_31884_, _31883_, _31880_);
  and (_31885_, _31884_, _31877_);
  and (_31886_, _31885_, _31870_);
  and (_31887_, _31886_, _31855_);
  and (_31888_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  and (_31889_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nor (_31890_, _31889_, _31888_);
  and (_31891_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_31892_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nor (_31893_, _31892_, _31891_);
  and (_31894_, _31893_, _31890_);
  and (_31895_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  and (_31896_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nor (_31897_, _31896_, _31895_);
  and (_31898_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_31899_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nor (_31900_, _31899_, _31898_);
  and (_31901_, _31900_, _31897_);
  and (_31902_, _31901_, _31894_);
  and (_31903_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_31904_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor (_31905_, _31904_, _31903_);
  and (_31906_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  and (_31907_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nor (_31908_, _31907_, _31906_);
  and (_31909_, _31908_, _31905_);
  and (_31910_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_31911_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor (_31912_, _31911_, _31910_);
  and (_31913_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  and (_31914_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nor (_31915_, _31914_, _31913_);
  and (_31916_, _31915_, _31912_);
  and (_31917_, _31916_, _31909_);
  and (_31918_, _31917_, _31902_);
  and (_31919_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  and (_31920_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nor (_31921_, _31920_, _31919_);
  and (_31922_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_31923_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nor (_31924_, _31923_, _31922_);
  and (_31925_, _31924_, _31921_);
  and (_31926_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  and (_31927_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor (_31928_, _31927_, _31926_);
  and (_31929_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  and (_31930_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nor (_31931_, _31930_, _31929_);
  and (_31932_, _31931_, _31928_);
  and (_31933_, _31932_, _31925_);
  and (_31934_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_31935_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nor (_31936_, _31935_, _31934_);
  and (_31937_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  and (_31938_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor (_31939_, _31938_, _31937_);
  and (_31940_, _31939_, _31936_);
  and (_31941_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_31942_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nor (_31943_, _31942_, _31941_);
  and (_31944_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  and (_31945_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nor (_31946_, _31945_, _31944_);
  and (_31947_, _31946_, _31943_);
  and (_31948_, _31947_, _31940_);
  and (_31949_, _31948_, _31933_);
  and (_31950_, _31949_, _31918_);
  and (_31951_, _31950_, _31887_);
  and (_31952_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  and (_31953_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nor (_31954_, _31953_, _31952_);
  and (_31955_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_31956_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nor (_31957_, _31956_, _31955_);
  and (_31958_, _31957_, _31954_);
  and (_31959_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  and (_31960_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nor (_31961_, _31960_, _31959_);
  and (_31962_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_31963_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nor (_31964_, _31963_, _31962_);
  and (_31965_, _31964_, _31961_);
  and (_31966_, _31965_, _31958_);
  and (_31967_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_31968_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor (_31969_, _31968_, _31967_);
  and (_31970_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_31971_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor (_31972_, _31971_, _31970_);
  and (_31973_, _31972_, _31969_);
  and (_31974_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_31975_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor (_31976_, _31975_, _31974_);
  and (_31977_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  and (_31978_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor (_31979_, _31978_, _31977_);
  and (_31980_, _31979_, _31976_);
  and (_31981_, _31980_, _31973_);
  and (_31982_, _31981_, _31966_);
  and (_31983_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  and (_31984_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor (_31985_, _31984_, _31983_);
  and (_31986_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_31987_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor (_31988_, _31987_, _31986_);
  and (_31989_, _31988_, _31985_);
  and (_31990_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  and (_31991_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor (_31992_, _31991_, _31990_);
  and (_31993_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_31994_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nor (_31995_, _31994_, _31993_);
  and (_31996_, _31995_, _31992_);
  and (_31997_, _31996_, _31989_);
  and (_31998_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_31999_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nor (_32000_, _31999_, _31998_);
  and (_32001_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  and (_32002_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor (_32003_, _32002_, _32001_);
  and (_32004_, _32003_, _32000_);
  and (_32005_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_32006_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nor (_32007_, _32006_, _32005_);
  and (_32008_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  and (_32009_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nor (_32010_, _32009_, _32008_);
  and (_32011_, _32010_, _32007_);
  and (_32012_, _32011_, _32004_);
  and (_32013_, _32012_, _31997_);
  and (_32014_, _32013_, _31982_);
  and (_32015_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  and (_32016_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nor (_32017_, _32016_, _32015_);
  and (_32018_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_32019_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nor (_32020_, _32019_, _32018_);
  and (_32021_, _32020_, _32017_);
  and (_32022_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  and (_32023_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nor (_32024_, _32023_, _32022_);
  and (_32025_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_32026_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nor (_32027_, _32026_, _32025_);
  and (_32028_, _32027_, _32024_);
  and (_32029_, _32028_, _32021_);
  and (_32030_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_32031_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor (_32032_, _32031_, _32030_);
  and (_32033_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  and (_32034_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor (_32035_, _32034_, _32033_);
  and (_32036_, _32035_, _32032_);
  and (_32037_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_32038_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor (_32039_, _32038_, _32037_);
  and (_32040_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  and (_32041_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nor (_32042_, _32041_, _32040_);
  and (_32043_, _32042_, _32039_);
  and (_32044_, _32043_, _32036_);
  and (_32045_, _32044_, _32029_);
  and (_32046_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_32047_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_32048_, _32047_, _32046_);
  and (_32049_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_32050_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_32051_, _32050_, _32049_);
  and (_32052_, _32051_, _32048_);
  and (_32053_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_32054_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_32055_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_32056_, _32055_, _32054_);
  nor (_32057_, _32056_, _32053_);
  and (_32058_, _32057_, _32052_);
  and (_32059_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_32060_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_32061_, _32060_, _32059_);
  and (_32062_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_32063_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_32064_, _32063_, _32062_);
  and (_32065_, _32064_, _32061_);
  and (_32066_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_32067_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_32068_, _32067_, _32066_);
  and (_32069_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_32070_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_32071_, _32070_, _32069_);
  and (_32072_, _32071_, _32068_);
  and (_32073_, _32072_, _32065_);
  and (_32074_, _32073_, _32058_);
  and (_32075_, _32074_, _32045_);
  and (_32076_, _32075_, _32014_);
  and (_32077_, _32076_, _31951_);
  and (_32078_, _32077_, _31824_);
  and (_32079_, _32078_, _31569_);
  nor (_32080_, _32079_, _31566_);
  or (_32081_, _32080_, _31567_);
  nor (_32082_, _30529_, _30527_);
  and (_32083_, _32079_, _21570_);
  and (_32084_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  not (_32085_, _32084_);
  and (_32086_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  and (_32087_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_32088_, _32087_, _32086_);
  and (_32089_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_32090_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or (_32091_, _32090_, _32089_);
  or (_32092_, _32091_, _32088_);
  and (_32093_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  and (_32094_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_32095_, _32094_, _32093_);
  and (_32096_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_32097_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_32098_, _32097_, _32096_);
  or (_32099_, _32098_, _32095_);
  or (_32100_, _32099_, _32092_);
  and (_32101_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  and (_32102_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_32103_, _32102_, _32101_);
  and (_32104_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  and (_32105_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_32106_, _32105_, _32104_);
  or (_32107_, _32106_, _32103_);
  and (_32108_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_32109_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_32110_, _32109_, _32108_);
  and (_32111_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  and (_32112_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_32113_, _32112_, _32111_);
  or (_32114_, _32113_, _32110_);
  or (_32115_, _32114_, _32107_);
  or (_32116_, _32115_, _32100_);
  and (_32117_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  and (_32118_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_32119_, _32118_, _32117_);
  and (_32120_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and (_32121_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_32122_, _32121_, _32120_);
  or (_32123_, _32122_, _32119_);
  and (_32124_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  and (_32125_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_32126_, _32125_, _32124_);
  and (_32127_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  and (_32128_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or (_32129_, _32128_, _32127_);
  or (_32130_, _32129_, _32126_);
  or (_32131_, _32130_, _32123_);
  and (_32132_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_32133_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_32134_, _32133_, _32132_);
  and (_32135_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_32136_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_32137_, _32136_, _32135_);
  or (_32138_, _32137_, _32134_);
  and (_32139_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and (_32140_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  or (_32141_, _32140_, _32139_);
  and (_32142_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_32143_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_32144_, _32143_, _32142_);
  or (_32145_, _32144_, _32141_);
  or (_32146_, _32145_, _32138_);
  or (_32147_, _32146_, _32131_);
  or (_32148_, _32147_, _32116_);
  and (_32149_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  and (_32150_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_32151_, _32150_, _32149_);
  and (_32152_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_32153_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_32154_, _32153_, _32152_);
  or (_32155_, _32154_, _32151_);
  and (_32156_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  and (_32157_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nor (_32158_, _32157_, _32156_);
  and (_32159_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_32160_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nor (_32161_, _32160_, _32159_);
  nand (_32162_, _32161_, _32158_);
  or (_32163_, _32162_, _32155_);
  and (_32164_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_32165_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_32166_, _32165_, _32164_);
  and (_32167_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  and (_32168_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  or (_32169_, _32168_, _32167_);
  or (_32170_, _32169_, _32166_);
  and (_32171_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  and (_32172_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_32173_, _32172_, _32171_);
  and (_32174_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_32175_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_32176_, _32175_, _32174_);
  or (_32177_, _32176_, _32173_);
  or (_32178_, _32177_, _32170_);
  or (_32179_, _32178_, _32163_);
  and (_32180_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_32181_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_32182_, _32181_, _32180_);
  and (_32183_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_32184_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_32185_, _32184_, _32183_);
  or (_32186_, _32185_, _32182_);
  and (_32187_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and (_32188_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_32189_, _32188_, _32187_);
  and (_32190_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  and (_32191_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_32192_, _32191_, _32190_);
  or (_32193_, _32192_, _32189_);
  or (_32194_, _32193_, _32186_);
  and (_32195_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_32196_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  or (_32197_, _32196_, _32195_);
  and (_32198_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_32199_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or (_32200_, _32199_, _32198_);
  or (_32201_, _32200_, _32197_);
  and (_32202_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  and (_32203_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_32204_, _32203_, _32202_);
  and (_32205_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_32206_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  or (_32207_, _32206_, _32205_);
  or (_32208_, _32207_, _32204_);
  or (_32209_, _32208_, _32201_);
  or (_32210_, _32209_, _32194_);
  or (_32211_, _32210_, _32179_);
  or (_32212_, _32211_, _32148_);
  and (_32213_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_32214_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nor (_32215_, _32214_, _32213_);
  and (_32216_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  and (_32217_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_32218_, _32217_, _32216_);
  nand (_32219_, _32218_, _32215_);
  and (_32220_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_32221_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_32222_, _32221_, _32220_);
  and (_32223_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  and (_32224_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_32225_, _32224_, _32223_);
  or (_32226_, _32225_, _32222_);
  or (_32227_, _32226_, _32219_);
  and (_32228_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_32229_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_32230_, _32229_, _32228_);
  and (_32231_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  and (_32232_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_32233_, _32232_, _32231_);
  or (_32234_, _32233_, _32230_);
  and (_32235_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_32236_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_32237_, _32236_, _32235_);
  and (_32238_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_32239_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_32240_, _32239_, _32238_);
  or (_32241_, _32240_, _32237_);
  or (_32242_, _32241_, _32234_);
  or (_32243_, _32242_, _32227_);
  and (_32244_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_32245_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_32246_, _32245_, _32244_);
  and (_32247_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_32248_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_32249_, _32248_, _32247_);
  or (_32250_, _32249_, _32246_);
  and (_32251_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  and (_32252_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_32253_, _32252_, _32251_);
  and (_32254_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_32255_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_32256_, _32255_, _32254_);
  or (_32257_, _32256_, _32253_);
  or (_32258_, _32257_, _32250_);
  and (_32259_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_32260_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_32261_, _32260_, _32259_);
  and (_32262_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_32263_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_32264_, _32263_, _32262_);
  or (_32265_, _32264_, _32261_);
  and (_32266_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  and (_32267_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_32268_, _32267_, _32266_);
  and (_32269_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_32270_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_32271_, _32270_, _32269_);
  or (_32272_, _32271_, _32268_);
  or (_32273_, _32272_, _32265_);
  or (_32274_, _32273_, _32258_);
  or (_32275_, _32274_, _32243_);
  and (_32276_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_32277_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_32278_, _32277_, _32276_);
  and (_32279_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  and (_32280_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_32281_, _32280_, _32279_);
  or (_32282_, _32281_, _32278_);
  and (_32283_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  and (_32284_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_32285_, _32284_, _32283_);
  and (_32286_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  and (_32287_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or (_32288_, _32287_, _32286_);
  or (_32289_, _32288_, _32285_);
  or (_32290_, _32289_, _32282_);
  and (_32291_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_32292_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor (_32293_, _32292_, _32291_);
  and (_32294_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  and (_32295_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor (_32296_, _32295_, _32294_);
  nand (_32297_, _32296_, _32293_);
  and (_32298_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_32299_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_32300_, _32299_, _32298_);
  and (_32301_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_32302_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_32303_, _32302_, _32301_);
  or (_32304_, _32303_, _32300_);
  or (_32305_, _32304_, _32297_);
  or (_32306_, _32305_, _32290_);
  and (_32307_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_32308_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_32309_, _32308_, _32307_);
  and (_32310_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_32311_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_32312_, _32311_, _32310_);
  or (_32313_, _32312_, _32309_);
  and (_32314_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_32315_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or (_32316_, _32315_, _32314_);
  and (_32317_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_32318_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_32319_, _32318_, _32317_);
  or (_32320_, _32319_, _32316_);
  or (_32321_, _32320_, _32313_);
  and (_32322_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_32323_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_32324_, _32323_, _32322_);
  and (_32325_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  and (_32326_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_32327_, _32326_, _32325_);
  or (_32328_, _32327_, _32324_);
  and (_32329_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  and (_32330_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_32331_, _32330_, _32329_);
  and (_32332_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_32333_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_32334_, _32333_, _32332_);
  or (_32335_, _32334_, _32331_);
  or (_32336_, _32335_, _32328_);
  or (_32337_, _32336_, _32321_);
  or (_32338_, _32337_, _32306_);
  or (_32339_, _32338_, _32275_);
  or (_32340_, _32339_, _32212_);
  and (_32341_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_32342_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_32343_, _32342_, _32341_);
  and (_32344_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_32345_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_32346_, _32345_, _32344_);
  or (_32347_, _32346_, _32343_);
  and (_32348_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  and (_32349_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_32350_, _32349_, _32348_);
  and (_32351_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_32352_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_32353_, _32352_, _32351_);
  or (_32354_, _32353_, _32350_);
  or (_32355_, _32354_, _32347_);
  and (_32356_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  and (_32357_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or (_32358_, _32357_, _32356_);
  and (_32359_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  and (_32360_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or (_32361_, _32360_, _32359_);
  or (_32362_, _32361_, _32358_);
  and (_32363_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  and (_32364_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_32365_, _32364_, _32363_);
  and (_32366_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  and (_32367_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or (_32368_, _32367_, _32366_);
  or (_32369_, _32368_, _32365_);
  or (_32370_, _32369_, _32362_);
  or (_32371_, _32370_, _32355_);
  and (_32372_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_32373_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_32374_, _32373_, _32372_);
  and (_32375_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_32376_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_32377_, _32376_, _32375_);
  or (_32378_, _32377_, _32374_);
  and (_32379_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_32380_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nor (_32381_, _32380_, _32379_);
  and (_32382_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  and (_32383_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nor (_32384_, _32383_, _32382_);
  nand (_32385_, _32384_, _32381_);
  or (_32386_, _32385_, _32378_);
  and (_32387_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  and (_32388_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_32389_, _32388_, _32387_);
  and (_32390_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_32391_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_32392_, _32391_, _32390_);
  or (_32393_, _32392_, _32389_);
  and (_32394_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_32395_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_32396_, _32395_, _32394_);
  and (_32397_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  and (_32398_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_32399_, _32398_, _32397_);
  or (_32400_, _32399_, _32396_);
  or (_32401_, _32400_, _32393_);
  or (_32402_, _32401_, _32386_);
  or (_32403_, _32402_, _32371_);
  and (_32404_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_32405_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_32406_, _32405_, _32404_);
  and (_32407_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  and (_32408_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_32409_, _32408_, _32407_);
  or (_32410_, _32409_, _32406_);
  and (_32411_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_32412_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor (_32413_, _32412_, _32411_);
  and (_32414_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  and (_32415_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nor (_32416_, _32415_, _32414_);
  nand (_32417_, _32416_, _32413_);
  or (_32418_, _32417_, _32410_);
  and (_32419_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_32420_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  and (_32421_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or (_32422_, _32421_, _32420_);
  or (_32423_, _32422_, _32419_);
  and (_32424_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and (_32425_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_32426_, _32425_, _32424_);
  and (_32427_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_32428_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or (_32429_, _32428_, _32427_);
  or (_32430_, _32429_, _32426_);
  or (_32431_, _32430_, _32423_);
  or (_32432_, _32431_, _32418_);
  and (_32433_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  and (_32434_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor (_32435_, _32434_, _32433_);
  and (_32436_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and (_32437_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nor (_32438_, _32437_, _32436_);
  nand (_32439_, _32438_, _32435_);
  and (_32440_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_32441_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  or (_32442_, _32441_, _32440_);
  and (_32443_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_32444_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_32445_, _32444_, _32443_);
  or (_32446_, _32445_, _32442_);
  or (_32447_, _32446_, _32439_);
  and (_32448_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  and (_32449_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_32450_, _32449_, _32448_);
  and (_32451_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and (_32452_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_32453_, _32452_, _32451_);
  or (_32454_, _32453_, _32450_);
  and (_32455_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and (_32456_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_32457_, _32456_, _32455_);
  and (_32458_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  and (_32459_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_32460_, _32459_, _32458_);
  or (_32461_, _32460_, _32457_);
  or (_32462_, _32461_, _32454_);
  or (_32463_, _32462_, _32447_);
  or (_32464_, _32463_, _32432_);
  or (_32465_, _32464_, _32403_);
  and (_32466_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_32467_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nor (_32468_, _32467_, _32466_);
  and (_32469_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and (_32470_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor (_32471_, _32470_, _32469_);
  nand (_32472_, _32471_, _32468_);
  and (_32473_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_32474_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_32475_, _32474_, _32473_);
  and (_32476_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_32477_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  or (_32478_, _32477_, _32476_);
  or (_32479_, _32478_, _32475_);
  or (_32480_, _32479_, _32472_);
  and (_32481_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_32482_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor (_32483_, _32482_, _32481_);
  and (_32484_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_32485_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nor (_32486_, _32485_, _32484_);
  nand (_32487_, _32486_, _32483_);
  and (_32488_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  and (_32489_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_32490_, _32489_, _32488_);
  and (_32491_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_32492_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_32493_, _32492_, _32491_);
  or (_32494_, _32493_, _32490_);
  or (_32495_, _32494_, _32487_);
  or (_32496_, _32495_, _32480_);
  and (_32497_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  and (_32498_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nor (_32499_, _32498_, _32497_);
  and (_32500_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  and (_32501_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_32502_, _32501_, _32500_);
  nand (_32503_, _32502_, _32499_);
  and (_32504_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_32505_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_32506_, _32505_, _32504_);
  and (_32507_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  and (_32508_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_32509_, _32508_, _32507_);
  or (_32510_, _32509_, _32506_);
  or (_32511_, _32510_, _32503_);
  and (_32512_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  and (_32513_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nor (_32514_, _32513_, _32512_);
  and (_32515_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_32516_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor (_32517_, _32516_, _32515_);
  nand (_32518_, _32517_, _32514_);
  and (_32519_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  and (_32520_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_32521_, _32520_, _32519_);
  and (_32522_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  and (_32523_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_32524_, _32523_, _32522_);
  or (_32525_, _32524_, _32521_);
  or (_32526_, _32525_, _32518_);
  or (_32527_, _32526_, _32511_);
  or (_32528_, _32527_, _32496_);
  and (_32529_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_32530_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_32531_, _32530_, _32529_);
  and (_32532_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_32533_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_32534_, _32533_, _32532_);
  or (_32535_, _32534_, _32531_);
  and (_32536_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  and (_32537_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_32538_, _32537_, _32536_);
  and (_32539_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_32540_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  or (_32541_, _32540_, _32539_);
  or (_32542_, _32541_, _32538_);
  or (_32543_, _32542_, _32535_);
  and (_32544_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  and (_32545_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_32546_, _32545_, _32544_);
  and (_32547_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  and (_32548_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_32549_, _32548_, _32547_);
  or (_32550_, _32549_, _32546_);
  and (_32551_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  and (_32552_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nor (_32553_, _32552_, _32551_);
  and (_32554_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_32555_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nor (_32556_, _32555_, _32554_);
  nand (_32557_, _32556_, _32553_);
  or (_32558_, _32557_, _32550_);
  or (_32559_, _32558_, _32543_);
  and (_32560_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  and (_32561_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_32562_, _32561_, _32560_);
  and (_32563_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  and (_32564_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or (_32565_, _32564_, _32563_);
  or (_32566_, _32565_, _32562_);
  and (_32567_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_32568_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_32569_, _32568_, _32567_);
  and (_32570_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_32571_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_32572_, _32571_, _32570_);
  or (_32573_, _32572_, _32569_);
  or (_32574_, _32573_, _32566_);
  and (_32575_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and (_32576_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  or (_32577_, _32576_, _32575_);
  and (_32578_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_32579_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or (_32580_, _32579_, _32578_);
  or (_32581_, _32580_, _32577_);
  and (_32582_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_32583_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_32584_, _32583_, _32582_);
  and (_32585_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and (_32586_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_32587_, _32586_, _32585_);
  or (_32588_, _32587_, _32584_);
  or (_32589_, _32588_, _32581_);
  or (_32590_, _32589_, _32574_);
  or (_32591_, _32590_, _32559_);
  or (_32592_, _32591_, _32528_);
  or (_32593_, _32592_, _32465_);
  nor (_32594_, _32593_, _32340_);
  and (_32595_, _32594_, _32085_);
  nor (_32596_, _30010_, iram_op1_reg[5]);
  nor (_32597_, _32596_, _31043_);
  and (_32598_, _32597_, _32595_);
  or (_32599_, _32598_, _32083_);
  or (_32600_, _32599_, _32082_);
  nor (_32601_, _32597_, _32595_);
  and (_32602_, _28973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  not (_32603_, _32602_);
  and (_32604_, _28848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_32605_, _28845_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor (_32606_, _32605_, _32604_);
  and (_32607_, _28852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  and (_32608_, _28855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor (_32609_, _32608_, _32607_);
  and (_32610_, _32609_, _32606_);
  and (_32611_, _28954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_32612_, _28957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nor (_32613_, _32612_, _32611_);
  and (_32614_, _28644_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_32615_, _28645_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor (_32616_, _32615_, _32614_);
  and (_32617_, _32616_, _32613_);
  and (_32618_, _32617_, _32610_);
  and (_32619_, _28916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  and (_32620_, _28915_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nor (_32621_, _32620_, _32619_);
  and (_32622_, _28545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_32623_, _28546_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nor (_32624_, _32623_, _32622_);
  and (_32625_, _32624_, _32621_);
  and (_32626_, _28846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  and (_32627_, _28894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nor (_32628_, _32627_, _32626_);
  and (_32629_, _28853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_32630_, _28856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nor (_32631_, _32630_, _32629_);
  and (_32632_, _32631_, _32628_);
  and (_32633_, _32632_, _32625_);
  and (_32634_, _32633_, _32618_);
  and (_32635_, _28564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  and (_32636_, _28563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nor (_32637_, _32636_, _32635_);
  and (_32638_, _28566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_32639_, _28892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor (_32640_, _32639_, _32638_);
  and (_32641_, _32640_, _32637_);
  and (_32642_, _28700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  and (_32643_, _28679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nor (_32644_, _32643_, _32642_);
  and (_32645_, _28895_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  and (_32646_, _28703_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nor (_32647_, _32646_, _32645_);
  and (_32648_, _32647_, _32644_);
  and (_32649_, _32648_, _32641_);
  and (_32650_, _28616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_32651_, _28891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nor (_32652_, _32651_, _32650_);
  and (_32653_, _28901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  and (_32654_, _28500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nor (_32655_, _32654_, _32653_);
  and (_32656_, _32655_, _32652_);
  and (_32657_, _28693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_32658_, _28692_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nor (_32659_, _32658_, _32657_);
  and (_32660_, _28501_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and (_32661_, _28699_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nor (_32662_, _32661_, _32660_);
  and (_32663_, _32662_, _32659_);
  and (_32664_, _32663_, _32656_);
  and (_32665_, _32664_, _32649_);
  and (_32666_, _32665_, _32634_);
  and (_32667_, _28427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_32668_, _28435_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor (_32669_, _32668_, _32667_);
  and (_32670_, _28515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and (_32671_, _28516_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nor (_32672_, _32671_, _32670_);
  and (_32673_, _32672_, _32669_);
  and (_32674_, _28806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_32675_, _28796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor (_32676_, _32675_, _32674_);
  and (_32677_, _28807_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and (_32678_, _28830_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nor (_32679_, _32678_, _32677_);
  and (_32680_, _32679_, _32676_);
  and (_32681_, _32680_, _32673_);
  and (_32682_, _28432_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and (_32683_, _28481_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nor (_32684_, _32683_, _32682_);
  and (_32685_, _28480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_32686_, _28831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nor (_32687_, _32686_, _32685_);
  and (_32688_, _32687_, _32684_);
  and (_32689_, _28803_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and (_32690_, _28450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nor (_32691_, _32690_, _32689_);
  and (_32692_, _28448_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_32693_, _28804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nor (_32694_, _32693_, _32692_);
  and (_32695_, _32694_, _32691_);
  and (_32696_, _32695_, _32688_);
  and (_32697_, _32696_, _32681_);
  and (_32698_, _28696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  and (_32699_, _28879_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nor (_32700_, _32699_, _32698_);
  and (_32701_, _28899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_32702_, _28702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nor (_32703_, _32702_, _32701_);
  and (_32704_, _32703_, _32700_);
  and (_32705_, _28717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_32706_, _28695_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nor (_32707_, _32706_, _32705_);
  and (_32708_, _28902_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  and (_32709_, _28898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nor (_32710_, _32709_, _32708_);
  and (_32711_, _32710_, _32707_);
  and (_32712_, _32711_, _32704_);
  and (_32713_, _28708_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  and (_32714_, _28677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nor (_32715_, _32714_, _32713_);
  and (_32716_, _28718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_32717_, _28714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nor (_32718_, _32717_, _32716_);
  and (_32719_, _32718_, _32715_);
  and (_32720_, _28680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  and (_32721_, _28880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor (_32722_, _32721_, _32720_);
  and (_32723_, _28876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_32724_, _28715_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor (_32725_, _32724_, _32723_);
  and (_32726_, _32725_, _32722_);
  and (_32727_, _32726_, _32719_);
  and (_32728_, _32727_, _32712_);
  and (_32729_, _32728_, _32697_);
  and (_32730_, _32729_, _32666_);
  and (_32731_, _28486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  and (_32732_, _28496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nor (_32733_, _32732_, _32731_);
  and (_32734_, _28491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_32735_, _28497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor (_32736_, _32735_, _32734_);
  and (_32737_, _32736_, _32733_);
  and (_32738_, _28474_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  and (_32739_, _28518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nor (_32740_, _32739_, _32738_);
  and (_32741_, _28799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_32742_, _28510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nor (_32743_, _32742_, _32741_);
  and (_32744_, _32743_, _32740_);
  and (_32745_, _32744_, _32737_);
  and (_32746_, _28468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_32747_, _28519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor (_32748_, _32747_, _32746_);
  and (_32749_, _28797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  and (_32750_, _28471_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor (_32751_, _32750_, _32749_);
  and (_32752_, _32751_, _32748_);
  and (_32753_, _28613_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_32754_, _28493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor (_32755_, _32754_, _32753_);
  and (_32756_, _28488_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_32757_, _28477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor (_32758_, _32757_, _32756_);
  and (_32759_, _32758_, _32755_);
  and (_32760_, _32759_, _32752_);
  and (_32761_, _32760_, _32745_);
  and (_32762_, _28636_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and (_32763_, _28637_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nor (_32764_, _32763_, _32762_);
  and (_32765_, _28639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_32766_, _28640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nor (_32767_, _32766_, _32765_);
  and (_32768_, _32767_, _32764_);
  and (_32769_, _28860_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and (_32770_, _28861_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nor (_32771_, _32770_, _32769_);
  and (_32772_, _28590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_32773_, _28947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nor (_32774_, _32773_, _32772_);
  and (_32775_, _32774_, _32771_);
  and (_32776_, _32775_, _32768_);
  and (_32777_, _28464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_32778_, _28462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nor (_32779_, _32778_, _32777_);
  and (_32780_, _28950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and (_32781_, _28570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nor (_32782_, _32781_, _32780_);
  and (_32783_, _32782_, _32779_);
  and (_32784_, _28946_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_32785_, _28589_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nor (_32786_, _32785_, _32784_);
  and (_32787_, _28578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and (_32788_, _28949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nor (_32789_, _32788_, _32787_);
  and (_32790_, _32789_, _32786_);
  and (_32791_, _32790_, _32783_);
  and (_32792_, _32791_, _32776_);
  and (_32793_, _32792_, _32761_);
  and (_32794_, _28629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_32795_, _28630_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor (_32796_, _32795_, _32794_);
  and (_32797_, _28633_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  and (_32798_, _28632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor (_32799_, _32798_, _32797_);
  and (_32800_, _32799_, _32796_);
  and (_32801_, _28652_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  and (_32802_, _28651_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nor (_32803_, _32802_, _32801_);
  and (_32804_, _28655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_32805_, _28573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nor (_32806_, _32805_, _32804_);
  and (_32807_, _32806_, _32803_);
  and (_32808_, _32807_, _32800_);
  and (_32809_, _28768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  and (_32810_, _28765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nor (_32811_, _32810_, _32809_);
  and (_32812_, _28760_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_32813_, _28767_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nor (_32814_, _32813_, _32812_);
  and (_32815_, _32814_, _32811_);
  and (_32816_, _28557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  and (_32817_, _28919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nor (_32818_, _32817_, _32816_);
  and (_32819_, _28550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_32820_, _28918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor (_32821_, _32820_, _32819_);
  and (_32822_, _32821_, _32818_);
  and (_32823_, _32822_, _32815_);
  and (_32824_, _32823_, _32808_);
  and (_32825_, _28548_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and (_32826_, _28764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nor (_32827_, _32826_, _32825_);
  and (_32828_, _28531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  and (_32829_, _28553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nor (_32830_, _32829_, _32828_);
  and (_32831_, _32830_, _32827_);
  and (_32832_, _28911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and (_32833_, _28912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nor (_32834_, _32833_, _32832_);
  and (_32835_, _28908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and (_32836_, _28909_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nor (_32837_, _32836_, _32835_);
  and (_32838_, _32837_, _32834_);
  and (_32839_, _32838_, _32831_);
  and (_32840_, _28558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  and (_32841_, _28526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nor (_32842_, _32841_, _32840_);
  and (_32843_, _28532_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and (_32844_, _28574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor (_32845_, _32844_, _32843_);
  and (_32846_, _32845_, _32842_);
  and (_32847_, _28587_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  and (_32848_, _28567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nor (_32849_, _32848_, _32847_);
  and (_32850_, _28586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and (_32851_, _28571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nor (_32852_, _32851_, _32850_);
  and (_32853_, _32852_, _32849_);
  and (_32854_, _32853_, _32846_);
  and (_32855_, _32854_, _32839_);
  and (_32856_, _32855_, _32824_);
  and (_32857_, _32856_, _32793_);
  and (_32858_, _32857_, _32730_);
  and (_32859_, _28614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  and (_32860_, _28617_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nor (_32861_, _32860_, _32859_);
  and (_32862_, _28884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_32863_, _28877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nor (_32864_, _32863_, _32862_);
  and (_32865_, _32864_, _32861_);
  and (_32866_, _28871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  and (_32867_, _28789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor (_32868_, _32867_, _32866_);
  and (_32869_, _28793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  and (_32870_, _28800_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nor (_32871_, _32870_, _32869_);
  and (_32872_, _32871_, _32868_);
  and (_32873_, _32872_, _32865_);
  and (_32874_, _28535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_32875_, _28823_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nor (_32876_, _32875_, _32874_);
  and (_32877_, _28583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  and (_32878_, _28536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nor (_32879_, _32878_, _32877_);
  and (_32880_, _32879_, _32876_);
  and (_32881_, _28456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_32882_, _28684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nor (_32883_, _32882_, _32881_);
  and (_32884_, _28453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  and (_32885_, _28683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nor (_32886_, _32885_, _32884_);
  and (_32887_, _32886_, _32883_);
  and (_32888_, _32887_, _32880_);
  and (_32889_, _32888_, _32873_);
  and (_32890_, _28602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_32891_, _28886_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor (_32892_, _32891_, _32890_);
  and (_32893_, _28883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  and (_32894_, _28887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor (_32895_, _32894_, _32893_);
  and (_32896_, _32895_, _32892_);
  and (_32897_, _28792_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_32898_, _28620_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor (_32899_, _32898_, _32897_);
  and (_32900_, _28623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_32901_, _28601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor (_32902_, _32901_, _32900_);
  and (_32903_, _32902_, _32899_);
  and (_32904_, _32903_, _32896_);
  and (_32905_, _28506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  and (_32906_, _28507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nor (_32907_, _32906_, _32905_);
  and (_32908_, _28669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_32909_, _28511_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nor (_32910_, _32909_, _32908_);
  and (_32911_, _32910_, _32907_);
  and (_32912_, _28662_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  and (_32913_, _28812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nor (_32914_, _32913_, _32912_);
  and (_32915_, _28813_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_32916_, _28665_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor (_32917_, _32916_, _32915_);
  and (_32918_, _32917_, _32914_);
  and (_32919_, _32918_, _32911_);
  and (_32920_, _32919_, _32904_);
  and (_32921_, _32920_, _32889_);
  and (_32922_, _28783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_32923_, _28782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor (_32924_, _32923_, _32922_);
  and (_32925_, _28757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  and (_32926_, _28758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor (_32927_, _32926_, _32925_);
  and (_32928_, _32927_, _32924_);
  and (_32929_, _28779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_32930_, _28780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor (_32931_, _32930_, _32929_);
  and (_32932_, _28773_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  and (_32933_, _28748_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nor (_32934_, _32933_, _32932_);
  and (_32935_, _32934_, _32931_);
  and (_32936_, _32935_, _32928_);
  and (_32937_, _28668_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  and (_32938_, _28661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nor (_32939_, _32938_, _32937_);
  and (_32940_, _28672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_32941_, _28958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor (_32942_, _32941_, _32940_);
  and (_32943_, _32942_, _32939_);
  and (_32944_, _28961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  and (_32945_, _28647_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nor (_32946_, _32945_, _32944_);
  and (_32947_, _28671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_32948_, _28648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nor (_32949_, _32948_, _32947_);
  and (_32950_, _32949_, _32946_);
  and (_32951_, _32950_, _32943_);
  and (_32952_, _32951_, _32936_);
  and (_32953_, _28964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_32954_, _28955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor (_32955_, _32954_, _32953_);
  and (_32956_, _28664_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  and (_32957_, _28815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nor (_32958_, _32957_, _32956_);
  and (_32959_, _32958_, _32955_);
  and (_32960_, _28965_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  and (_32961_, _28962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor (_32962_, _32961_, _32960_);
  and (_32963_, _28654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  and (_32964_, _28942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nor (_32965_, _32964_, _32963_);
  and (_32966_, _32965_, _32962_);
  and (_32967_, _32966_, _32959_);
  and (_32968_, _28737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  and (_32969_, _28733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor (_32970_, _32969_, _32968_);
  and (_32971_, _28736_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_32972_, _28442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nor (_32973_, _32972_, _32971_);
  and (_32974_, _32973_, _32970_);
  and (_32975_, _28749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_32976_, _28752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nor (_32977_, _32976_, _32975_);
  and (_32978_, _28734_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  and (_32979_, _28751_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nor (_32980_, _32979_, _32978_);
  and (_32981_, _32980_, _32977_);
  and (_32982_, _32981_, _32974_);
  and (_32983_, _32982_, _32967_);
  and (_32984_, _32983_, _32952_);
  and (_32985_, _32984_, _32921_);
  and (_32986_, _28606_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_32987_, _28863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor (_32988_, _32987_, _32986_);
  and (_32989_, _28790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  and (_32990_, _28864_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor (_32991_, _32990_, _32989_);
  and (_32992_, _32991_, _32988_);
  and (_32993_, _28621_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_32994_, _28599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor (_32995_, _32994_, _32993_);
  and (_32996_, _28605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  and (_32997_, _28624_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nor (_32998_, _32997_, _32996_);
  and (_32999_, _32998_, _32995_);
  and (_33000_, _32999_, _32992_);
  and (_33001_, _28827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  and (_33002_, _28744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nor (_33003_, _33002_, _33001_);
  and (_33004_, _28745_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_33005_, _28819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nor (_33006_, _33005_, _33004_);
  and (_33007_, _33006_, _33003_);
  and (_33008_, _28686_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  and (_33009_, _28676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nor (_33010_, _33009_, _33008_);
  and (_33011_, _28741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_33012_, _28687_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nor (_33013_, _33012_, _33011_);
  and (_33014_, _33013_, _33010_);
  and (_33015_, _33014_, _33007_);
  and (_33016_, _33015_, _33000_);
  and (_33017_, _28529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_33018_, _28943_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nor (_33019_, _33018_, _33017_);
  and (_33020_, _28940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  and (_33021_, _28939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nor (_33022_, _33021_, _33020_);
  and (_33023_, _33022_, _33019_);
  and (_33024_, _28742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_33025_, _28820_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nor (_33026_, _33025_, _33024_);
  and (_33027_, _28828_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  and (_33028_, _28580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nor (_33029_, _33028_, _33027_);
  and (_33030_, _33029_, _33026_);
  and (_33031_, _33030_, _33023_);
  and (_33032_, _28608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  and (_33033_, _28555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nor (_33034_, _33033_, _33032_);
  and (_33035_, _28609_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_33036_, _28597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nor (_33037_, _33036_, _33035_);
  and (_33038_, _33037_, _33034_);
  and (_33039_, _28849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  and (_33040_, _28867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nor (_33041_, _33040_, _33039_);
  and (_33042_, _28868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_33043_, _28870_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nor (_33044_, _33043_, _33042_);
  and (_33045_, _33044_, _33041_);
  and (_33046_, _33045_, _33038_);
  and (_33047_, _33046_, _33031_);
  and (_33048_, _33047_, _33016_);
  and (_33049_, _28834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  and (_33050_, _28707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nor (_33051_, _33050_, _33049_);
  and (_33052_, _28837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_33053_, _28835_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nor (_33054_, _33053_, _33052_);
  and (_33055_, _33054_, _33051_);
  and (_33056_, _28710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  and (_33057_, _28838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nor (_33058_, _33057_, _33056_);
  and (_33059_, _28822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_33060_, _28711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nor (_33061_, _33060_, _33059_);
  and (_33062_, _33061_, _33058_);
  and (_33063_, _33062_, _33055_);
  and (_33064_, _28923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_33065_, _28924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nor (_33066_, _33065_, _33064_);
  and (_33067_, _28927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  and (_33068_, _28934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor (_33069_, _33068_, _33067_);
  and (_33070_, _33069_, _33066_);
  and (_33071_, _28931_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_33072_, _28729_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor (_33073_, _33072_, _33071_);
  and (_33074_, _28933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  and (_33075_, _28930_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nor (_33076_, _33075_, _33074_);
  and (_33077_, _33076_, _33073_);
  and (_33078_, _33077_, _33070_);
  and (_33079_, _33078_, _33063_);
  and (_33080_, _28539_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_33081_, _28582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_33082_, _33081_, _33080_);
  and (_33083_, _28540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_33084_, _29456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_33085_, _33084_, _33083_);
  and (_33086_, _33085_, _33082_);
  and (_33087_, _29460_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_33088_, _29462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_33089_, _29464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_33090_, _33089_, _33088_);
  nor (_33091_, _33090_, _33087_);
  and (_33092_, _33091_, _33086_);
  and (_33093_, _28772_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_33094_, _28775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_33095_, _33094_, _33093_);
  and (_33096_, _28776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_33097_, _28926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_33098_, _33097_, _33096_);
  and (_33099_, _33098_, _33095_);
  and (_33100_, _28761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_33101_, _28727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_33102_, _33101_, _33100_);
  and (_33103_, _28730_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_33104_, _28726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_33105_, _33104_, _33103_);
  and (_33106_, _33105_, _33102_);
  and (_33107_, _33106_, _33099_);
  and (_33108_, _33107_, _33092_);
  and (_33109_, _33108_, _33079_);
  and (_33110_, _33109_, _33048_);
  and (_33111_, _33110_, _32985_);
  and (_33112_, _33111_, _32858_);
  and (_33113_, _33112_, _32603_);
  nor (_33114_, _31043_, iram_op1_reg[6]);
  nor (_33115_, _33114_, _31044_);
  nor (_33116_, _33115_, _33113_);
  or (_33117_, _33116_, _32601_);
  and (_33118_, _31047_, _31042_);
  and (_33119_, _33115_, _33113_);
  or (_33120_, _33119_, _33118_);
  or (_33121_, _33120_, _33117_);
  or (_33122_, _33121_, _32600_);
  or (_33123_, _33122_, _32081_);
  or (_33124_, _33123_, _31051_);
  and (_33125_, pc_inc_dir_r, _28439_);
  and (_33126_, _33125_, _28364_);
  and (property_invalid_inc_dir_iram, _33126_, _33124_);
  buf (_38319_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7]);
  buf (_38312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0]);
  buf (_38313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1]);
  buf (_38314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2]);
  buf (_38315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3]);
  buf (_38316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4]);
  buf (_38317_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5]);
  buf (_38318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6]);
  buf (_38996_, _39040_);
  buf (_36894_[7], _36865_[7]);
  buf (_36895_[7], _36866_[7]);
  buf (_36906_[7], _36865_[7]);
  buf (_36907_[7], _36866_[7]);
  buf (_36894_[0], _36865_[0]);
  buf (_36894_[1], _36865_[1]);
  buf (_36894_[2], _36865_[2]);
  buf (_36894_[3], _36865_[3]);
  buf (_36894_[4], _36865_[4]);
  buf (_36894_[5], _36865_[5]);
  buf (_36894_[6], _36865_[6]);
  buf (_36895_[0], _36866_[0]);
  buf (_36895_[1], _36866_[1]);
  buf (_36895_[2], _36866_[2]);
  buf (_36895_[3], _36866_[3]);
  buf (_36895_[4], _36866_[4]);
  buf (_36895_[5], _36866_[5]);
  buf (_36895_[6], _36866_[6]);
  buf (_36906_[0], _36865_[0]);
  buf (_36906_[1], _36865_[1]);
  buf (_36906_[2], _36865_[2]);
  buf (_36906_[3], _36865_[3]);
  buf (_36906_[4], _36865_[4]);
  buf (_36906_[5], _36865_[5]);
  buf (_36906_[6], _36865_[6]);
  buf (_36907_[0], _36866_[0]);
  buf (_36907_[1], _36866_[1]);
  buf (_36907_[2], _36866_[2]);
  buf (_36907_[3], _36866_[3]);
  buf (_36907_[4], _36866_[4]);
  buf (_36907_[5], _36866_[5]);
  buf (_36907_[6], _36866_[6]);
  buf (_38990_, _36880_);
  buf (_36926_, _36880_);
  dff (iram_op1[0], _00003_[0]);
  dff (iram_op1[1], _00003_[1]);
  dff (iram_op1[2], _00003_[2]);
  dff (iram_op1[3], _00003_[3]);
  dff (iram_op1[4], _00003_[4]);
  dff (iram_op1[5], _00003_[5]);
  dff (iram_op1[6], _00003_[6]);
  dff (iram_op1[7], _00003_[7]);
  dff (op1_out_r[0], _00005_[0]);
  dff (op1_out_r[1], _00005_[1]);
  dff (op1_out_r[2], _00005_[2]);
  dff (op1_out_r[3], _00005_[3]);
  dff (op1_out_r[4], _00005_[4]);
  dff (op1_out_r[5], _00005_[5]);
  dff (op1_out_r[6], _00005_[6]);
  dff (op1_out_r[7], _00005_[7]);
  dff (cy_reg, _00001_);
  dff (acc_reg[0], _00000_[0]);
  dff (acc_reg[1], _00000_[1]);
  dff (acc_reg[2], _00000_[2]);
  dff (acc_reg[3], _00000_[3]);
  dff (acc_reg[4], _00000_[4]);
  dff (acc_reg[5], _00000_[5]);
  dff (acc_reg[6], _00000_[6]);
  dff (acc_reg[7], _00000_[7]);
  dff (iram_op1_reg[0], _00004_[0]);
  dff (iram_op1_reg[1], _00004_[1]);
  dff (iram_op1_reg[2], _00004_[2]);
  dff (iram_op1_reg[3], _00004_[3]);
  dff (iram_op1_reg[4], _00004_[4]);
  dff (iram_op1_reg[5], _00004_[5]);
  dff (iram_op1_reg[6], _00004_[6]);
  dff (iram_op1_reg[7], _00004_[7]);
  dff (pc_change_r, _00006_);
  dff (pc_inc_acc_r, _00007_);
  dff (pc_inc_dir_r, _00008_);
  dff (first_instr, _00002_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _36730_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _36731_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _36732_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _36733_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _36734_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _36735_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _36736_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _36737_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _36858_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _36729_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _36729_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _36729_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _36729_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _36729_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _36729_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _36729_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _36729_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _36729_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _36729_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _36729_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _36729_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _36729_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _36729_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _36729_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _36786_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _36787_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _36788_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _36789_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _36790_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _36791_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _36792_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _36793_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _36794_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _36795_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _36796_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _36797_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _36798_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _36799_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _36800_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _36801_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _36802_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _36803_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _36804_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _36805_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _36806_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _36807_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _36808_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _36809_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _36810_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _36811_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _36812_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _36813_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _36814_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _36815_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _36816_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _36857_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _36817_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _36818_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _36819_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _36820_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _36821_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _36822_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _36823_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _36824_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _36825_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _36826_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _36827_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _36828_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _36829_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _36830_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _36831_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _36832_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _36833_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _36834_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _36835_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _36836_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _36837_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _36838_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _36839_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _36840_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _36841_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _36842_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _36843_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _36844_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _36845_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _36846_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _36847_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _36848_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _36849_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _36850_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _36851_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _36852_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _36853_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _36854_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _36855_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _36856_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _36738_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _36739_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _36740_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _36741_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _36742_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _36743_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _36744_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _36745_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _36746_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _36747_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _36748_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _36749_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _36750_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _36751_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _36752_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _36753_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _36754_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _36755_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _36756_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _36757_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _36758_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _36759_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _36760_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _36761_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _36762_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _36763_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _36764_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _36765_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _36766_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _36767_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _36768_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _36769_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _36770_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _36771_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _36772_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _36773_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _36774_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _36775_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _36776_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _36777_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _36778_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _36779_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _36780_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _36781_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _36782_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _36783_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _36784_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _36785_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _36860_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _36860_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _36860_[2]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _36860_[3]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _36860_[4]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _36860_[5]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _36859_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _36859_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _36861_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _36861_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _36861_[2]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _36861_[3]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _36861_[4]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _36861_[5]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _36861_[6]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _36861_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _36862_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _36862_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _36863_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _36863_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _36863_[2]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _36863_[3]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _36863_[4]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _36863_[5]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _36863_[6]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _36863_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _36863_[8]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _36863_[9]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _36863_[10]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _36863_[11]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _36863_[12]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _36863_[13]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _36863_[14]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _36863_[15]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _36864_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _36864_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _36864_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _36864_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _36864_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _36864_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _36864_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _36864_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _36865_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _36865_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _36865_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _36865_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _36865_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _36865_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _36865_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _36865_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _36866_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _36866_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _36866_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _36866_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _36866_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _36866_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _36866_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _36866_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _36867_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _36867_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _36867_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _36868_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _36868_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _36868_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _36869_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _36869_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _36870_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _36870_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _36870_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _36870_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _36870_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _36870_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _36870_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _36870_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _36871_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _36872_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _36872_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _36873_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _36873_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _36874_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _36874_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _36874_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _36875_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _36875_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _36875_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _36876_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _36876_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _36877_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _36877_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _36877_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _36877_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _36878_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _36878_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _36879_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _36880_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _36881_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _36881_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _36881_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _36881_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _36881_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _36881_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _36881_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _36881_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _36882_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _36882_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _36882_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _36882_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _36882_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _36882_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _36882_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _36882_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _36883_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _36883_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _36883_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _36883_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _36883_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _36883_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _36883_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _36883_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _36884_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _36884_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _36884_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _36884_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _36884_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _36884_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _36884_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _36884_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _36885_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _36885_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _36885_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _36885_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _36885_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _36885_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _36885_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _36885_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _36886_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _36886_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _36886_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _36886_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _36886_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _36886_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _36886_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _36886_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _36887_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _36887_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _36887_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _36887_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _36887_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _36887_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _36887_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _36887_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _36888_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _36888_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _36888_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _36888_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _36888_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _36888_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _36888_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _36888_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _36892_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _36892_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _36892_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _36892_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _36892_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _36889_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _36889_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _36889_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _36889_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _36889_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _36889_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _36889_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _36889_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _36889_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _36889_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _36889_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _36889_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _36889_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _36889_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _36889_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _36889_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _36890_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _36890_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _36890_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _36890_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _36890_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _36890_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _36890_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _36890_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _36890_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _36890_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _36890_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _36890_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _36890_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _36890_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _36890_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _36890_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _36913_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _36913_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _36913_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _36913_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _36913_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _36913_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _36913_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _36913_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _36913_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _36913_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _36913_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _36913_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _36913_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _36913_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _36913_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _36913_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _36913_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _36913_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _36913_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _36913_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _36913_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _36913_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _36913_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _36913_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _36913_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _36913_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _36913_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _36913_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _36913_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _36913_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _36913_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _36913_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _36891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _36893_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _36893_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _36893_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _36893_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _36893_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _36893_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _36893_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _36893_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _36894_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _36894_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _36894_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _36894_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _36894_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _36894_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _36894_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _36894_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _36895_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _36895_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _36895_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _36895_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _36895_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _36895_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _36895_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _36895_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _36896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _36897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _36898_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36898_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _36898_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _36898_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _36898_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _36898_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _36898_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _36898_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _36899_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _36899_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36899_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _36899_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _36899_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _36899_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _36899_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _36899_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _36899_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _36899_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _36899_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _36899_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _36899_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _36899_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _36899_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _36899_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _36900_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _36900_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _36900_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _36900_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _36900_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _36900_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _36900_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _36900_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _36900_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _36900_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _36900_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _36900_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _36900_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _36900_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _36900_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _36900_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _36901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _36903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _36902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _36904_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _36904_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _36904_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _36904_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _36904_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _36904_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _36904_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _36904_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _36905_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36905_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _36905_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _36906_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _36906_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _36906_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _36906_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _36906_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _36906_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _36906_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _36906_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _36907_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _36907_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _36907_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _36907_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _36907_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _36907_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _36907_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _36907_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _36908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _36909_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _36909_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _36909_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _36909_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _36909_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _36909_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _36909_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _36909_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _36910_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _36911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _36912_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _36912_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _36912_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _36912_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _36914_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _36914_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _36914_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _36914_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _36914_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _36914_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _36914_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _36914_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _36914_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _36914_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _36914_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _36914_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _36914_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _36914_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _36914_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _36914_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _36914_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _36914_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _36914_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _36914_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _36914_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _36914_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _36914_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _36914_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _36914_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _36914_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _36914_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _36914_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _36914_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _36914_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _36914_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _36914_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _36915_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _36915_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _36915_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _36915_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _36915_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _36915_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _36915_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _36915_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _36916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _36917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _36918_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _36918_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _36918_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _36918_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _36918_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _36918_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _36918_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _36918_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _36918_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _36918_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _36918_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _36918_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _36918_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _36918_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _36918_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _36918_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _36919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _36920_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _36921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _36922_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _36922_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _36922_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _36922_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _36922_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _36922_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _36922_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _36922_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _36922_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _36922_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _36922_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _36922_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _36922_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _36922_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _36922_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _36922_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _36923_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _36924_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _36925_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _36925_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _36925_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _36925_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _36925_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _36925_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _36925_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _36925_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _36926_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _36927_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _36927_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _36927_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _37136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _37137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _37138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _37139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _37140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _37141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _37142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _37143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _37128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _37129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _37130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _37131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _37132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _37133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _37134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _37135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _37120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _37121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _37122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _37123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _37124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _37125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _37126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _37127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _37112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _37113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _37114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _37115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _37116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _37117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _37118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _37119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _37096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _37097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _37098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _37099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _37100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _37101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _37102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _37103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _37088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _37089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _37090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _37091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _37092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _37093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _37094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _37095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _37080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _37081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _37082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _37083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _37084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _37085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _37086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _37087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _37072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _37073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _37074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _37075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _37076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _37077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _37078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _37079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _37184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _37185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _37186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _37187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _37188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _37189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _37190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _37191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _37064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _37065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _37066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _37067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _37068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _37069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _37070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _37071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _37056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _37057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _37058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _37059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _37060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _37061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _37062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _37063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _37048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _37049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _37050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _37051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _37052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _37053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _37054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _37055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _37040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _37041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _37042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _37043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _37044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _37045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _37046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _37047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _37032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _37033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _37034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _37035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _37036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _37037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _37038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _37039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _37024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _37025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _37026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _37027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _37028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _37029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _37030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _37031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _37008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _37009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _37010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _37011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _37012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _37013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _37014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _37015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _37000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _37001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _37002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _37003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _37004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _37005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _37006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _37007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _37200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _37201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _37202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _37203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _37204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _37205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _37206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _37207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _37272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _37273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _37274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _37275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _37276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _37277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _37278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _37279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _37264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _37265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _37266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _37267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _37268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _37269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _37270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _37271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _37256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _37257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _37258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _37259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _37260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _37261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _37262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _37263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _37480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _37481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _37482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _37483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _37484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _37485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _37486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _37487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _37472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _37473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _37474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _37475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _37476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _37477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _37478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _37479_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _37464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _37465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _37466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _37467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _37468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _37469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _37470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _37471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _37448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _37449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _37450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _37451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _37452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _37453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _37454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _37455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _37440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _37441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _37442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _37443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _37444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _37445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _37446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _37447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _37432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _37433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _37434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _37435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _37436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _37437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _37438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _37439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _37424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _37425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _37426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _37427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _37428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _37429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _37430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _37431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _37416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _37417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _37418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _37419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _37420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _37421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _37422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _37423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _37408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _37409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _37410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _37411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _37412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _37413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _37414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _37415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _37400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _37401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _37402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _37403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _37404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _37405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _37406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _37407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _37928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _37929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _37930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _37931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _37932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _37933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _37934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _37935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _37920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _37921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _37922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _37923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _37924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _37925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _37926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _37927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _37912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _37913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _37914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _37915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _37916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _37917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _37918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _37919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _37896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _37897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _37898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _37899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _37900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _37901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _37902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _37903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _37888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _37889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _37890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _37891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _37892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _37893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _37894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _37895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _37880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _37881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _37882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _37883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _37884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _37885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _37886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _37887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _37872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _37873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _37874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _37875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _37876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _37877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _37878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _37879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _37864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _37865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _37866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _37867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _37868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _37869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _37870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _37871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _38016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _38017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _38018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _38019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _38020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _38021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _38022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _38023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _38008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _38009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _38010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _38011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _38012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _38013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _38014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _38015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _38000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _38001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _38002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _38003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _38004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _38005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _38006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _38007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _37984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _37985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _37986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _37987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _37988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _37989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _37990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _37991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _37704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _37705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _37706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _37707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _37708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _37709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _37710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _37711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _38064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _38065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _38066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _38067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _38068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _38069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _38070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _38071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _38056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _38057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _38058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _38059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _38060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _38061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _38062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _38063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _37688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _37689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _37690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _37691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _37692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _37693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _37694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _37695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _37696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _37697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _37698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _37699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _37700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _37701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _37702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _37703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _37672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _37673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _37674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _37675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _37676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _37677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _37678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _37679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _37680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _37681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _37682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _37683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _37684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _37685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _37686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _37687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _37664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _37665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _37666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _37667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _37668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _37669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _37670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _37671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _37656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _37657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _37658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _37659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _37660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _37661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _37662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _37663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _37648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _37649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _37650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _37651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _37652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _37653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _37654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _37655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _37624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _37625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _37626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _37627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _37628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _37629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _37630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _37631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _37640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _37641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _37642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _37643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _37644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _37645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _37646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _37647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _37816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _37817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _37818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _37819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _37820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _37821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _37822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _37823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _36928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _36929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _36930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _36931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _36932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _36933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _36934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _36935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _38536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _38537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _38538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _38539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _38540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _38541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _38542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _38543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _38448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _38449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _38450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _38451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _38452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _38453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _38454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _38455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _38360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _38361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _38362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _38363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _38364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _38365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _38366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _38367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _38800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _38801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _38802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _38803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _38804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _38805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _38806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _38807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _38712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _38713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _38714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _38715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _38716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _38717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _38718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _38719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _38624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _38625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _38626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _38627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _38628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _38629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _38630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _38631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _38920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _38921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _38922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _38923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _38924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _38925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _38926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _38927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _38912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _38913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _38914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _38915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _38916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _38917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _38918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _38919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _38904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _38905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _38906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _38907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _38908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _38909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _38910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _38911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _38896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _38897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _38898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _38899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _38900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _38901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _38902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _38903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _38880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _38881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _38882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _38883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _38884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _38885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _38886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _38887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _38872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _38873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _38874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _38875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _38876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _38877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _38878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _38879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _38864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _38865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _38866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _38867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _38868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _38869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _38870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _38871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _38856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _38857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _38858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _38859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _38860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _38861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _38862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _38863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _38848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _38849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _38850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _38851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _38852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _38853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _38854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _38855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _38840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _38841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _38842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _38843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _38844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _38845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _38846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _38847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _38832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _38833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _38834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _38835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _38836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _38837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _38838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _38839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _38824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _38825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _38826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _38827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _38828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _38829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _38830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _38831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _38816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _38817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _38818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _38819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _38820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _38821_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _38822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _38823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _38808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _38809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _38810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _38811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _38812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _38813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _38814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _38815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _38792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _38793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _38794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _38795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _38796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _38797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _38798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _38799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _38784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _38785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _38786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _38787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _38788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _38789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _38790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _38791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _38776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _38777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _38778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _38779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _38780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _38781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _38782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _38783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _38768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _38769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _38770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _38771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _38772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _38773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _38774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _38775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _38760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _38761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _38762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _38763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _38764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _38765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _38766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _38767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _38752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _38753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _38754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _38755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _38756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _38757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _38758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _38759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _38744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _38745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _38746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _38747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _38748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _38749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _38750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _38751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _38736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _38737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _38738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _38739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _38740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _38741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _38742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _38743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _38728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _38729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _38730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _38731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _38732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _38733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _38734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _38735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _38720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _38721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _38722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _38723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _38724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _38725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _38726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _38727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _38704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _38705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _38706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _38707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _38708_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _38709_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _38710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _38711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _38696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _38697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _38698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _38699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _38700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _38701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _38702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _38703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _38688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _38689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _38690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _38691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _38692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _38693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _38694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _38695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _38680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _38681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _38682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _38683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _38684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _38685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _38686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _38687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _38672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _38673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _38674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _38675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _38676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _38677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _38678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _38679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _38664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _38665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _38666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _38667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _38668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _38669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _38670_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _38671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _38656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _38657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _38658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _38659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _38660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _38661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _38662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _38663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _38648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _38649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _38650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _38651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _38652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _38653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _38654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _38655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _38640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _38641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _38642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _38643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _38644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _38645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _38646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _38647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _38632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _38633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _38634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _38635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _38636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _38637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _38638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _38639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _38616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _38617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _38618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _38619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _38620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _38621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _38622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _38623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _38608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _38609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _38610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _38611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _38612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _38613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _38614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _38615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _38600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _38601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _38602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _38603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _38604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _38605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _38606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _38607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _38592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _38593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _38594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _38595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _38596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _38597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _38598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _38599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _38584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _38585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _38586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _38587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _38588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _38589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _38590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _38591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _38576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _38577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _38578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _38579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _38580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _38581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _38582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _38583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _38568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _38569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _38570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _38571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _38572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _38573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _38574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _38575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _38560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _38561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _38562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _38563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _38564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _38565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _38566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _38567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _38552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _38553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _38554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _38555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _38556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _38557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _38558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _38559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _38544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _38545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _38546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _38547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _38548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _38549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _38550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _38551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _38528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _38529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _38530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _38531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _38532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _38533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _38534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _38535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _38520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _38521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _38522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _38523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _38524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _38525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _38526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _38527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _38512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _38513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _38514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _38515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _38516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _38517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _38518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _38519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _38504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _38505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _38506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _38507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _38508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _38509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _38510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _38511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _38496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _38497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _38498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _38499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _38500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _38501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _38502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _38503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _38488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _38489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _38490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _38491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _38492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _38493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _38494_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _38495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _38480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _38481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _38482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _38483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _38484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _38485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _38486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _38487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _38472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _38473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _38474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _38475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _38476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _38477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _38478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _38479_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _38464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _38465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _38466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _38467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _38468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _38469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _38470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _38471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _38456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _38457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _38458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _38459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _38460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _38461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _38462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _38463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _38440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _38441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _38442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _38443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _38444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _38445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _38446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _38447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _38432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _38433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _38434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _38435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _38436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _38437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _38438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _38439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _38424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _38425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _38426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _38427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _38428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _38429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _38430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _38431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _38416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _38417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _38418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _38419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _38420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _38421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _38422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _38423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _38408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _38409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _38410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _38411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _38412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _38413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _38414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _38415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _38400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _38401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _38402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _38403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _38404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _38405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _38406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _38407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _38392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _38393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _38394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _38395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _38396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _38397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _38398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _38399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _38384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _38385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _38386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _38387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _38388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _38389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _38390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _38391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _38376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _38377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _38378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _38379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _38380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _38381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _38382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _38383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _38368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _38369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _38370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _38371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _38372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _38373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _38374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _38375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _38352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _38353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _38354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _38355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _38356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _38357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _38358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _38359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _38344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _38345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _38346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _38347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _38348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _38349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _38350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _38351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _38336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _38337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _38338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _38339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _38340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _38341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _38342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _38343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _38328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _38329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _38330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _38331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _38332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _38333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _38334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _38335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _38320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _38321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _38322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _38323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _38324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _38325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _38326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _38327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _38256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _38257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _38258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _38259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _38260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _38261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _38262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _38263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _38168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _38169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _38170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _38171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _38172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _38173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _38174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _38175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _38080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _38081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _38082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _38083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _38084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _38085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _38086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _38087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _37992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _37993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _37994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _37995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _37996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _37997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _37998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _37999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _37904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _37905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _37906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _37907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _37908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _37909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _37910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _37911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _37808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _37809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _37810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _37811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _37812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _37813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _37814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _37815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _37720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _37721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _37722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _37723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _37724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _37725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _37726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _37727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _37632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _37633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _37634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _37635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _37636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _37637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _37638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _37639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _37544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _37545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _37546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _37547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _37548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _37549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _37550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _37551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _37456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _37457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _37458_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _37459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _37460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _37461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _37462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _37463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _37368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _37369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _37370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _37371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _37372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _37373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _37374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _37375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _37280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _37281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _37282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _37283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _37284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _37285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _37286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _37287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _37192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _37193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _37194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _37195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _37196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _37197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _37198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _37199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _37104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _37105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _37106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _37107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _37108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _37109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _37110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _37111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _37016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _37017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _37018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _37019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _37020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _37021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _37022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _37023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _38976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _38977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _38978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _38979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _38980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _38981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _38982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _38983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _38888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _38889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _38890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _38891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _38892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _38893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _38894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _38895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _38048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _38049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _38050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _38051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _38052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _38053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _38054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _38055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _37976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _37977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _37978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _37979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _37980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _37981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _37982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _37983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _37856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _37857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _37858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _37859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _37860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _37861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _37862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _37863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _37848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _37849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _37850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _37851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _37852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _37853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _37854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _37855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _37840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _37841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _37842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _37843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _37844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _37845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _37846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _37847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _37832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _37833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _37834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _37835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _37836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _37837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _37838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _37839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _37824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _37825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _37826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _37827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _37828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _37829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _37830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _37831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _37800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _37801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _37802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _37803_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _37804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _37805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _37806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _37807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _37792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _37793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _37794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _37795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _37796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _37797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _37798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _37799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _37784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _37785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _37786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _37787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _37788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _37789_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _37790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _37791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _37776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _37777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _37778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _37779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _37780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _37781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _37782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _37783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _37768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _37769_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _37770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _37771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _37772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _37773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _37774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _37775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _37760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _37761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _37762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _37763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _37764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _37765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _37766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _37767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _37752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _37753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _37754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _37755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _37756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _37757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _37758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _37759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _37744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _37745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _37746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _37747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _37748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _37749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _37750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _37751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _37736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _37737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _37738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _37739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _37740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _37741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _37742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _37743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _37728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _37729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _37730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _37731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _37732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _37733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _37734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _37735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _37712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _37713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _37714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _37715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _37716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _37717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _37718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _37719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _37392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _37393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _37394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _37395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _37396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _37397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _37398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _37399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _37512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _37513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _37514_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _37515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _37516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _37517_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _37518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _37519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _37384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _37385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _37386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _37387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _37388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _37389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _37390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _37391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _37504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _37505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _37506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _37507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _37508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _37509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _37510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _37511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _37376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _37377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _37378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _37379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _37380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _37381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _37382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _37383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _37496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _37497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _37498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _37499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _37500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _37501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _37502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _37503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _37360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _37361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _37362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _37363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _37364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _37365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _37366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _37367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _37488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _37489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _37490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _37491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _37492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _37493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _37494_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _37495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _37352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _37353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _37354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _37355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _37356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _37357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _37358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _37359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _37344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _37345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _37346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _37347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _37348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _37349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _37350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _37351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _37336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _37337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _37338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _37339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _37340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _37341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _37342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _37343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _37328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _37329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _37330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _37331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _37332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _37333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _37334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _37335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _37320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _37321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _37322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _37323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _37324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _37325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _37326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _37327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _37312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _37313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _37314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _37315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _37316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _37317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _37318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _37319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _37304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _37305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _37306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _37307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _37308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _37309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _37310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _37311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _37296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _37297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _37298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _37299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _37300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _37301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _37302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _37303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _37288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _37289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _37290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _37291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _37292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _37293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _37294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _37295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _37248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _37249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _37250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _37251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _37252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _37253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _37254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _37255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _36992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _36993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _36994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _36995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _36996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _36997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _36998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _36999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _36984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _36985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _36986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _36987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _36988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _36989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _36990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _36991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _36976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _36977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _36978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _36979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _36980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _36981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _36982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _36983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _36968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _36969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _36970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _36971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _36972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _36973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _36974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _36975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _36960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _36961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _36962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _36963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _36964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _36965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _36966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _36967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _37176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _37177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _37178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _37179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _37180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _37181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _37182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _37183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _36952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _36953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _36954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _36955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _36956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _36957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _36958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _36959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _36944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _36945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _36946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _36947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _36948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _36949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _36950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _36951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _36936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _36937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _36938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _36939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _36940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _36941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _36942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _36943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _38968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _38969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _38970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _38971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _38972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _38973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _38974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _38975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _38960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _38961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _38962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _38963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _38964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _38965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _38966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _38967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _37168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _37169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _37170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _37171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _37172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _37173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _37174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _37175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _38952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _38953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _38954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _38955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _38956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _38957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _38958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _38959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _38944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _38945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _38946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _38947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _38948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _38949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _38950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _38951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _37160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _37161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _37162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _37163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _37164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _37165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _37166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _37167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _38936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _38937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _38938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _38939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _38940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _38941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _38942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _38943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _38928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _38929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _38930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _38931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _38932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _38933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _38934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _38935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _38232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _38233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _38234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _38235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _38236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _38237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _38238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _38239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _38240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _38241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _38242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _38243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _38244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _38245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _38246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _38247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _38136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _38137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _38138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _38139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _38140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _38141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _38142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _38143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _38144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _38145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _38146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _38147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _38148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _38149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _38150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _38151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _37944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _37945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _37946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _37947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _37948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _37949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _37950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _37951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _37616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _37617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _37618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _37619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _37620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _37621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _37622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _37623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _37552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _37553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _37554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _37555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _37556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _37557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _37558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _37559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _37152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _37153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _37154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _37155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _37156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _37157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _37158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _37159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _37144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _37145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _37146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _37147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _37148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _37149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _37150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _37151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _37608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _37609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _37610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _37611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _37612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _37613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _37614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _37615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _37592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _37593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _37594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _37595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _37596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _37597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _37598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _37599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _37600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _37601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _37602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _37603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _37604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _37605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _37606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _37607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _37576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _37577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _37578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _37579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _37580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _37581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _37582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _37583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _37584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _37585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _37586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _37587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _37588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _37589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _37590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _37591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _37560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _37561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _37562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _37563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _37564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _37565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _37566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _37567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _37568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _37569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _37570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _37571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _37572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _37573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _37574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _37575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _37536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _37537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _37538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _37539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _37540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _37541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _37542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _37543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _37528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _37529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _37530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _37531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _37532_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _37533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _37534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _37535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _37520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _37521_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _37522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _37523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _37524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _37525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _37526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _37527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _37232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _37233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _37234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _37235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _37236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _37237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _37238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _37239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _37240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _37241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _37242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _37243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _37244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _37245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _37246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _37247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _37224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _37225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _37226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _37227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _37228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _37229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _37230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _37231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _37216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _37217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _37218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _37219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _37220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _37221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _37222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _37223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _37208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _37209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _37210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _37211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _37212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _37213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _37214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _37215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [0], _38312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [1], _38313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [2], _38314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [3], _38315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [4], _38316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [5], _38317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [6], _38318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[256] [7], _38319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _38304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _38305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _38306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _38307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _38308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _38309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _38310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _38311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _38288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _38289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _38290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _38291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _38292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _38293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _38294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _38295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _38296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _38297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _38298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _38299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _38300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _38301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _38302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _38303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _38280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _38281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _38282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _38283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _38284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _38285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _38286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _38287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _38272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _38273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _38274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _38275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _38276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _38277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _38278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _38279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _38248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _38249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _38250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _38251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _38252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _38253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _38254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _38255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _38264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _38265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _38266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _38267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _38268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _38269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _38270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _38271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _38224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _38225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _38226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _38227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _38228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _38229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _38230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _38231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _38216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _38217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _38218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _38219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _38220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _38221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _38222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _38223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _38200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _38201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _38202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _38203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _38204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _38205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _38206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _38207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _38208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _38209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _38210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _38211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _38212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _38213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _38214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _38215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _38192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _38193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _38194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _38195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _38196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _38197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _38198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _38199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _38184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _38185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _38186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _38187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _38188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _38189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _38190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _38191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _38176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _38177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _38178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _38179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _38180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _38181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _38182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _38183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _38160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _38161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _38162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _38163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _38164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _38165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _38166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _38167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _38152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _38153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _38154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _38155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _38156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _38157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _38158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _38159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _38120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _38121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _38122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _38123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _38124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _38125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _38126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _38127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _38128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _38129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _38130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _38131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _38132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _38133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _38134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _38135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _38112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _38113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _38114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _38115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _38116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _38117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _38118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _38119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _38104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _38105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _38106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _38107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _38108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _38109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _38110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _38111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _38096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _38097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _38098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _38099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _38100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _38101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _38102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _38103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _38088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _38089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _38090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _38091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _38092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _38093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _38094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _38095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _38072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _38073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _38074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _38075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _38076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _38077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _38078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _38079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _38040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _38041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _38042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _38043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _38044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _38045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _38046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _38047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _38032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _38033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _38034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _38035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _38036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _38037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _38038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _38039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _38024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _38025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _38026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _38027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _38028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _38029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _38030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _38031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _37936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _37937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _37938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _37939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _37940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _37941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _37942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _37943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _37968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _37969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _37970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _37971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _37972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _37973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _37974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _37975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _37952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _37953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _37954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _37955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _37956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _37957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _37958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _37959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _37960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _37961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _37962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _37963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _37964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _37965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _37966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _37967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _38984_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _38984_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _38984_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _38984_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _38984_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _38984_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _38984_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _38984_[7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _38985_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _38986_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _38986_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _38986_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _38986_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _38987_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _38988_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _38989_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _38989_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _38989_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _38989_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _38989_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _38989_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _38989_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _38989_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _38990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _38991_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _38991_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _38991_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _38991_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _38991_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _38991_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _38991_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _38991_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _38992_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _38992_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _38992_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _38992_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _38992_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _38992_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _38992_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _38992_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _38993_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _38993_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _38993_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _38993_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _38993_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _38993_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _38993_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _38993_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _38994_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _38994_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _38994_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _38994_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _38994_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _38994_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _38994_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _38994_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _38995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _38996_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _38997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _38998_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _38998_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _38998_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _38998_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _38998_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _38998_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _38998_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _38998_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _38999_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _38999_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _39000_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _39001_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _39001_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _39001_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _39002_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _39002_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _39002_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _39003_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _39003_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _39004_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _39004_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _39005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _39006_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _39007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _39008_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _39009_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _39009_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _39009_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39009_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _39010_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _39010_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _39010_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _39010_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _39010_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _39010_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _39010_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _39010_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _39011_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _39011_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _39011_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _39011_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _39011_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _39011_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _39011_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _39011_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _39012_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _39012_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _39012_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _39012_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _39012_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _39012_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _39012_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _39012_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _39013_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _39013_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _39013_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _39013_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _39013_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _39013_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _39013_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _39013_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _39014_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _39014_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _39014_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _39014_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _39014_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _39014_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _39014_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _39014_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _39015_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _39015_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _39015_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _39015_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _39015_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _39015_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _39015_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _39015_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _39016_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _39016_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _39016_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _39016_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _39016_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _39016_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _39016_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _39017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _39018_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _39018_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _39018_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _39018_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _39018_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _39018_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _39018_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _39018_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39020_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _39021_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _39021_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _39021_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _39021_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _39021_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _39021_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _39021_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _39021_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _39022_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _39022_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _39022_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _39022_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _39022_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _39022_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _39022_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _39022_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _39023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _39024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _39025_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _39025_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _39025_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _39025_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _39025_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _39025_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _39025_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _39025_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _39026_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _39026_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _39026_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _39026_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _39026_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _39026_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _39026_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _39026_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _39027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _39028_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _39028_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _39028_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _39028_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39028_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _39028_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _39028_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _39028_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _39029_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _39030_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _39031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _39032_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _39033_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _39033_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _39033_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _39033_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _39033_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _39033_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _39033_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _39033_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _39034_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _39034_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _39034_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _39034_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _39034_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _39034_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _39034_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _39034_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _39035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _39036_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _39036_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _39036_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _39036_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _39036_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _39036_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _39036_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _39036_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _39037_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _39037_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _39037_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _39037_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _39037_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _39037_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _39037_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _39037_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _39038_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _39039_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _39039_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _39039_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _39039_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _39039_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _39039_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _39039_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _39039_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _39049_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _39049_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _39049_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _39049_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _39049_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _39049_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _39049_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _39049_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _39049_[8]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _39049_[9]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _39049_[10]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _39049_[11]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _39040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _39041_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _39042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _39043_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _39044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _39045_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _39046_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _39046_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _39047_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _39047_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _39047_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _39047_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _39048_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _39048_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _39048_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _39048_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _39048_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _39048_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _39048_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _39048_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _39050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _39051_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _39052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _39053_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _39054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _39055_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _39055_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _39055_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _39055_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _39056_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _39056_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _39056_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _39056_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _39056_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _39056_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _39056_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _39056_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _39056_[8]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _39056_[9]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _39056_[10]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _39057_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _39057_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _39057_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _39057_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _39057_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _39057_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _39057_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _39057_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _39058_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _39058_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _39058_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _39058_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _39058_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _39058_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _39058_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _39058_[7]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 );
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 );
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.uart_int , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tc2_int , \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
