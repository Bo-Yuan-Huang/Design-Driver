
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire [7:0] _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  input [34:0] ABINPUT;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire eq_state;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire \oc8051_golden_model_1.n1046 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire \oc8051_golden_model_1.n1063 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1157 ;
  wire [3:0] \oc8051_golden_model_1.n1159 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire [3:0] \oc8051_golden_model_1.n1167 ;
  wire \oc8051_golden_model_1.n1214 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [2:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1265 ;
  wire [1:0] \oc8051_golden_model_1.n1266 ;
  wire [7:0] \oc8051_golden_model_1.n1267 ;
  wire [6:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1276 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire [7:0] \oc8051_golden_model_1.n1284 ;
  wire \oc8051_golden_model_1.n1300 ;
  wire [7:0] \oc8051_golden_model_1.n1301 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1360 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [8:0] \oc8051_golden_model_1.n1367 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [4:0] \oc8051_golden_model_1.n1374 ;
  wire \oc8051_golden_model_1.n1375 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire \oc8051_golden_model_1.n1384 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire \oc8051_golden_model_1.n1401 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [8:0] \oc8051_golden_model_1.n1424 ;
  wire \oc8051_golden_model_1.n1425 ;
  wire [4:0] \oc8051_golden_model_1.n1430 ;
  wire \oc8051_golden_model_1.n1431 ;
  wire \oc8051_golden_model_1.n1439 ;
  wire [7:0] \oc8051_golden_model_1.n1440 ;
  wire [6:0] \oc8051_golden_model_1.n1441 ;
  wire \oc8051_golden_model_1.n1456 ;
  wire [7:0] \oc8051_golden_model_1.n1457 ;
  wire [8:0] \oc8051_golden_model_1.n1459 ;
  wire [8:0] \oc8051_golden_model_1.n1461 ;
  wire \oc8051_golden_model_1.n1462 ;
  wire [3:0] \oc8051_golden_model_1.n1463 ;
  wire [4:0] \oc8051_golden_model_1.n1464 ;
  wire [4:0] \oc8051_golden_model_1.n1466 ;
  wire \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1468 ;
  wire \oc8051_golden_model_1.n1475 ;
  wire [7:0] \oc8051_golden_model_1.n1476 ;
  wire [6:0] \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [7:0] \oc8051_golden_model_1.n1493 ;
  wire [8:0] \oc8051_golden_model_1.n1496 ;
  wire \oc8051_golden_model_1.n1497 ;
  wire \oc8051_golden_model_1.n1504 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [8:0] \oc8051_golden_model_1.n1509 ;
  wire [8:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [4:0] \oc8051_golden_model_1.n1513 ;
  wire [4:0] \oc8051_golden_model_1.n1515 ;
  wire \oc8051_golden_model_1.n1516 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1524 ;
  wire [7:0] \oc8051_golden_model_1.n1525 ;
  wire [6:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [4:0] \oc8051_golden_model_1.n1544 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [6:0] \oc8051_golden_model_1.n1547 ;
  wire [7:0] \oc8051_golden_model_1.n1548 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [7:0] \oc8051_golden_model_1.n1559 ;
  wire [6:0] \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [6:0] \oc8051_golden_model_1.n1563 ;
  wire [7:0] \oc8051_golden_model_1.n1564 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire [8:0] \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire \oc8051_golden_model_1.n1586 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire [8:0] \oc8051_golden_model_1.n1593 ;
  wire \oc8051_golden_model_1.n1594 ;
  wire [4:0] \oc8051_golden_model_1.n1595 ;
  wire [4:0] \oc8051_golden_model_1.n1597 ;
  wire \oc8051_golden_model_1.n1598 ;
  wire \oc8051_golden_model_1.n1605 ;
  wire [7:0] \oc8051_golden_model_1.n1606 ;
  wire [6:0] \oc8051_golden_model_1.n1607 ;
  wire \oc8051_golden_model_1.n1622 ;
  wire [7:0] \oc8051_golden_model_1.n1623 ;
  wire [8:0] \oc8051_golden_model_1.n1627 ;
  wire \oc8051_golden_model_1.n1628 ;
  wire [4:0] \oc8051_golden_model_1.n1630 ;
  wire \oc8051_golden_model_1.n1631 ;
  wire \oc8051_golden_model_1.n1638 ;
  wire [7:0] \oc8051_golden_model_1.n1639 ;
  wire [6:0] \oc8051_golden_model_1.n1640 ;
  wire \oc8051_golden_model_1.n1655 ;
  wire [7:0] \oc8051_golden_model_1.n1656 ;
  wire [8:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire [4:0] \oc8051_golden_model_1.n1663 ;
  wire \oc8051_golden_model_1.n1664 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire [7:0] \oc8051_golden_model_1.n1672 ;
  wire [6:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1688 ;
  wire [7:0] \oc8051_golden_model_1.n1689 ;
  wire [8:0] \oc8051_golden_model_1.n1693 ;
  wire \oc8051_golden_model_1.n1694 ;
  wire [4:0] \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1697 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire [6:0] \oc8051_golden_model_1.n1706 ;
  wire \oc8051_golden_model_1.n1721 ;
  wire [7:0] \oc8051_golden_model_1.n1722 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire [6:0] \oc8051_golden_model_1.n1748 ;
  wire [7:0] \oc8051_golden_model_1.n1749 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1821 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1838 ;
  wire [7:0] \oc8051_golden_model_1.n1839 ;
  wire \oc8051_golden_model_1.n1855 ;
  wire [7:0] \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1879 ;
  wire [6:0] \oc8051_golden_model_1.n1880 ;
  wire [7:0] \oc8051_golden_model_1.n1881 ;
  wire \oc8051_golden_model_1.n1936 ;
  wire [7:0] \oc8051_golden_model_1.n1937 ;
  wire \oc8051_golden_model_1.n1953 ;
  wire [7:0] \oc8051_golden_model_1.n1954 ;
  wire \oc8051_golden_model_1.n1970 ;
  wire [7:0] \oc8051_golden_model_1.n1971 ;
  wire \oc8051_golden_model_1.n1987 ;
  wire [7:0] \oc8051_golden_model_1.n1988 ;
  wire \oc8051_golden_model_1.n2085 ;
  wire [7:0] \oc8051_golden_model_1.n2086 ;
  wire \oc8051_golden_model_1.n2102 ;
  wire [7:0] \oc8051_golden_model_1.n2103 ;
  wire \oc8051_golden_model_1.n2119 ;
  wire [7:0] \oc8051_golden_model_1.n2120 ;
  wire \oc8051_golden_model_1.n2136 ;
  wire [7:0] \oc8051_golden_model_1.n2137 ;
  wire \oc8051_golden_model_1.n2141 ;
  wire [6:0] \oc8051_golden_model_1.n2142 ;
  wire [7:0] \oc8051_golden_model_1.n2143 ;
  wire [6:0] \oc8051_golden_model_1.n2144 ;
  wire [7:0] \oc8051_golden_model_1.n2145 ;
  wire \oc8051_golden_model_1.n2160 ;
  wire [7:0] \oc8051_golden_model_1.n2161 ;
  wire \oc8051_golden_model_1.n2200 ;
  wire [7:0] \oc8051_golden_model_1.n2201 ;
  wire [6:0] \oc8051_golden_model_1.n2202 ;
  wire [7:0] \oc8051_golden_model_1.n2203 ;
  wire [3:0] \oc8051_golden_model_1.n2210 ;
  wire \oc8051_golden_model_1.n2211 ;
  wire [7:0] \oc8051_golden_model_1.n2212 ;
  wire [6:0] \oc8051_golden_model_1.n2213 ;
  wire \oc8051_golden_model_1.n2228 ;
  wire [7:0] \oc8051_golden_model_1.n2229 ;
  wire [7:0] \oc8051_golden_model_1.n2441 ;
  wire \oc8051_golden_model_1.n2444 ;
  wire \oc8051_golden_model_1.n2446 ;
  wire \oc8051_golden_model_1.n2452 ;
  wire [7:0] \oc8051_golden_model_1.n2453 ;
  wire [6:0] \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire \oc8051_golden_model_1.n2474 ;
  wire \oc8051_golden_model_1.n2476 ;
  wire \oc8051_golden_model_1.n2482 ;
  wire [7:0] \oc8051_golden_model_1.n2483 ;
  wire [6:0] \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire \oc8051_golden_model_1.n2504 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire \oc8051_golden_model_1.n2512 ;
  wire [7:0] \oc8051_golden_model_1.n2513 ;
  wire [6:0] \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire \oc8051_golden_model_1.n2534 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire \oc8051_golden_model_1.n2559 ;
  wire [7:0] \oc8051_golden_model_1.n2560 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire [6:0] \oc8051_golden_model_1.n2564 ;
  wire [7:0] \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire [7:0] \oc8051_golden_model_1.n2568 ;
  wire [15:0] \oc8051_golden_model_1.n2572 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire [6:0] \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire [7:0] \oc8051_golden_model_1.n2600 ;
  wire [6:0] \oc8051_golden_model_1.n2601 ;
  wire [7:0] \oc8051_golden_model_1.n2602 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire \oc8051_golden_model_1.n2666 ;
  wire [7:0] \oc8051_golden_model_1.n2667 ;
  wire [6:0] \oc8051_golden_model_1.n2668 ;
  wire [7:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [6:0] \oc8051_golden_model_1.n2695 ;
  wire [7:0] \oc8051_golden_model_1.n2696 ;
  wire [3:0] \oc8051_golden_model_1.n2697 ;
  wire [7:0] \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2713 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire [7:0] \oc8051_golden_model_1.n2734 ;
  wire [6:0] \oc8051_golden_model_1.n2735 ;
  wire \oc8051_golden_model_1.n2750 ;
  wire [7:0] \oc8051_golden_model_1.n2751 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2756 ;
  wire \oc8051_golden_model_1.n2757 ;
  wire \oc8051_golden_model_1.n2758 ;
  wire \oc8051_golden_model_1.n2759 ;
  wire \oc8051_golden_model_1.n2766 ;
  wire [7:0] \oc8051_golden_model_1.n2767 ;
  wire \oc8051_golden_model_1.n2768 ;
  wire \oc8051_golden_model_1.n2769 ;
  wire \oc8051_golden_model_1.n2770 ;
  wire \oc8051_golden_model_1.n2771 ;
  wire \oc8051_golden_model_1.n2772 ;
  wire \oc8051_golden_model_1.n2773 ;
  wire \oc8051_golden_model_1.n2774 ;
  wire \oc8051_golden_model_1.n2775 ;
  wire \oc8051_golden_model_1.n2782 ;
  wire [7:0] \oc8051_golden_model_1.n2783 ;
  wire [7:0] \oc8051_golden_model_1.n2815 ;
  wire [6:0] \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire [7:0] \oc8051_golden_model_1.n2837 ;
  wire [6:0] \oc8051_golden_model_1.n2838 ;
  wire \oc8051_golden_model_1.n2853 ;
  wire [7:0] \oc8051_golden_model_1.n2854 ;
  wire [7:0] \oc8051_golden_model_1.n2858 ;
  wire [3:0] \oc8051_golden_model_1.n2859 ;
  wire [7:0] \oc8051_golden_model_1.n2860 ;
  wire \oc8051_golden_model_1.n2861 ;
  wire \oc8051_golden_model_1.n2862 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2865 ;
  wire \oc8051_golden_model_1.n2866 ;
  wire \oc8051_golden_model_1.n2867 ;
  wire \oc8051_golden_model_1.n2868 ;
  wire \oc8051_golden_model_1.n2875 ;
  wire [7:0] \oc8051_golden_model_1.n2876 ;
  wire \oc8051_golden_model_1.n2894 ;
  wire [7:0] \oc8051_golden_model_1.n2895 ;
  wire [7:0] \oc8051_golden_model_1.n2896 ;
  wire \oc8051_golden_model_1.n2912 ;
  wire [7:0] \oc8051_golden_model_1.n2913 ;
  wire [7:0] \oc8051_golden_model_1.n2914 ;
  wire \oc8051_golden_model_1.rst ;
  wire [34:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.des1 ;
  wire [7:0] \oc8051_top_1.des2 ;
  wire \oc8051_top_1.desAc ;
  wire \oc8051_top_1.desCy ;
  wire \oc8051_top_1.desOv ;
  wire [7:0] \oc8051_top_1.des_acc ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.des ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.data_in ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.alu ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des_acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_dat ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_in ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat2 ;
  wire \oc8051_top_1.oc8051_sfr1.desAc ;
  wire \oc8051_top_1.oc8051_sfr1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.des_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire [7:0] \oc8051_top_1.sub_result ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire [7:0] \oc8051_top_1.wr_dat ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire p1_valid_r;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire property_valid_psw_1_r;
  wire property_valid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  wire regs_always_zero;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_39026_, rst);
  not (_15675_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_15686_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15697_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15686_);
  and (_15708_, _15697_, _15675_);
  and (_15719_, \oc8051_top_1.oc8051_decoder1.wr , _15686_);
  not (_15730_, _15719_);
  nor (_15741_, _15730_, _15708_);
  and (_15752_, _15741_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_15763_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_15774_, _15763_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_15785_, _15774_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_15796_, _15785_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_15807_, _15796_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_15817_, _15807_);
  and (_15828_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15686_);
  and (_15839_, _15828_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_15850_, _15839_, _15675_);
  not (_15861_, _15850_);
  nor (_15872_, _15796_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_15883_, _15872_, _15861_);
  and (_15894_, _15883_, _15817_);
  not (_15904_, _15894_);
  and (_15915_, _15839_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_15926_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_15937_, _15828_, _15926_);
  and (_15948_, _15937_, _15675_);
  and (_15959_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_15970_, _15959_, _15915_);
  nor (_15981_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_15992_, _15981_, _15697_);
  and (_16002_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_16013_, _15937_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_16034_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_16035_, _16034_, _16002_);
  and (_16046_, _16035_, _15970_);
  and (_16057_, _16046_, _15904_);
  and (_16068_, _15807_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_16079_, _16068_);
  nor (_16089_, _15807_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_16100_, _16089_, _15861_);
  and (_16111_, _16100_, _16079_);
  not (_16122_, _16111_);
  and (_16133_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_16144_, _16133_, _15915_);
  and (_16155_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_16166_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_16177_, _16166_, _16155_);
  and (_16187_, _16177_, _16144_);
  and (_16198_, _16187_, _16122_);
  nor (_16209_, _16198_, _16057_);
  not (_16220_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_16231_, _16068_, _16220_);
  and (_16242_, _16068_, _16220_);
  nor (_16253_, _16242_, _16231_);
  nor (_16264_, _16253_, _15861_);
  not (_16275_, _16264_);
  and (_16285_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_16296_, _16285_);
  not (_16307_, _15915_);
  and (_16318_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_16329_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_16340_, _16329_, _16318_);
  and (_16351_, _16340_, _16307_);
  and (_16362_, _16351_, _16296_);
  and (_16372_, _16362_, _16275_);
  not (_16383_, _16372_);
  not (_16394_, _15785_);
  nor (_16405_, _15774_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_16416_, _16405_, _15861_);
  and (_16427_, _16416_, _16394_);
  not (_16438_, _16427_);
  and (_16449_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_16460_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_16470_, _16460_, _16449_);
  and (_16481_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_16492_, _15981_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_16503_, _16492_, _15697_);
  and (_16514_, _16503_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_16525_, _16514_, _16481_);
  and (_16536_, _16525_, _16470_);
  and (_16547_, _16536_, _16438_);
  not (_16557_, _16547_);
  and (_16568_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_16579_, _16568_);
  and (_16590_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_16601_, _16590_, _15915_);
  and (_16612_, _16601_, _16579_);
  nor (_16623_, _15785_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_16634_, _16623_);
  nor (_16644_, _15861_, _15796_);
  and (_16665_, _16644_, _16634_);
  and (_16666_, _16503_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_16677_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_16688_, _16677_, _16666_);
  not (_16699_, _16688_);
  nor (_16710_, _16699_, _16665_);
  and (_16721_, _16710_, _16612_);
  nor (_16732_, _16721_, _16557_);
  and (_16742_, _16732_, _16383_);
  and (_16753_, _16742_, _16209_);
  nor (_16764_, _15763_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_16775_, _16764_, _15774_);
  and (_16786_, _16775_, _15850_);
  and (_16797_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_16808_, _16797_, _16786_);
  and (_16819_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_16829_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_16840_, _16503_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_16851_, _16840_, _16829_);
  nor (_16862_, _16851_, _16819_);
  and (_16873_, _16862_, _16808_);
  not (_16884_, _16873_);
  not (_16895_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_16906_, _15850_, _16895_);
  and (_16917_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_16927_, _16917_, _16906_);
  and (_16938_, _16503_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  not (_16949_, _16938_);
  and (_16960_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_16971_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_16982_, _16971_, _16960_);
  and (_16993_, _16982_, _16949_);
  and (_17004_, _16993_, _16927_);
  and (_17015_, _16013_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_17025_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_17046_, _17025_, _15763_);
  and (_17047_, _17046_, _15850_);
  nor (_17058_, _17047_, _17015_);
  and (_17069_, _15992_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_17080_, _16503_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_17091_, _15948_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_17102_, _17091_, _17080_);
  nor (_17112_, _17102_, _17069_);
  and (_17123_, _17112_, _17058_);
  nor (_17134_, _17123_, _17004_);
  and (_17145_, _17134_, _16884_);
  and (_17156_, _17145_, _16753_);
  or (_17167_, _17156_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_17178_, ABINPUT[0]);
  nand (_17189_, _17156_, _17178_);
  and (_17200_, _17189_, _17167_);
  and (_17211_, _17200_, _15752_);
  not (_17221_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_17232_, _15741_, _17221_);
  and (_17243_, _17123_, _17004_);
  and (_17254_, _17243_, _16873_);
  and (_17265_, _17254_, _16753_);
  and (_17276_, _17265_, ABINPUT[26]);
  nor (_17287_, _17265_, _17221_);
  or (_17298_, _17287_, _17276_);
  not (_17309_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_17320_, _15741_, _17309_);
  and (_17330_, _17320_, _17298_);
  or (_17341_, _17330_, _17232_);
  or (_17352_, _17341_, _17211_);
  and (_05324_, _17352_, _39026_);
  not (_17373_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_17384_, _17265_, _17373_);
  and (_17395_, _17254_, ABINPUT[0]);
  and (_17406_, _17395_, _16753_);
  or (_17417_, _17406_, _17384_);
  and (_17428_, _17417_, _15752_);
  nor (_17439_, _15741_, _17373_);
  and (_17459_, _17265_, ABINPUT[19]);
  or (_17460_, _17459_, _17384_);
  and (_17471_, _17460_, _17320_);
  or (_17482_, _17471_, _17439_);
  or (_17493_, _17482_, _17428_);
  and (_29071_, _17493_, _39026_);
  not (_17514_, _17004_);
  and (_17525_, _17123_, _17514_);
  and (_17536_, _17525_, _16873_);
  nand (_17547_, _17536_, _16753_);
  and (_17558_, _17547_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_17568_, _17536_, ABINPUT[0]);
  and (_17579_, _17568_, _16753_);
  or (_17590_, _17579_, _17558_);
  and (_17601_, _17590_, _15752_);
  not (_17612_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_17623_, _15741_, _17612_);
  and (_17634_, _17265_, ABINPUT[20]);
  nor (_17645_, _17265_, _17612_);
  or (_17656_, _17645_, _17634_);
  and (_17667_, _17656_, _17320_);
  or (_17677_, _17667_, _17623_);
  or (_17688_, _17677_, _17601_);
  and (_29180_, _17688_, _39026_);
  nor (_17709_, _17123_, _17514_);
  and (_17720_, _17709_, _16873_);
  nand (_17731_, _17720_, _16753_);
  and (_17742_, _17731_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_17753_, _17720_, ABINPUT[0]);
  and (_17764_, _17753_, _16753_);
  or (_17775_, _17764_, _17742_);
  and (_17786_, _17775_, _15752_);
  not (_17796_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor (_17807_, _15741_, _17796_);
  and (_17818_, _17265_, ABINPUT[21]);
  nor (_17829_, _17265_, _17796_);
  or (_17840_, _17829_, _17818_);
  and (_17851_, _17840_, _17320_);
  or (_17862_, _17851_, _17807_);
  or (_17883_, _17862_, _17786_);
  and (_29289_, _17883_, _39026_);
  and (_17894_, _17134_, _16873_);
  nand (_17904_, _17894_, _16753_);
  and (_17915_, _17904_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_17926_, _17894_, ABINPUT[0]);
  and (_17937_, _17926_, _16753_);
  or (_17948_, _17937_, _17915_);
  and (_17959_, _17948_, _15752_);
  not (_17970_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_17981_, _15741_, _17970_);
  and (_17992_, _17265_, ABINPUT[22]);
  nor (_18003_, _17265_, _17970_);
  or (_18013_, _18003_, _17992_);
  and (_18024_, _18013_, _17320_);
  or (_18035_, _18024_, _17981_);
  or (_18046_, _18035_, _17959_);
  and (_29398_, _18046_, _39026_);
  and (_18067_, _17243_, _16884_);
  nand (_18078_, _18067_, _16753_);
  and (_18089_, _18078_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_18100_, _18067_, ABINPUT[0]);
  and (_18111_, _18100_, _16753_);
  or (_18122_, _18111_, _18089_);
  and (_18132_, _18122_, _15752_);
  not (_18143_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_18154_, _15741_, _18143_);
  and (_18165_, _17265_, ABINPUT[23]);
  nor (_18176_, _17265_, _18143_);
  or (_18187_, _18176_, _18165_);
  and (_18198_, _18187_, _17320_);
  or (_18209_, _18198_, _18154_);
  or (_18220_, _18209_, _18132_);
  and (_29507_, _18220_, _39026_);
  and (_18240_, _17525_, _16884_);
  nand (_18251_, _18240_, _16753_);
  and (_18262_, _18251_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_18273_, _18240_, ABINPUT[0]);
  and (_18284_, _18273_, _16753_);
  or (_18295_, _18284_, _18262_);
  and (_18306_, _18295_, _15752_);
  not (_18317_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_18338_, _15741_, _18317_);
  and (_18339_, _17265_, ABINPUT[24]);
  nor (_18350_, _17265_, _18317_);
  or (_18360_, _18350_, _18339_);
  and (_18371_, _18360_, _17320_);
  or (_18382_, _18371_, _18338_);
  or (_18393_, _18382_, _18306_);
  and (_29616_, _18393_, _39026_);
  and (_18414_, _17709_, _16884_);
  nand (_18425_, _18414_, _16753_);
  and (_18436_, _18425_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_18447_, _18414_, ABINPUT[0]);
  and (_18458_, _18447_, _16753_);
  or (_18468_, _18458_, _18436_);
  and (_18479_, _18468_, _15752_);
  not (_18490_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_18501_, _15741_, _18490_);
  and (_18512_, _17265_, ABINPUT[25]);
  nor (_18523_, _17265_, _18490_);
  or (_18534_, _18523_, _18512_);
  and (_18545_, _18534_, _17320_);
  or (_18556_, _18545_, _18501_);
  or (_18567_, _18556_, _18479_);
  and (_29725_, _18567_, _39026_);
  and (_18587_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_18598_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_18609_, _18598_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_18620_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_18631_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_18642_, _18631_, _18620_);
  and (_18653_, _18598_, _15686_);
  and (_18664_, _18653_, _18642_);
  and (_18675_, _18642_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_18686_, _18675_, _18664_);
  and (_18697_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_18707_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_18718_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_18729_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_18740_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_18751_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18762_, _18751_, _18740_);
  and (_18773_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_18784_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18795_, _18784_, _18740_);
  and (_18816_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_18817_, _18816_, _18773_);
  not (_18827_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18838_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _18827_);
  and (_18849_, _18838_, _18740_);
  and (_18860_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not (_18871_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_18882_, _18871_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_18893_, _18882_, _18740_);
  and (_18904_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_18915_, _18904_, _18860_);
  nor (_18926_, _18751_, _18740_);
  and (_18937_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_18947_, _18751_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_18958_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_18969_, _18958_, _18937_);
  and (_18980_, _18969_, _18915_);
  and (_18991_, _18980_, _18817_);
  nor (_19002_, _18991_, _18729_);
  and (_19013_, _19002_, _18718_);
  nor (_19024_, _19013_, _18707_);
  nor (_19035_, _19024_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19046_, _19035_, _18697_);
  and (_19057_, _19046_, _18664_);
  nor (_19067_, _19057_, _18686_);
  and (_19078_, _18642_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_19089_, _19078_, _18664_);
  and (_19100_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19111_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_19122_, _18729_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19133_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_19144_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_19155_, _19144_, _19133_);
  and (_19166_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_19177_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_19188_, _19177_, _19166_);
  and (_19198_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_19209_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_19220_, _19209_, _19198_);
  and (_19231_, _19220_, _19188_);
  and (_19242_, _19231_, _19155_);
  nor (_19253_, _19242_, _19122_);
  nor (_19264_, _19253_, _19111_);
  nor (_19275_, _19264_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19286_, _19275_, _19100_);
  and (_19297_, _19286_, _18664_);
  nor (_19318_, _19297_, _19089_);
  not (_19319_, _19318_);
  nor (_19341_, _19319_, _19067_);
  and (_19342_, _18642_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_19364_, _19342_, _18664_);
  not (_19365_, _18664_);
  and (_19387_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_19388_, _19387_);
  and (_19399_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_19410_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_19421_, _19410_, _19399_);
  and (_19432_, _19421_, _19388_);
  and (_19443_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_19453_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_19464_, _19453_, _19443_);
  and (_19475_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_19486_, _19475_, _18729_);
  and (_19497_, _19486_, _19464_);
  and (_19508_, _19497_, _19432_);
  and (_19519_, _19508_, _18718_);
  nor (_19530_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _18718_);
  nor (_19541_, _19530_, _19519_);
  nor (_19552_, _19541_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_19563_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_19574_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _19563_);
  nor (_19584_, _19574_, _19552_);
  nor (_19595_, _19584_, _19365_);
  nor (_19606_, _19595_, _19364_);
  and (_19617_, _19606_, _19341_);
  and (_19628_, _18642_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_19639_, _19628_, _18664_);
  and (_19650_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19661_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19672_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_19682_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_19693_, _19682_, _19672_);
  and (_19704_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_19715_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_19726_, _19715_, _19704_);
  and (_19737_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_19748_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_19759_, _19748_, _19737_);
  and (_19770_, _19759_, _19726_);
  and (_19781_, _19770_, _19693_);
  nor (_19792_, _19781_, _18729_);
  and (_19802_, _19792_, _18718_);
  or (_19813_, _19802_, _19661_);
  and (_19824_, _19813_, _19563_);
  nor (_19835_, _19824_, _19650_);
  and (_19846_, _19835_, _18664_);
  nor (_19857_, _19846_, _19639_);
  not (_19868_, _19857_);
  and (_19879_, _18642_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_19890_, _19879_, _18664_);
  and (_19901_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19911_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19922_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_19933_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_19944_, _19933_, _19922_);
  and (_19955_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_19966_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_19977_, _19966_, _19955_);
  and (_19988_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_19999_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_20010_, _19999_, _19988_);
  and (_20020_, _20010_, _19977_);
  and (_20031_, _20020_, _19944_);
  nor (_20042_, _20031_, _19122_);
  or (_20053_, _20042_, _19911_);
  and (_20064_, _20053_, _19563_);
  nor (_20075_, _20064_, _19901_);
  and (_20086_, _20075_, _18664_);
  nor (_20097_, _20086_, _19890_);
  and (_20108_, _18642_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_20119_, _20108_, _18664_);
  and (_20129_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_20140_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_20151_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_20162_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_20173_, _20162_, _20151_);
  and (_20184_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_20195_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_20206_, _20195_, _20184_);
  and (_20217_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_20228_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_20238_, _20228_, _20217_);
  and (_20249_, _20238_, _20206_);
  and (_20260_, _20249_, _20173_);
  nor (_20271_, _20260_, _19122_);
  nor (_20282_, _20271_, _20140_);
  nor (_20293_, _20282_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_20304_, _20293_, _20129_);
  and (_20315_, _20304_, _18664_);
  nor (_20326_, _20315_, _20119_);
  nor (_20337_, _20326_, _20097_);
  and (_20347_, _20337_, _19868_);
  and (_20358_, _20347_, _19617_);
  and (_20369_, _19606_, _19318_);
  and (_20380_, _18642_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_20391_, _20380_, _18664_);
  and (_20402_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_20413_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_20424_, _20413_, _20402_);
  and (_20435_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_20446_, _20435_, _18729_);
  and (_20456_, _20446_, _20424_);
  and (_20467_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_20478_, _20467_);
  and (_20489_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_20500_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_20511_, _20500_, _20489_);
  and (_20522_, _20511_, _20478_);
  and (_20533_, _20522_, _20456_);
  and (_20544_, _20533_, _18718_);
  nor (_20555_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _18718_);
  nor (_20565_, _20555_, _20544_);
  nor (_20576_, _20565_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_20587_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _19563_);
  nor (_20598_, _20587_, _20576_);
  nor (_20609_, _20598_, _19365_);
  nor (_20620_, _20609_, _20391_);
  not (_20631_, _20620_);
  nor (_20642_, _20631_, _19067_);
  and (_20653_, _20642_, _20369_);
  not (_20664_, _20326_);
  nor (_20674_, _20664_, _20097_);
  and (_20685_, _20674_, _19857_);
  and (_20696_, _20685_, _20653_);
  or (_20707_, _20696_, _20358_);
  and (_20718_, _20326_, _20097_);
  and (_20729_, _20718_, _19868_);
  and (_20740_, _20729_, _19617_);
  and (_20751_, _20674_, _19868_);
  and (_20762_, _20751_, _20620_);
  and (_20773_, _20762_, _19617_);
  or (_20784_, _20773_, _20740_);
  or (_20794_, _20784_, _20707_);
  and (_20805_, _20097_, _19868_);
  and (_20816_, _20805_, _20664_);
  and (_20827_, _20816_, _20653_);
  and (_20838_, _20337_, _19857_);
  and (_20849_, _20838_, _19617_);
  or (_20860_, _20849_, _20827_);
  or (_20871_, _19318_, _19067_);
  and (_20882_, _18642_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_20893_, _20882_, _18664_);
  and (_20903_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20914_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20925_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_20936_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_20947_, _20936_, _20925_);
  and (_20958_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_20969_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_20980_, _20969_, _20958_);
  and (_20991_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_21002_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_21012_, _21002_, _20991_);
  and (_21023_, _21012_, _20980_);
  and (_21034_, _21023_, _20947_);
  nor (_21045_, _21034_, _18729_);
  and (_21056_, _21045_, _18718_);
  or (_21067_, _21056_, _20914_);
  and (_21078_, _21067_, _19563_);
  nor (_21089_, _21078_, _20903_);
  and (_21100_, _21089_, _18664_);
  nor (_21111_, _21100_, _20893_);
  or (_21121_, _21111_, _19606_);
  nor (_21132_, _21121_, _20871_);
  and (_21143_, _20729_, _20620_);
  and (_21154_, _21143_, _21132_);
  and (_21165_, _20751_, _20631_);
  and (_21176_, _21165_, _19617_);
  or (_21187_, _21176_, _21154_);
  or (_21198_, _21187_, _20860_);
  nor (_21209_, _21198_, _20794_);
  not (_21220_, _19606_);
  nor (_21230_, _20871_, _21220_);
  and (_21241_, _21230_, _21111_);
  and (_21252_, _20631_, _19857_);
  and (_21263_, _21252_, _20674_);
  and (_21274_, _21263_, _21241_);
  not (_21285_, _21274_);
  and (_21296_, _21241_, _20762_);
  and (_21307_, _20097_, _19857_);
  and (_21318_, _21307_, _20664_);
  and (_21329_, _21318_, _20620_);
  and (_21339_, _21329_, _21241_);
  nor (_21350_, _21339_, _21296_);
  and (_21361_, _21350_, _21285_);
  and (_21372_, _20631_, _19617_);
  and (_21383_, _21307_, _20326_);
  nor (_21394_, _21383_, _20816_);
  not (_21405_, _21394_);
  and (_21416_, _21405_, _21372_);
  not (_21427_, _21416_);
  not (_21438_, _21111_);
  and (_21448_, _21230_, _21438_);
  and (_21459_, _21448_, _20838_);
  and (_21470_, _21318_, _21372_);
  nor (_21481_, _21470_, _21459_);
  and (_21492_, _21481_, _21427_);
  and (_21503_, _21492_, _21361_);
  and (_21514_, _21503_, _21209_);
  nor (_21525_, _21514_, _18609_);
  not (_21536_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_21547_, \oc8051_top_1.oc8051_decoder1.state [1], _15686_);
  and (_21557_, _21547_, _21536_);
  and (_21568_, _21557_, _21318_);
  and (_21579_, _21568_, _21132_);
  and (_21590_, _21459_, _21547_);
  and (_21601_, _21590_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_21612_, _21601_, _21579_);
  nor (_21623_, _21612_, _21525_);
  nor (_21634_, _21623_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_21645_, _21634_, _18587_);
  and (_21656_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_21667_, _21252_, _20337_);
  and (_21677_, _21667_, _21132_);
  not (_21688_, _21677_);
  and (_21699_, _20620_, _19857_);
  and (_21710_, _21699_, _20337_);
  and (_21721_, _21710_, _21132_);
  and (_21732_, _20620_, _20347_);
  and (_21743_, _21732_, _21132_);
  nor (_21754_, _21743_, _21721_);
  and (_21765_, _21754_, _21688_);
  and (_21776_, _21220_, _19341_);
  and (_21786_, _21776_, _21111_);
  and (_21797_, _21252_, _20718_);
  and (_21808_, _21797_, _21786_);
  and (_21819_, _21699_, _20674_);
  and (_21830_, _21786_, _21819_);
  nor (_21841_, _21830_, _21808_);
  and (_21852_, _21841_, _21765_);
  and (_21863_, _21448_, _21165_);
  and (_21874_, _20816_, _20620_);
  and (_21885_, _21230_, _21874_);
  nor (_21895_, _21885_, _21863_);
  not (_21906_, _21895_);
  nor (_21917_, _21874_, _20838_);
  not (_21928_, _21786_);
  nor (_21939_, _21928_, _21917_);
  nor (_21950_, _21939_, _21906_);
  and (_21961_, _20631_, _20347_);
  and (_21972_, _21961_, _21786_);
  and (_21983_, _21263_, _19617_);
  nor (_21994_, _21983_, _21972_);
  and (_22005_, _21994_, _21950_);
  and (_22016_, _22005_, _21852_);
  and (_22027_, _21263_, _21132_);
  and (_22038_, _20816_, _20631_);
  and (_22049_, _22038_, _21786_);
  nor (_22060_, _22049_, _22027_);
  and (_22071_, _22038_, _21241_);
  and (_22082_, _22038_, _21448_);
  nor (_22093_, _22082_, _22071_);
  and (_22104_, _22093_, _22060_);
  and (_22115_, _21448_, _21819_);
  and (_22126_, _20729_, _20631_);
  and (_22137_, _22126_, _21448_);
  nor (_22148_, _22137_, _22115_);
  and (_22159_, _21786_, _21143_);
  and (_22170_, _21786_, _21732_);
  nor (_22181_, _22170_, _22159_);
  and (_22192_, _22181_, _22148_);
  and (_22203_, _21448_, _21329_);
  and (_22214_, _21132_, _21819_);
  nor (_22225_, _22214_, _22203_);
  and (_22236_, _22225_, _22192_);
  and (_22247_, _22236_, _22104_);
  and (_22258_, _21132_, _20729_);
  not (_22269_, _22258_);
  and (_22280_, _21318_, _20631_);
  and (_22291_, _22280_, _21241_);
  and (_22302_, _22280_, _21448_);
  nor (_22313_, _22302_, _22291_);
  and (_22324_, _22313_, _22269_);
  and (_22335_, _21448_, _21143_);
  and (_22346_, _21448_, _21263_);
  nor (_22357_, _22346_, _22335_);
  and (_22368_, _20631_, _19067_);
  and (_22379_, _22368_, _20685_);
  nor (_22390_, _22379_, _21459_);
  and (_22401_, _21786_, _20762_);
  not (_22412_, _22401_);
  and (_22423_, _22412_, _22390_);
  and (_22434_, _22423_, _22357_);
  and (_22445_, _21448_, _20762_);
  and (_22456_, _21786_, _21165_);
  nor (_22467_, _22456_, _22445_);
  and (_22478_, _21786_, _22280_);
  and (_22489_, _22126_, _21786_);
  nor (_22500_, _22489_, _22478_);
  and (_22511_, _22500_, _22467_);
  and (_22522_, _22511_, _22434_);
  and (_22533_, _22522_, _22324_);
  and (_22544_, _22533_, _22247_);
  and (_22555_, _22544_, _22016_);
  nor (_22566_, _22555_, _18609_);
  and (_22577_, _21132_, _20838_);
  and (_22588_, _22577_, _20631_);
  or (_22599_, _21743_, _22588_);
  and (_22610_, _22599_, _21557_);
  and (_22621_, _20664_, _20097_);
  and (_22632_, _21132_, _22621_);
  and (_22643_, _22632_, _21557_);
  or (_22654_, _22643_, _21601_);
  or (_22665_, _22654_, _22610_);
  nor (_22676_, _22665_, _22566_);
  nor (_22687_, _22676_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22698_, _22687_, _21656_);
  nor (_22709_, _22698_, _21645_);
  and (_22720_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_22731_, _18609_);
  and (_22742_, _21776_, _21438_);
  and (_22753_, _22742_, _21165_);
  and (_22764_, _22742_, _21263_);
  nor (_22775_, _22764_, _22753_);
  nor (_22786_, _22775_, _22731_);
  and (_22797_, _22775_, _21361_);
  nor (_22808_, _22797_, _18609_);
  or (_22819_, _22808_, _22643_);
  nor (_22830_, _22819_, _22786_);
  nor (_22841_, _22830_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22852_, _22841_, _22720_);
  and (_22863_, _22852_, _39026_);
  and (_35268_, _22863_, _22709_);
  not (_22884_, _17320_);
  and (_22895_, _16383_, _16198_);
  and (_22906_, _16721_, _16057_);
  and (_22917_, _22906_, _22895_);
  and (_22928_, _22917_, _16547_);
  nand (_22939_, _22928_, _17536_);
  nor (_22950_, _22939_, _22884_);
  and (_22961_, _22950_, ABINPUT[10]);
  nor (_22972_, _22950_, _16220_);
  nor (_22983_, _22972_, _22961_);
  not (_22994_, _22983_);
  not (_23005_, _22950_);
  and (_23016_, _23005_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_23027_, _22950_, ABINPUT[9]);
  nor (_23038_, _23027_, _23016_);
  and (_23049_, _23005_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_23060_, _22950_, ABINPUT[8]);
  nor (_23071_, _23060_, _23049_);
  and (_23082_, _23005_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_23093_, _22950_, ABINPUT[7]);
  nor (_23104_, _23093_, _23082_);
  and (_23115_, _23005_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_23126_, _22950_, ABINPUT[6]);
  nor (_23137_, _23126_, _23115_);
  and (_23148_, _23005_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_23159_, _22950_, ABINPUT[5]);
  nor (_23170_, _23159_, _23148_);
  and (_23181_, _23005_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_23192_, _22950_, ABINPUT[4]);
  nor (_23203_, _23192_, _23181_);
  nor (_23214_, _22950_, _16895_);
  and (_23225_, _22950_, ABINPUT[3]);
  nor (_23236_, _23225_, _23214_);
  and (_23247_, _23236_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_23258_, _23247_, _23203_);
  and (_23269_, _23258_, _23170_);
  and (_23280_, _23269_, _23137_);
  and (_23291_, _23280_, _23104_);
  and (_23302_, _23291_, _23071_);
  and (_23313_, _23302_, _23038_);
  and (_23324_, _23313_, _22994_);
  nor (_23335_, _23313_, _22994_);
  nor (_23346_, _23335_, _23324_);
  and (_23357_, _23346_, _15861_);
  nor (_23367_, _23357_, _16264_);
  nor (_23378_, _23367_, _22950_);
  nor (_23389_, _23378_, _22961_);
  nor (_35488_, _23389_, rst);
  not (_23410_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_23421_, _23236_, _23410_);
  nor (_23432_, _23236_, _23410_);
  nor (_23443_, _23432_, _23421_);
  and (_23454_, _23443_, _15861_);
  nor (_23465_, _23454_, _16906_);
  nor (_23475_, _23465_, _22950_);
  nor (_23486_, _23475_, _23225_);
  nand (_38077_, _23486_, _39026_);
  nor (_23507_, _23247_, _23203_);
  nor (_23518_, _23507_, _23258_);
  nor (_23529_, _23518_, _15850_);
  nor (_23540_, _23529_, _17047_);
  nor (_23551_, _23540_, _22950_);
  nor (_23562_, _23551_, _23192_);
  nand (_38086_, _23562_, _39026_);
  nor (_23583_, _23258_, _23170_);
  nor (_23594_, _23583_, _23269_);
  nor (_23605_, _23594_, _15850_);
  nor (_23616_, _23605_, _16786_);
  nor (_23627_, _23616_, _22950_);
  nor (_23638_, _23627_, _23159_);
  nand (_38094_, _23638_, _39026_);
  nor (_23659_, _23269_, _23137_);
  nor (_23670_, _23659_, _23280_);
  nor (_23681_, _23670_, _15850_);
  nor (_23692_, _23681_, _16427_);
  nor (_23702_, _23692_, _22950_);
  nor (_23713_, _23702_, _23126_);
  nor (_38103_, _23713_, rst);
  nor (_23734_, _23280_, _23104_);
  nor (_23745_, _23734_, _23291_);
  nor (_23756_, _23745_, _15850_);
  nor (_23767_, _23756_, _16665_);
  nor (_23778_, _23767_, _22950_);
  nor (_23789_, _23778_, _23093_);
  nor (_38111_, _23789_, rst);
  nor (_23810_, _23291_, _23071_);
  nor (_23820_, _23810_, _23302_);
  nor (_23831_, _23820_, _15850_);
  nor (_23842_, _23831_, _15894_);
  nor (_23853_, _23842_, _22950_);
  nor (_23864_, _23853_, _23060_);
  nor (_38119_, _23864_, rst);
  nor (_23885_, _23302_, _23038_);
  nor (_23896_, _23885_, _23313_);
  nor (_23907_, _23896_, _15850_);
  nor (_23918_, _23907_, _16111_);
  nor (_23928_, _23918_, _22950_);
  nor (_23939_, _23928_, _23027_);
  nor (_38128_, _23939_, rst);
  and (_23960_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15686_);
  and (_23971_, _23960_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_23982_, _17894_, _16547_);
  nand (_23993_, _23982_, _22917_);
  nor (_24004_, _23993_, _22884_);
  or (_24015_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_24026_, ABINPUT[26]);
  nand (_24037_, _24004_, _24026_);
  and (_24047_, _24037_, _24015_);
  or (_24058_, _24047_, _23971_);
  not (_24069_, ABINPUT[18]);
  nand (_24080_, _23971_, _24069_);
  and (_24091_, _24080_, _39026_);
  and (_40187_, _24091_, _24058_);
  and (_24112_, _22928_, _17720_);
  and (_24123_, _24112_, _17320_);
  nor (_24134_, _24123_, _23971_);
  and (_24145_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_24156_, _24134_, _24026_);
  or (_24167_, _24156_, _24145_);
  and (_40208_, _24167_, _39026_);
  or (_24188_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_24199_, ABINPUT[19]);
  nand (_24210_, _24004_, _24199_);
  and (_24220_, _24210_, _24188_);
  or (_24231_, _24220_, _23971_);
  not (_24242_, ABINPUT[11]);
  nand (_24253_, _23971_, _24242_);
  and (_24264_, _24253_, _39026_);
  and (_41219_, _24264_, _24231_);
  or (_24285_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_24295_, ABINPUT[20]);
  nand (_24306_, _24004_, _24295_);
  and (_24317_, _24306_, _24285_);
  or (_24328_, _24317_, _23971_);
  not (_24339_, ABINPUT[12]);
  nand (_24350_, _23971_, _24339_);
  and (_24361_, _24350_, _39026_);
  and (_41228_, _24361_, _24328_);
  or (_24381_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_24392_, ABINPUT[21]);
  nand (_24403_, _24004_, _24392_);
  and (_24414_, _24403_, _24381_);
  or (_24425_, _24414_, _23971_);
  not (_24436_, ABINPUT[13]);
  nand (_24447_, _23971_, _24436_);
  and (_24458_, _24447_, _39026_);
  and (_41236_, _24458_, _24425_);
  or (_24478_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_24489_, ABINPUT[22]);
  nand (_24500_, _24004_, _24489_);
  and (_24511_, _24500_, _24478_);
  or (_24522_, _24511_, _23971_);
  not (_24533_, ABINPUT[14]);
  nand (_24544_, _23971_, _24533_);
  and (_24554_, _24544_, _39026_);
  and (_41245_, _24554_, _24522_);
  or (_24575_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_24586_, ABINPUT[23]);
  nand (_24597_, _24004_, _24586_);
  and (_24608_, _24597_, _24575_);
  or (_24619_, _24608_, _23971_);
  not (_24630_, ABINPUT[15]);
  nand (_24640_, _23971_, _24630_);
  and (_24651_, _24640_, _39026_);
  and (_41254_, _24651_, _24619_);
  or (_24672_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_24683_, ABINPUT[24]);
  nand (_24694_, _24004_, _24683_);
  and (_24705_, _24694_, _24672_);
  or (_24716_, _24705_, _23971_);
  not (_24726_, ABINPUT[16]);
  nand (_24737_, _23971_, _24726_);
  and (_24748_, _24737_, _39026_);
  and (_41263_, _24748_, _24716_);
  or (_24769_, _24004_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_24780_, ABINPUT[25]);
  nand (_24791_, _24004_, _24780_);
  and (_24802_, _24791_, _24769_);
  or (_24812_, _24802_, _23971_);
  not (_24823_, ABINPUT[17]);
  nand (_24834_, _23971_, _24823_);
  and (_24845_, _24834_, _39026_);
  and (_41272_, _24845_, _24812_);
  and (_24866_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_24877_, _24134_, _24199_);
  or (_24888_, _24877_, _24866_);
  and (_41280_, _24888_, _39026_);
  and (_24908_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_24919_, _24134_, _24295_);
  or (_24930_, _24919_, _24908_);
  and (_41289_, _24930_, _39026_);
  and (_24951_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nor (_24962_, _24134_, _24392_);
  or (_24973_, _24962_, _24951_);
  and (_41297_, _24973_, _39026_);
  and (_24993_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_25004_, _24134_, _24489_);
  or (_25015_, _25004_, _24993_);
  and (_41306_, _25015_, _39026_);
  and (_25036_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_25047_, _24134_, _24586_);
  or (_25058_, _25047_, _25036_);
  and (_41314_, _25058_, _39026_);
  and (_25078_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_25089_, _24134_, _24683_);
  or (_25100_, _25089_, _25078_);
  and (_41323_, _25100_, _39026_);
  and (_25121_, _24134_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_25132_, _24134_, _24780_);
  or (_25143_, _25132_, _25121_);
  and (_41331_, _25143_, _39026_);
  nor (_25163_, _16372_, _16198_);
  and (_25174_, _16732_, _16057_);
  and (_25185_, _25174_, _25163_);
  and (_25196_, _25185_, _15752_);
  and (_25207_, _17145_, ABINPUT[0]);
  not (_25218_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25229_, _17145_, _25218_);
  nor (_25239_, _25229_, _25207_);
  nand (_25250_, _25239_, _25196_);
  nor (_25261_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_25272_, _25261_, ABINPUT[0]);
  nand (_25283_, _25261_, _25218_);
  and (_25294_, _25283_, _25272_);
  or (_25305_, _25294_, _25196_);
  and (_25316_, _25305_, _25250_);
  and (_25326_, _17320_, _17254_);
  and (_25337_, _25326_, _25185_);
  not (_25348_, _25337_);
  and (_25359_, _25348_, _25316_);
  and (_25370_, _25337_, ABINPUT[10]);
  or (_25381_, _25370_, _25359_);
  and (_01572_, _25381_, _39026_);
  nand (_25402_, _25196_, _17536_);
  and (_25413_, _25402_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_25423_, _25196_, _17568_);
  or (_25434_, _25423_, _25337_);
  or (_25445_, _25434_, _25413_);
  not (_25456_, ABINPUT[4]);
  nand (_25467_, _25337_, _25456_);
  and (_25478_, _25467_, _25445_);
  and (_06388_, _25478_, _39026_);
  not (_25499_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_25510_, _17720_, _25499_);
  nor (_25520_, _25510_, _17753_);
  nand (_25531_, _25520_, _25196_);
  and (_25542_, ABINPUT[2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_25553_, _25499_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_25564_, _25553_, _25542_);
  or (_25575_, _25564_, _25196_);
  and (_25586_, _25575_, _25531_);
  and (_25597_, _25586_, _25348_);
  and (_25608_, _25337_, ABINPUT[5]);
  or (_25619_, _25608_, _25597_);
  and (_06399_, _25619_, _39026_);
  nand (_25639_, _25196_, _17894_);
  and (_25650_, _25639_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_25661_, _25196_, _17926_);
  or (_25672_, _25661_, _25650_);
  and (_25683_, _25672_, _25348_);
  and (_25694_, _25337_, ABINPUT[6]);
  or (_25705_, _25694_, _25683_);
  and (_06410_, _25705_, _39026_);
  nand (_25726_, _25196_, _18067_);
  and (_25737_, _25726_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_25747_, _25196_, _18100_);
  or (_25758_, _25747_, _25737_);
  and (_25769_, _25758_, _25348_);
  and (_25780_, _25337_, ABINPUT[7]);
  or (_25791_, _25780_, _25769_);
  and (_06421_, _25791_, _39026_);
  nand (_25812_, _25196_, _18240_);
  and (_25823_, _25812_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_25834_, _25196_, _18273_);
  or (_25845_, _25834_, _25337_);
  or (_25856_, _25845_, _25823_);
  not (_25866_, ABINPUT[8]);
  nand (_25877_, _25337_, _25866_);
  and (_25888_, _25877_, _25856_);
  and (_06432_, _25888_, _39026_);
  not (_25909_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_25920_, _18414_, _25909_);
  nor (_25931_, _25920_, _18447_);
  nand (_25942_, _25931_, _25196_);
  and (_25953_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_25964_, _25953_, ABINPUT[1]);
  nor (_25975_, _25953_, _25909_);
  or (_25985_, _25975_, _25964_);
  or (_25996_, _25985_, _25196_);
  and (_26007_, _25996_, _25942_);
  and (_26018_, _26007_, _25348_);
  and (_26029_, _25337_, ABINPUT[9]);
  or (_26040_, _26029_, _26018_);
  and (_06443_, _26040_, _39026_);
  not (_26061_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_26072_, _23960_, _26061_);
  and (_26083_, _26072_, ABINPUT[18]);
  nor (_26093_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26104_, _26093_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_26115_, _17254_, _16547_);
  not (_26126_, _16057_);
  and (_26137_, _16721_, _26126_);
  and (_26148_, _26137_, _25163_);
  and (_26159_, _26148_, _26115_);
  and (_26170_, _26159_, _17320_);
  nor (_26181_, _26170_, _26104_);
  nor (_26192_, _26181_, _24026_);
  not (_26203_, _26181_);
  and (_26213_, _16721_, _16547_);
  not (_26224_, _15752_);
  nor (_26235_, _26224_, _16372_);
  and (_26246_, _26235_, _16209_);
  and (_26257_, _26246_, _26213_);
  nand (_26268_, _26257_, _17145_);
  and (_26279_, _26268_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_26290_, _26213_, _16209_);
  and (_26300_, _26235_, _26290_);
  and (_26311_, _26300_, _25207_);
  nor (_26322_, _26311_, _26279_);
  nor (_26333_, _26322_, _26203_);
  nor (_26344_, _26333_, _26192_);
  nor (_26355_, _26344_, _26072_);
  nor (_26366_, _26355_, _26083_);
  nor (_07163_, _26366_, rst);
  and (_26387_, _26072_, ABINPUT[11]);
  or (_26398_, _26072_, _24199_);
  nor (_26408_, _26398_, _26181_);
  nor (_26419_, _26408_, _26387_);
  not (_26430_, _26072_);
  and (_26441_, _26181_, _26430_);
  not (_26452_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_26463_, _26300_, _17254_);
  nor (_26474_, _26463_, _26452_);
  and (_26485_, _26257_, _17395_);
  nor (_26496_, _26485_, _26474_);
  not (_26507_, _26496_);
  and (_26518_, _26507_, _26441_);
  not (_26528_, _26518_);
  and (_26539_, _26528_, _26419_);
  nor (_08869_, _26539_, rst);
  and (_26560_, _26072_, ABINPUT[12]);
  nor (_26571_, _26181_, _24295_);
  nand (_26582_, _26257_, _17536_);
  and (_26593_, _26582_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_26604_, _26300_, _17568_);
  nor (_26615_, _26604_, _26593_);
  nor (_26626_, _26615_, _26203_);
  nor (_26637_, _26626_, _26571_);
  nor (_26647_, _26637_, _26072_);
  nor (_26658_, _26647_, _26560_);
  nor (_08880_, _26658_, rst);
  and (_26679_, _26072_, ABINPUT[13]);
  not (_26690_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_26701_, _26300_, _17720_);
  nor (_26712_, _26701_, _26690_);
  and (_26723_, _26300_, _17753_);
  nor (_26734_, _26723_, _26712_);
  and (_26745_, _26734_, _26181_);
  nor (_26756_, _26181_, ABINPUT[21]);
  or (_26767_, _26756_, _26745_);
  nor (_26778_, _26767_, _26072_);
  nor (_26788_, _26778_, _26679_);
  nor (_08891_, _26788_, rst);
  and (_26809_, _26072_, _24533_);
  and (_26820_, _26441_, _26257_);
  and (_26831_, _26820_, _17926_);
  not (_26842_, _26831_);
  nand (_26853_, _26257_, _17894_);
  and (_26864_, _26853_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_26875_, _26864_, _26441_);
  nor (_26886_, _26181_, _24489_);
  nor (_26897_, _26886_, _26875_);
  and (_26908_, _26897_, _26842_);
  and (_26918_, _26908_, _26430_);
  nor (_26929_, _26918_, _26809_);
  and (_08902_, _26929_, _39026_);
  and (_26950_, _26072_, _24630_);
  nor (_26961_, _26181_, _24586_);
  or (_26972_, _26961_, _26072_);
  not (_26983_, _26972_);
  not (_26994_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_27005_, _26300_, _18067_);
  nor (_27016_, _27005_, _26994_);
  and (_27027_, _27016_, _26441_);
  and (_27038_, _26820_, _18100_);
  nor (_27048_, _27038_, _27027_);
  and (_27059_, _27048_, _26983_);
  nor (_27070_, _27059_, _26950_);
  and (_08913_, _27070_, _39026_);
  and (_27091_, _26072_, ABINPUT[16]);
  nor (_27102_, _26072_, _24683_);
  or (_27113_, _27102_, _26441_);
  not (_27124_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_27135_, _18240_, _27124_);
  or (_27146_, _27135_, _18273_);
  and (_27156_, _27146_, _26820_);
  not (_27167_, _26300_);
  nand (_27178_, _27167_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_27189_, _27178_, _26181_);
  or (_27200_, _27189_, _27156_);
  and (_27211_, _27200_, _27113_);
  or (_27222_, _27211_, _27091_);
  and (_08924_, _27222_, _39026_);
  and (_27243_, _26072_, _24823_);
  and (_27254_, _26820_, _18447_);
  not (_27264_, _27254_);
  not (_27275_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_27286_, _26300_, _18414_);
  nor (_27297_, _27286_, _27275_);
  and (_27308_, _27297_, _26441_);
  nor (_27319_, _26181_, _24780_);
  nor (_27330_, _27319_, _27308_);
  and (_27341_, _27330_, _27264_);
  and (_27352_, _27341_, _26430_);
  nor (_27363_, _27352_, _27243_);
  and (_08935_, _27363_, _39026_);
  and (_27383_, _22928_, _17145_);
  or (_27394_, _27383_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand (_27405_, _27383_, _17178_);
  and (_27416_, _27405_, _15752_);
  and (_27427_, _27416_, _27394_);
  not (_27438_, ABINPUT[10]);
  and (_27449_, _22917_, _26115_);
  nand (_27460_, _27449_, _27438_);
  or (_27471_, _27449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_27482_, _27471_, _17320_);
  and (_27492_, _27482_, _27460_);
  not (_27503_, _15741_);
  and (_27514_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_27525_, _27514_, rst);
  or (_27536_, _27525_, _27492_);
  or (_19308_, _27536_, _27427_);
  and (_27557_, _25174_, _22895_);
  nand (_27568_, _27557_, _17145_);
  and (_27579_, _27568_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_27590_, _27557_, _25207_);
  or (_27601_, _27590_, _27579_);
  and (_27611_, _27601_, _15752_);
  and (_27622_, _27557_, _17254_);
  and (_27633_, _27622_, ABINPUT[10]);
  not (_27644_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_27655_, _27622_, _27644_);
  or (_27666_, _27655_, _27633_);
  and (_27677_, _27666_, _17320_);
  nor (_27688_, _15741_, _27644_);
  or (_27699_, _27688_, rst);
  or (_27710_, _27699_, _27677_);
  or (_19330_, _27710_, _27611_);
  and (_27730_, _26137_, _22895_);
  and (_27741_, _27730_, _26115_);
  and (_27752_, _27741_, ABINPUT[10]);
  not (_27763_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_27774_, _27741_, _27763_);
  or (_27785_, _27774_, _27752_);
  and (_27796_, _27785_, _17320_);
  and (_27807_, _27730_, _16547_);
  nor (_27818_, _17145_, _27763_);
  or (_27829_, _27818_, _25207_);
  and (_27839_, _27829_, _27807_);
  nor (_27850_, _27807_, _27763_);
  or (_27861_, _27850_, _27839_);
  and (_27872_, _27861_, _15752_);
  nor (_27883_, _15741_, _27763_);
  or (_27894_, _27883_, rst);
  or (_27905_, _27894_, _27872_);
  or (_19353_, _27905_, _27796_);
  nor (_27925_, _16721_, _16057_);
  and (_27936_, _22895_, _27925_);
  and (_27947_, _27936_, _26115_);
  and (_27958_, _27947_, ABINPUT[10]);
  not (_27969_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_27980_, _27947_, _27969_);
  or (_27991_, _27980_, _27958_);
  and (_28001_, _27991_, _17320_);
  nor (_28012_, _17145_, _27969_);
  or (_28023_, _28012_, _25207_);
  and (_28034_, _16198_, _26126_);
  and (_28045_, _28034_, _16742_);
  and (_28056_, _28045_, _28023_);
  nor (_28067_, _28045_, _27969_);
  or (_28078_, _28067_, _28056_);
  and (_28089_, _28078_, _15752_);
  nor (_28099_, _15741_, _27969_);
  or (_28110_, _28099_, rst);
  or (_28121_, _28110_, _28089_);
  or (_19376_, _28121_, _28001_);
  not (_28142_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_28153_, _27449_, _28142_);
  and (_28164_, _22928_, _17395_);
  or (_28175_, _28164_, _28153_);
  and (_28185_, _28175_, _15752_);
  and (_28196_, _27449_, ABINPUT[3]);
  or (_28207_, _28196_, _28153_);
  and (_28218_, _28207_, _17320_);
  nor (_28229_, _15741_, _28142_);
  or (_28240_, _28229_, rst);
  or (_28251_, _28240_, _28218_);
  or (_38290_, _28251_, _28185_);
  nand (_28271_, _27449_, _25456_);
  or (_28282_, _27449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_28293_, _28282_, _17320_);
  and (_28304_, _28293_, _28271_);
  and (_28315_, _22928_, _17568_);
  and (_28326_, _22939_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_28337_, _28326_, _28315_);
  and (_28348_, _28337_, _15752_);
  and (_28358_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_28369_, _28358_, rst);
  or (_28380_, _28369_, _28348_);
  or (_38292_, _28380_, _28304_);
  not (_28401_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_28412_, _24112_, _28401_);
  and (_28423_, _22928_, _17753_);
  or (_28434_, _28423_, _28412_);
  and (_28444_, _28434_, _15752_);
  nor (_28455_, _27449_, _28401_);
  and (_28466_, _27449_, ABINPUT[5]);
  or (_28477_, _28466_, _28455_);
  and (_28488_, _28477_, _17320_);
  nor (_28499_, _15741_, _28401_);
  or (_28510_, _28499_, rst);
  or (_28521_, _28510_, _28488_);
  or (_38294_, _28521_, _28444_);
  not (_28541_, ABINPUT[6]);
  nand (_28552_, _27449_, _28541_);
  or (_28563_, _27449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_28574_, _28563_, _17320_);
  and (_28585_, _28574_, _28552_);
  and (_28596_, _23993_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_28607_, _22928_, _17926_);
  or (_28617_, _28607_, _28596_);
  and (_28628_, _28617_, _15752_);
  and (_28639_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_28650_, _28639_, rst);
  or (_28661_, _28650_, _28628_);
  or (_38296_, _28661_, _28585_);
  and (_28682_, _22928_, _18067_);
  or (_28693_, _28682_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_28703_, _28682_, _17178_);
  and (_28714_, _28703_, _15752_);
  and (_28725_, _28714_, _28693_);
  not (_28736_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_28747_, _27449_, _28736_);
  and (_28758_, _27449_, ABINPUT[7]);
  or (_28769_, _28758_, _28747_);
  and (_28780_, _28769_, _17320_);
  nor (_28790_, _15741_, _28736_);
  or (_28801_, _28790_, rst);
  or (_28812_, _28801_, _28780_);
  or (_38298_, _28812_, _28725_);
  nand (_28833_, _22928_, _18240_);
  and (_28844_, _28833_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_28855_, _22928_, _18273_);
  or (_28866_, _28855_, _28844_);
  and (_28876_, _28866_, _15752_);
  not (_28887_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_28898_, _27449_, _28887_);
  and (_28909_, _27449_, ABINPUT[8]);
  or (_28920_, _28909_, _28898_);
  and (_28931_, _28920_, _17320_);
  nor (_28942_, _15741_, _28887_);
  or (_28953_, _28942_, rst);
  or (_28963_, _28953_, _28931_);
  or (_38300_, _28963_, _28876_);
  nand (_28984_, _22928_, _18414_);
  and (_28995_, _28984_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_29006_, _22928_, _18447_);
  or (_29017_, _29006_, _28995_);
  and (_29028_, _29017_, _15752_);
  not (_29039_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_29049_, _27449_, _29039_);
  and (_29060_, _27449_, ABINPUT[9]);
  or (_29072_, _29060_, _29049_);
  and (_29083_, _29072_, _17320_);
  nor (_29094_, _15741_, _29039_);
  or (_29105_, _29094_, rst);
  or (_29116_, _29105_, _29083_);
  or (_38302_, _29116_, _29028_);
  and (_29136_, _15752_, ABINPUT[0]);
  and (_29147_, _17320_, ABINPUT[3]);
  or (_29158_, _29147_, _29136_);
  and (_29169_, _29158_, _27622_);
  not (_29181_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_29192_, _15741_, _29181_);
  or (_29203_, _29192_, rst);
  nand (_29214_, _15741_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_29224_, _29214_, _27622_);
  or (_29235_, _29224_, _29203_);
  or (_38304_, _29235_, _29169_);
  nand (_29256_, _27557_, _17536_);
  and (_29267_, _29256_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_29278_, _27557_, _17568_);
  or (_29290_, _29278_, _29267_);
  and (_29301_, _29290_, _15752_);
  and (_29311_, _27622_, ABINPUT[4]);
  not (_29322_, _27622_);
  and (_29333_, _29322_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_29344_, _29333_, _29311_);
  and (_29355_, _29344_, _17320_);
  and (_29366_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_29377_, _29366_, rst);
  or (_29388_, _29377_, _29355_);
  or (_38306_, _29388_, _29301_);
  nand (_29409_, _27557_, _17720_);
  and (_29420_, _29409_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_29431_, _27557_, _17753_);
  or (_29442_, _29431_, _29420_);
  and (_29453_, _29442_, _15752_);
  not (_29464_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_29475_, _27622_, _29464_);
  and (_29485_, _27622_, ABINPUT[5]);
  or (_29496_, _29485_, _29475_);
  and (_29508_, _29496_, _17320_);
  nor (_29519_, _15741_, _29464_);
  or (_29530_, _29519_, rst);
  or (_29541_, _29530_, _29508_);
  or (_38308_, _29541_, _29453_);
  nand (_29562_, _27557_, _17894_);
  and (_29572_, _29562_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_29583_, _27557_, _17926_);
  or (_29594_, _29583_, _29572_);
  and (_29605_, _29594_, _15752_);
  and (_29617_, _27622_, ABINPUT[6]);
  and (_29628_, _29322_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_29639_, _29628_, _29617_);
  and (_29650_, _29639_, _17320_);
  and (_29660_, _27503_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_29671_, _29660_, rst);
  or (_29682_, _29671_, _29650_);
  or (_38310_, _29682_, _29605_);
  nand (_29703_, _27557_, _18067_);
  and (_29714_, _29703_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_29726_, _27557_, _18100_);
  or (_29737_, _29726_, _29714_);
  and (_29747_, _29737_, _15752_);
  not (_29758_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_29769_, _27622_, _29758_);
  and (_29780_, _27622_, ABINPUT[7]);
  or (_29791_, _29780_, _29769_);
  and (_29802_, _29791_, _17320_);
  nor (_29813_, _15741_, _29758_);
  or (_29824_, _29813_, rst);
  or (_29834_, _29824_, _29802_);
  or (_38312_, _29834_, _29747_);
  nand (_29855_, _27557_, _18240_);
  and (_29866_, _29855_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_29877_, _27557_, _18273_);
  or (_29888_, _29877_, _29866_);
  and (_29899_, _29888_, _15752_);
  not (_29910_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_29920_, _27622_, _29910_);
  and (_29931_, _27622_, ABINPUT[8]);
  or (_29942_, _29931_, _29920_);
  and (_29953_, _29942_, _17320_);
  nor (_29964_, _15741_, _29910_);
  or (_29975_, _29964_, rst);
  or (_29986_, _29975_, _29953_);
  or (_38314_, _29986_, _29899_);
  nand (_30006_, _27557_, _18414_);
  and (_30017_, _30006_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_30028_, _27557_, _18447_);
  or (_30039_, _30028_, _30017_);
  and (_30050_, _30039_, _15752_);
  not (_30061_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_30072_, _27622_, _30061_);
  and (_30083_, _27622_, ABINPUT[9]);
  or (_30093_, _30083_, _30072_);
  and (_30104_, _30093_, _17320_);
  nor (_30115_, _15741_, _30061_);
  or (_30126_, _30115_, rst);
  or (_30137_, _30126_, _30104_);
  or (_38316_, _30137_, _30050_);
  and (_30158_, _27741_, ABINPUT[3]);
  not (_30169_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_30179_, _27741_, _30169_);
  or (_30190_, _30179_, _30158_);
  and (_30201_, _30190_, _17320_);
  nor (_30212_, _27807_, _30169_);
  nor (_30223_, _17254_, _30169_);
  or (_30234_, _30223_, _17395_);
  and (_30245_, _30234_, _27807_);
  or (_30256_, _30245_, _30212_);
  and (_30266_, _30256_, _15752_);
  nor (_30277_, _15741_, _30169_);
  or (_30288_, _30277_, rst);
  or (_30299_, _30288_, _30266_);
  or (_38318_, _30299_, _30201_);
  and (_30320_, _27741_, ABINPUT[4]);
  not (_30331_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_30341_, _27741_, _30331_);
  or (_30352_, _30341_, _30320_);
  and (_30363_, _30352_, _17320_);
  nor (_30374_, _17536_, _30331_);
  or (_30385_, _30374_, _17568_);
  and (_30396_, _30385_, _27807_);
  nor (_30407_, _27807_, _30331_);
  or (_30418_, _30407_, _30396_);
  and (_30428_, _30418_, _15752_);
  nor (_30439_, _15741_, _30331_);
  or (_30450_, _30439_, rst);
  or (_30461_, _30450_, _30428_);
  or (_38320_, _30461_, _30363_);
  and (_30482_, _27741_, ABINPUT[5]);
  not (_30493_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_30504_, _27741_, _30493_);
  or (_30514_, _30504_, _30482_);
  and (_30525_, _30514_, _17320_);
  nor (_30536_, _17720_, _30493_);
  or (_30547_, _30536_, _17753_);
  and (_30558_, _30547_, _27807_);
  nor (_30569_, _27807_, _30493_);
  or (_30580_, _30569_, _30558_);
  and (_30591_, _30580_, _15752_);
  nor (_30601_, _15741_, _30493_);
  or (_30612_, _30601_, rst);
  or (_30623_, _30612_, _30591_);
  or (_38322_, _30623_, _30525_);
  and (_30644_, _27741_, ABINPUT[6]);
  not (_30655_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_30666_, _27741_, _30655_);
  or (_30677_, _30666_, _30644_);
  and (_30687_, _30677_, _17320_);
  nor (_30698_, _17894_, _30655_);
  or (_30709_, _30698_, _17926_);
  and (_30720_, _30709_, _27807_);
  nor (_30731_, _27807_, _30655_);
  or (_30742_, _30731_, _30720_);
  and (_30753_, _30742_, _15752_);
  nor (_30764_, _15741_, _30655_);
  or (_30775_, _30764_, rst);
  or (_30785_, _30775_, _30753_);
  or (_38324_, _30785_, _30687_);
  and (_30806_, _27741_, ABINPUT[7]);
  not (_30817_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_30828_, _27741_, _30817_);
  or (_30839_, _30828_, _30806_);
  and (_30850_, _30839_, _17320_);
  nor (_30861_, _18067_, _30817_);
  or (_30871_, _30861_, _18100_);
  and (_30882_, _30871_, _27807_);
  nor (_30893_, _27807_, _30817_);
  or (_30904_, _30893_, _30882_);
  and (_30915_, _30904_, _15752_);
  nor (_30926_, _15741_, _30817_);
  or (_30937_, _30926_, rst);
  or (_30948_, _30937_, _30915_);
  or (_38326_, _30948_, _30850_);
  and (_30969_, _27741_, ABINPUT[8]);
  not (_30980_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_30991_, _27741_, _30980_);
  or (_31002_, _30991_, _30969_);
  and (_31013_, _31002_, _17320_);
  nor (_31024_, _18240_, _30980_);
  or (_31035_, _31024_, _18273_);
  and (_31046_, _31035_, _27807_);
  nor (_31057_, _27807_, _30980_);
  or (_31068_, _31057_, _31046_);
  and (_31079_, _31068_, _15752_);
  nor (_31090_, _15741_, _30980_);
  or (_31101_, _31090_, rst);
  or (_31112_, _31101_, _31079_);
  or (_38328_, _31112_, _31013_);
  and (_31132_, _27741_, ABINPUT[9]);
  not (_31143_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_31154_, _27741_, _31143_);
  or (_31165_, _31154_, _31132_);
  and (_31176_, _31165_, _17320_);
  nor (_31187_, _18414_, _31143_);
  or (_31198_, _31187_, _18447_);
  and (_31209_, _31198_, _27807_);
  nor (_31220_, _27807_, _31143_);
  or (_31231_, _31220_, _31209_);
  and (_31242_, _31231_, _15752_);
  nor (_31253_, _15741_, _31143_);
  or (_31264_, _31253_, rst);
  or (_31275_, _31264_, _31242_);
  or (_38329_, _31275_, _31176_);
  and (_31296_, _27947_, ABINPUT[3]);
  not (_31307_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_31318_, _27947_, _31307_);
  or (_31329_, _31318_, _31296_);
  and (_31340_, _31329_, _17320_);
  nor (_31351_, _17254_, _31307_);
  or (_31362_, _31351_, _17395_);
  and (_31373_, _31362_, _28045_);
  nor (_31384_, _28045_, _31307_);
  or (_31395_, _31384_, _31373_);
  and (_31406_, _31395_, _15752_);
  nor (_31417_, _15741_, _31307_);
  or (_31428_, _31417_, rst);
  or (_31439_, _31428_, _31406_);
  or (_38331_, _31439_, _31340_);
  and (_31460_, _27947_, ABINPUT[4]);
  not (_31471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_31482_, _27947_, _31471_);
  or (_31493_, _31482_, _31460_);
  and (_31504_, _31493_, _17320_);
  nor (_31514_, _17536_, _31471_);
  or (_31525_, _31514_, _17568_);
  and (_31536_, _31525_, _28045_);
  nor (_31547_, _28045_, _31471_);
  or (_31558_, _31547_, _31536_);
  and (_31569_, _31558_, _15752_);
  nor (_31580_, _15741_, _31471_);
  or (_31591_, _31580_, rst);
  or (_31602_, _31591_, _31569_);
  or (_38333_, _31602_, _31504_);
  and (_31623_, _27947_, ABINPUT[5]);
  not (_31634_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_31645_, _27947_, _31634_);
  or (_31656_, _31645_, _31623_);
  and (_31667_, _31656_, _17320_);
  nor (_31678_, _17720_, _31634_);
  or (_31689_, _31678_, _17753_);
  and (_31700_, _31689_, _28045_);
  nor (_31711_, _28045_, _31634_);
  or (_31722_, _31711_, _31700_);
  and (_31733_, _31722_, _15752_);
  nor (_31744_, _15741_, _31634_);
  or (_31755_, _31744_, rst);
  or (_31766_, _31755_, _31733_);
  or (_38335_, _31766_, _31667_);
  and (_31787_, _27947_, ABINPUT[6]);
  not (_31798_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_31809_, _27947_, _31798_);
  or (_31820_, _31809_, _31787_);
  and (_31831_, _31820_, _17320_);
  nor (_31842_, _17894_, _31798_);
  or (_31853_, _31842_, _17926_);
  and (_31864_, _31853_, _28045_);
  nor (_31875_, _28045_, _31798_);
  or (_31886_, _31875_, _31864_);
  and (_31896_, _31886_, _15752_);
  nor (_31907_, _15741_, _31798_);
  or (_31918_, _31907_, rst);
  or (_31929_, _31918_, _31896_);
  or (_38337_, _31929_, _31831_);
  and (_31950_, _27947_, ABINPUT[7]);
  not (_31961_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_31972_, _27947_, _31961_);
  or (_31983_, _31972_, _31950_);
  and (_31994_, _31983_, _17320_);
  nor (_32005_, _18067_, _31961_);
  or (_32016_, _32005_, _18100_);
  and (_32027_, _32016_, _28045_);
  nor (_32038_, _28045_, _31961_);
  or (_32049_, _32038_, _32027_);
  and (_32060_, _32049_, _15752_);
  nor (_32071_, _15741_, _31961_);
  or (_32082_, _32071_, rst);
  or (_32093_, _32082_, _32060_);
  or (_38339_, _32093_, _31994_);
  and (_32114_, _27947_, ABINPUT[8]);
  not (_32125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_32136_, _27947_, _32125_);
  or (_32147_, _32136_, _32114_);
  and (_32158_, _32147_, _17320_);
  nor (_32169_, _18240_, _32125_);
  or (_32180_, _32169_, _18273_);
  and (_32191_, _32180_, _28045_);
  nor (_32202_, _28045_, _32125_);
  or (_32213_, _32202_, _32191_);
  and (_32224_, _32213_, _15752_);
  nor (_32235_, _15741_, _32125_);
  or (_32246_, _32235_, rst);
  or (_32256_, _32246_, _32224_);
  or (_38341_, _32256_, _32158_);
  and (_32277_, _27947_, ABINPUT[9]);
  not (_32288_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_32299_, _27947_, _32288_);
  or (_32310_, _32299_, _32277_);
  and (_32321_, _32310_, _17320_);
  nor (_32332_, _18414_, _32288_);
  or (_32343_, _32332_, _18447_);
  and (_32354_, _32343_, _28045_);
  nor (_32365_, _28045_, _32288_);
  or (_32376_, _32365_, _32354_);
  and (_32387_, _32376_, _15752_);
  nor (_32398_, _15741_, _32288_);
  or (_32409_, _32398_, rst);
  or (_32420_, _32409_, _32387_);
  or (_38343_, _32420_, _32321_);
  and (_32441_, _25326_, _16557_);
  and (_32452_, _32441_, _27730_);
  nor (_32463_, _26224_, _16547_);
  and (_32474_, _32463_, _27730_);
  and (_32485_, _32474_, _17145_);
  nand (_32496_, _32485_, _17178_);
  or (_32507_, _32485_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_32518_, _32507_, _32496_);
  or (_32529_, _32518_, _32452_);
  nand (_32540_, _32452_, _27438_);
  and (_32551_, _32540_, _39026_);
  and (_38937_, _32551_, _32529_);
  and (_32572_, _32441_, _27936_);
  not (_32583_, _16721_);
  and (_32594_, _32463_, _32583_);
  and (_32604_, _32594_, _16383_);
  and (_32615_, _32604_, _28034_);
  and (_32626_, _32615_, _17145_);
  nand (_32637_, _32626_, _17178_);
  or (_32648_, _32626_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_32659_, _32648_, _32637_);
  or (_32670_, _32659_, _32572_);
  nand (_32681_, _32572_, _27438_);
  and (_32692_, _32681_, _39026_);
  and (_38973_, _32692_, _32670_);
  and (_32733_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_32744_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _39026_);
  and (_38993_, _32744_, _32733_);
  not (_32765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_32776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _32765_);
  not (_32787_, _32776_);
  not (_32798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_32809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_32820_, _32809_, _32798_);
  not (_32831_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_32842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_32853_, _32842_, _32831_);
  nor (_32864_, _32853_, _32820_);
  not (_32875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_32886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_32897_, _32886_, _32875_);
  not (_32908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_32919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_32930_, _32919_, _32908_);
  nor (_32941_, _32930_, _32897_);
  and (_32952_, _32941_, _32864_);
  nor (_32963_, _32952_, _32787_);
  and (_32973_, _32809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_32984_, _32842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_32995_, _32984_, _32973_);
  and (_33006_, _32886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_33017_, _32919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_33028_, _33017_, _33006_);
  and (_33039_, _33028_, _32995_);
  nand (_33050_, _33039_, _32765_);
  or (_33061_, _33050_, _32963_);
  not (_33072_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _33072_);
  nand (_33094_, _33083_, _32733_);
  and (_33105_, _33094_, _39026_);
  and (_38995_, _33105_, _33061_);
  and (_33126_, _32897_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_33137_, _33126_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_33148_, _32864_);
  and (_33159_, _32930_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33170_, _33159_, _33148_);
  and (_33181_, _33170_, _33137_);
  and (_33192_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _33072_);
  and (_33203_, _33192_, _33148_);
  or (_33214_, _33203_, _33181_);
  and (_33225_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_33236_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _33072_);
  nor (_33247_, _33236_, _33225_);
  and (_33258_, _33247_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_33269_, _33258_, _32765_);
  nor (_33280_, _33269_, _33039_);
  not (_33291_, _33280_);
  and (_33302_, _33291_, _32963_);
  and (_33313_, _33302_, _33214_);
  or (_33324_, _33313_, _32733_);
  and (_33334_, _33006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_33345_, _32995_);
  or (_33356_, _33345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_33367_, _33356_, _33334_);
  not (_33378_, _33017_);
  and (_33389_, _33378_, _32995_);
  or (_33400_, _33192_, _33389_);
  and (_33411_, _33400_, _33367_);
  and (_33422_, _33411_, _33280_);
  nor (_33433_, _33280_, _32963_);
  and (_33444_, _33433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_33455_, _33444_, _33422_);
  or (_33466_, _33455_, _33324_);
  not (_33477_, _32733_);
  or (_33488_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_33499_, _33488_, _39026_);
  and (_38997_, _33499_, _33466_);
  and (_33520_, _32463_, _22917_);
  and (_33531_, _33520_, _17894_);
  nand (_33542_, _33531_, _17178_);
  and (_33553_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_33564_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _33072_);
  and (_33575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33586_, _33575_, _33564_);
  nor (_33597_, _33586_, _32765_);
  nand (_33608_, _33597_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_33619_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _33072_);
  and (_33630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33641_, _33630_, _33619_);
  nor (_33652_, _33641_, _32765_);
  and (_33663_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_33674_, _33663_, _33192_);
  nand (_33685_, _33674_, _33652_);
  or (_33695_, _33685_, _33608_);
  and (_33706_, _33695_, _33553_);
  or (_33717_, _33706_, _33531_);
  and (_33728_, _33717_, _33542_);
  and (_33739_, _32441_, _22917_);
  or (_33750_, _33739_, _33728_);
  nand (_33761_, _33739_, _28541_);
  and (_33772_, _33761_, _39026_);
  and (_39017_, _33772_, _33750_);
  not (_33793_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_33804_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _33793_);
  nor (_33815_, _33674_, _32765_);
  or (_33826_, _33815_, _33652_);
  or (_33837_, _33826_, _33608_);
  and (_33848_, _33837_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_33859_, _33848_, _33804_);
  nand (_33870_, _33520_, _17536_);
  and (_33881_, _33870_, _33859_);
  nor (_33892_, _33870_, _17178_);
  or (_33903_, _33892_, _33739_);
  or (_33914_, _33903_, _33881_);
  nand (_33925_, _33739_, _25456_);
  and (_33936_, _33925_, _39026_);
  and (_39019_, _33936_, _33914_);
  not (_33957_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_33968_, _33597_, _33957_);
  or (_33979_, _33968_, _33685_);
  and (_33990_, _33979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand (_34001_, _33520_, _18240_);
  and (_34012_, _34001_, _33990_);
  and (_34022_, _33520_, _18273_);
  or (_34033_, _34022_, _33739_);
  or (_34044_, _34033_, _34012_);
  nand (_34055_, _33739_, _25866_);
  and (_34066_, _34055_, _39026_);
  and (_39020_, _34066_, _34044_);
  nand (_34087_, _33815_, _33641_);
  or (_34098_, _34087_, _33968_);
  and (_34109_, _34098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand (_34120_, _33520_, _17145_);
  and (_34131_, _34120_, _34109_);
  and (_34142_, _33520_, _25207_);
  or (_34153_, _34142_, _33739_);
  or (_34164_, _34153_, _34131_);
  nand (_34175_, _33739_, _27438_);
  and (_34186_, _34175_, _39026_);
  and (_39022_, _34186_, _34164_);
  nand (_34207_, _33520_, _18414_);
  and (_34218_, _34207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_34229_, _33520_, _18447_);
  or (_34240_, _34229_, _33739_);
  or (_34251_, _34240_, _34218_);
  not (_34262_, ABINPUT[9]);
  nand (_34273_, _33739_, _34262_);
  and (_34284_, _34273_, _39026_);
  and (_39024_, _34284_, _34251_);
  and (_34305_, _33433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_34316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _33072_);
  nor (_34327_, _34316_, _33083_);
  nor (_34338_, _34327_, _33291_);
  or (_34349_, _34338_, _32733_);
  or (_34359_, _34349_, _34305_);
  or (_34370_, _34327_, _33477_);
  and (_34381_, _34370_, _39026_);
  and (_39028_, _34381_, _34359_);
  and (_34402_, _32897_, _33072_);
  or (_34413_, _34402_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_34424_, _32930_, _33072_);
  nor (_34435_, _34424_, _33148_);
  and (_34446_, _34435_, _34413_);
  and (_34457_, _33663_, _33148_);
  or (_34468_, _34457_, _34446_);
  and (_34479_, _34468_, _33302_);
  or (_34490_, _34479_, _32733_);
  and (_34501_, _33006_, _33072_);
  or (_34512_, _33345_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_34523_, _34512_, _34501_);
  or (_34534_, _33663_, _33389_);
  and (_34545_, _34534_, _34523_);
  and (_34556_, _34545_, _33280_);
  and (_34567_, _33433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_34578_, _34567_, _34556_);
  or (_34589_, _34578_, _34490_);
  or (_34600_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_34611_, _34600_, _39026_);
  and (_39030_, _34611_, _34589_);
  nor (_34632_, _32733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_34643_, _34632_, _33280_);
  nand (_34654_, _34632_, _32963_);
  and (_34665_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _39026_);
  nand (_34675_, _34665_, _34654_);
  nor (_39031_, _34675_, _34643_);
  nor (_34696_, _32733_, _33072_);
  and (_34707_, _34696_, _33280_);
  nand (_34718_, _34696_, _32963_);
  and (_34729_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _39026_);
  nand (_34740_, _34729_, _34718_);
  nor (_39033_, _34740_, _34707_);
  nor (_34771_, _33433_, _32733_);
  and (_34782_, _32733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_34793_, _34782_, _34771_);
  and (_40001_, _34793_, _39026_);
  and (_34814_, _32733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_34825_, _34814_, _34771_);
  and (_40003_, _34825_, _39026_);
  and (_34846_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _39026_);
  and (_40005_, _34846_, _32733_);
  not (_34867_, _32853_);
  nor (_34878_, _32897_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_34889_, _34878_, _32930_);
  or (_34900_, _34889_, _32820_);
  and (_34911_, _34900_, _34867_);
  and (_34922_, _34911_, _33302_);
  not (_34933_, _32984_);
  or (_34944_, _33006_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_34955_, _34944_, _33378_);
  or (_34966_, _34955_, _32973_);
  and (_34977_, _34966_, _34933_);
  and (_34987_, _34977_, _33280_);
  or (_34998_, _34987_, _32733_);
  or (_35009_, _34998_, _34922_);
  or (_35020_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_35031_, _35020_, _39026_);
  and (_40007_, _35031_, _35009_);
  nand (_35052_, _32864_, _32776_);
  or (_35063_, _35052_, _32941_);
  nor (_35074_, _35063_, _33280_);
  or (_35085_, _33028_, _33345_);
  nor (_35096_, _35085_, _33269_);
  or (_35107_, _35096_, _32733_);
  or (_35118_, _35107_, _35074_);
  or (_35129_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_35140_, _35129_, _39026_);
  and (_40009_, _35140_, _35118_);
  and (_35161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _39026_);
  and (_40011_, _35161_, _32733_);
  and (_35182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _39026_);
  and (_40013_, _35182_, _32733_);
  nand (_35203_, _34632_, _33433_);
  nor (_35214_, _33280_, _32733_);
  or (_35225_, _35214_, _33072_);
  and (_35236_, _35225_, _39026_);
  and (_40015_, _35236_, _35203_);
  not (_35257_, _34771_);
  and (_35269_, _35257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_35280_, _34501_);
  and (_35290_, _35280_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_35301_, _33017_, _33072_);
  or (_35312_, _35301_, _32973_);
  or (_35323_, _35312_, _35290_);
  not (_35334_, _32973_);
  or (_35345_, _33575_, _35334_);
  and (_35356_, _35345_, _35323_);
  or (_35367_, _35356_, _32984_);
  or (_35378_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _33072_);
  or (_35389_, _35378_, _34933_);
  and (_35400_, _35389_, _33280_);
  and (_35411_, _35400_, _35367_);
  not (_35422_, _34402_);
  and (_35433_, _35422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_35444_, _34424_, _32820_);
  or (_35455_, _35444_, _35433_);
  not (_35466_, _32820_);
  or (_35477_, _33575_, _35466_);
  and (_35489_, _35477_, _35455_);
  or (_35500_, _35489_, _32853_);
  or (_35511_, _35378_, _34867_);
  and (_35522_, _35511_, _33302_);
  and (_35533_, _35522_, _35500_);
  or (_35544_, _35533_, _35411_);
  and (_35555_, _35544_, _33477_);
  or (_35566_, _35555_, _35269_);
  and (_40017_, _35566_, _39026_);
  and (_35587_, _35422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_35597_, _35587_, _35444_);
  or (_35608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _33072_);
  or (_35619_, _35608_, _35466_);
  and (_35630_, _35619_, _34867_);
  and (_35641_, _35630_, _35597_);
  and (_35652_, _33630_, _32853_);
  or (_35663_, _35652_, _35641_);
  and (_35674_, _35663_, _33302_);
  and (_35685_, _35280_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_35696_, _35685_, _35312_);
  or (_35707_, _35608_, _35334_);
  and (_35718_, _35707_, _35696_);
  or (_35729_, _35718_, _32984_);
  or (_35740_, _33630_, _34933_);
  and (_35751_, _35740_, _33280_);
  and (_35762_, _35751_, _35729_);
  and (_35773_, _33433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_35784_, _35773_, _32733_);
  or (_35795_, _35784_, _35762_);
  or (_35806_, _35795_, _35674_);
  or (_35817_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_35828_, _35817_, _39026_);
  and (_40019_, _35828_, _35806_);
  and (_35849_, _35257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_35860_, _33334_);
  and (_35871_, _35860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_35882_, _33017_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_35893_, _35882_, _32973_);
  or (_35904_, _35893_, _35871_);
  or (_35911_, _33564_, _35334_);
  and (_35919_, _35911_, _35904_);
  or (_35927_, _35919_, _32984_);
  or (_35934_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_35942_, _35934_, _34933_);
  and (_35950_, _35942_, _33280_);
  and (_35957_, _35950_, _35927_);
  not (_35965_, _33126_);
  and (_35969_, _35965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_35970_, _33159_, _32820_);
  or (_35971_, _35970_, _35969_);
  or (_35976_, _33564_, _35466_);
  and (_35987_, _35976_, _35971_);
  or (_35998_, _35987_, _32853_);
  or (_36009_, _35934_, _34867_);
  and (_36020_, _36009_, _33302_);
  and (_36031_, _36020_, _35998_);
  or (_36042_, _36031_, _35957_);
  and (_36053_, _36042_, _33477_);
  or (_36064_, _36053_, _35849_);
  and (_40021_, _36064_, _39026_);
  and (_36085_, _35965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_36096_, _36085_, _35970_);
  or (_36107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_36118_, _36107_, _35466_);
  and (_36129_, _36118_, _34867_);
  and (_36140_, _36129_, _36096_);
  and (_36151_, _33619_, _32853_);
  or (_36162_, _36151_, _36140_);
  and (_36172_, _36162_, _33302_);
  and (_36183_, _35860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_36194_, _36183_, _35893_);
  or (_36204_, _36107_, _35334_);
  and (_36215_, _36204_, _36194_);
  or (_36226_, _36215_, _32984_);
  or (_36236_, _33619_, _34933_);
  and (_36247_, _36236_, _33280_);
  and (_36258_, _36247_, _36226_);
  and (_36269_, _33433_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_36280_, _36269_, _32733_);
  or (_36291_, _36280_, _36258_);
  or (_36302_, _36291_, _36172_);
  or (_36312_, _33477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_36323_, _36312_, _39026_);
  and (_40023_, _36323_, _36302_);
  and (_36344_, _34654_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_36355_, _36344_, _34643_);
  and (_40025_, _36355_, _39026_);
  and (_36376_, _34718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_36387_, _36376_, _34707_);
  and (_40027_, _36387_, _39026_);
  and (_36408_, _33520_, _17254_);
  nand (_36419_, _36408_, _17178_);
  or (_36430_, _36408_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_36441_, _36430_, _36419_);
  or (_36452_, _36441_, _33739_);
  not (_36463_, ABINPUT[3]);
  nand (_36474_, _33739_, _36463_);
  and (_36485_, _36474_, _39026_);
  and (_40029_, _36485_, _36452_);
  nand (_36506_, _33520_, _17720_);
  and (_36517_, _36506_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_36528_, _33520_, _17753_);
  or (_36539_, _36528_, _33739_);
  or (_36550_, _36539_, _36517_);
  not (_36561_, ABINPUT[5]);
  nand (_36572_, _33739_, _36561_);
  and (_36583_, _36572_, _39026_);
  and (_40031_, _36583_, _36550_);
  nand (_36604_, _33520_, _18067_);
  and (_36615_, _36604_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_36626_, _33520_, _18100_);
  or (_36637_, _36626_, _33739_);
  or (_36648_, _36637_, _36615_);
  not (_36659_, ABINPUT[7]);
  nand (_36670_, _33739_, _36659_);
  and (_36681_, _36670_, _39026_);
  and (_40033_, _36681_, _36648_);
  nand (_36702_, _32474_, _17254_);
  and (_36713_, _36702_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_36724_, _32474_, _17395_);
  or (_36735_, _36724_, _32452_);
  or (_36746_, _36735_, _36713_);
  nand (_36757_, _32452_, _36463_);
  and (_36768_, _36757_, _39026_);
  and (_40035_, _36768_, _36746_);
  nand (_36789_, _32474_, _17536_);
  and (_36800_, _36789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_36811_, _32474_, _17568_);
  or (_36822_, _36811_, _32452_);
  or (_36833_, _36822_, _36800_);
  nand (_36844_, _32452_, _25456_);
  and (_36855_, _36844_, _39026_);
  and (_40037_, _36855_, _36833_);
  and (_36876_, _32474_, _17720_);
  or (_36887_, _36876_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand (_36898_, _36876_, _17178_);
  and (_36909_, _36898_, _36887_);
  or (_36920_, _36909_, _32452_);
  nand (_36931_, _32452_, _36561_);
  and (_36942_, _36931_, _39026_);
  and (_40039_, _36942_, _36920_);
  nand (_36963_, _32474_, _17894_);
  and (_36974_, _36963_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_36985_, _32474_, _17926_);
  or (_36996_, _36985_, _32452_);
  or (_37007_, _36996_, _36974_);
  nand (_37018_, _32452_, _28541_);
  and (_37029_, _37018_, _39026_);
  and (_40041_, _37029_, _37007_);
  nand (_37050_, _32474_, _18067_);
  and (_37061_, _37050_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_37072_, _32474_, _18100_);
  or (_37083_, _37072_, _32452_);
  or (_37094_, _37083_, _37061_);
  nand (_37105_, _32452_, _36659_);
  and (_37116_, _37105_, _39026_);
  and (_40043_, _37116_, _37094_);
  nand (_37137_, _32474_, _18240_);
  and (_37148_, _37137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_37159_, _32474_, _18273_);
  or (_37170_, _37159_, _32452_);
  or (_37181_, _37170_, _37148_);
  nand (_37192_, _32452_, _25866_);
  and (_37203_, _37192_, _39026_);
  and (_40045_, _37203_, _37181_);
  nand (_37212_, _32474_, _18414_);
  and (_37223_, _37212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_37225_, _32474_, _18447_);
  or (_37226_, _37225_, _32452_);
  or (_37227_, _37226_, _37223_);
  nand (_37228_, _32452_, _34262_);
  and (_37229_, _37228_, _39026_);
  and (_40047_, _37229_, _37227_);
  nand (_37230_, _32615_, _17254_);
  and (_37231_, _37230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_37232_, _32615_, _17395_);
  or (_37233_, _37232_, _32572_);
  or (_37234_, _37233_, _37231_);
  nand (_37235_, _32572_, _36463_);
  and (_37236_, _37235_, _39026_);
  and (_40049_, _37236_, _37234_);
  nand (_37237_, _32615_, _17536_);
  and (_37238_, _37237_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_37239_, _32615_, _17568_);
  or (_37240_, _37239_, _32572_);
  or (_37241_, _37240_, _37238_);
  nand (_37242_, _32572_, _25456_);
  and (_37243_, _37242_, _39026_);
  and (_40051_, _37243_, _37241_);
  and (_37244_, _32615_, _17720_);
  or (_37245_, _37244_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_37246_, _37244_, _17178_);
  and (_37247_, _37246_, _37245_);
  or (_37248_, _37247_, _32572_);
  nand (_37249_, _32572_, _36561_);
  and (_37250_, _37249_, _39026_);
  and (_40053_, _37250_, _37248_);
  nand (_37251_, _32615_, _17894_);
  and (_37252_, _37251_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_37253_, _32615_, _17926_);
  or (_37254_, _37253_, _32572_);
  or (_37255_, _37254_, _37252_);
  nand (_37256_, _32572_, _28541_);
  and (_37257_, _37256_, _39026_);
  and (_40055_, _37257_, _37255_);
  nand (_37258_, _32615_, _18067_);
  and (_37259_, _37258_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_37260_, _32615_, _18100_);
  or (_37261_, _37260_, _32572_);
  or (_37262_, _37261_, _37259_);
  nand (_37263_, _32572_, _36659_);
  and (_37264_, _37263_, _39026_);
  and (_40057_, _37264_, _37262_);
  nand (_37265_, _32615_, _18240_);
  and (_37266_, _37265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_37267_, _32615_, _18273_);
  or (_37268_, _37267_, _32572_);
  or (_37269_, _37268_, _37266_);
  nand (_37270_, _32572_, _25866_);
  and (_37271_, _37270_, _39026_);
  and (_40059_, _37271_, _37269_);
  nand (_37272_, _32615_, _18414_);
  and (_37273_, _37272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_37274_, _32615_, _18447_);
  or (_37275_, _37274_, _32572_);
  or (_37276_, _37275_, _37273_);
  nand (_37277_, _32572_, _34262_);
  and (_37278_, _37277_, _39026_);
  and (_40061_, _37278_, _37276_);
  not (_37279_, _22852_);
  and (_37280_, _22852_, _21645_);
  not (_37281_, _37280_);
  nor (_37282_, _37281_, _22698_);
  not (_37283_, _18653_);
  and (_37284_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_37285_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_37286_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_37287_, _37286_, _37285_);
  and (_37288_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_37289_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_37290_, _37289_, _37288_);
  and (_37291_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_37292_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_37293_, _37292_, _37291_);
  and (_37294_, _37293_, _37290_);
  and (_37295_, _37294_, _37287_);
  nor (_37296_, _18729_, _37283_);
  not (_37297_, _37296_);
  nor (_37298_, _37297_, _37295_);
  nor (_37299_, _37298_, _37284_);
  not (_37300_, _37299_);
  and (_37301_, _37300_, _37282_);
  nor (_37302_, _37301_, _37279_);
  and (_37303_, _22852_, _22709_);
  not (_37304_, _23389_);
  and (_37305_, _37304_, _37303_);
  not (_37306_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_37307_, _15719_, _16351_);
  and (_37308_, _21111_, _17004_);
  nor (_37309_, _21111_, _17004_);
  nor (_37310_, _37309_, _37308_);
  and (_37311_, _37310_, _17123_);
  not (_37312_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_37313_, _25337_, _37312_);
  nor (_37314_, _37313_, _25694_);
  and (_37315_, _37314_, _16557_);
  nor (_37316_, _37314_, _16557_);
  nor (_37317_, _37316_, _37315_);
  and (_37318_, _37317_, _16873_);
  and (_37319_, _37318_, _37311_);
  and (_37320_, _37319_, _37307_);
  and (_37321_, _37320_, _37306_);
  nor (_37322_, _37314_, _21111_);
  and (_37323_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_37324_, _37314_, _21111_);
  and (_37325_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_37326_, _37325_, _37323_);
  nor (_37327_, _37314_, _21438_);
  and (_37328_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_37329_, _37314_, _21438_);
  and (_37330_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_37331_, _37330_, _37328_);
  and (_37332_, _37331_, _37326_);
  nor (_37333_, _37332_, _37321_);
  and (_37334_, _37321_, ABINPUT[10]);
  nor (_37335_, _37334_, _37333_);
  not (_37336_, _37335_);
  not (_37337_, _21645_);
  and (_37338_, _22698_, _37337_);
  and (_37339_, _37338_, _22852_);
  and (_37340_, _37339_, _37336_);
  nor (_37341_, _37340_, _37305_);
  and (_37342_, _37341_, _37302_);
  nor (_37343_, _21677_, _22445_);
  and (_37344_, _37343_, _22357_);
  and (_37345_, _21754_, _22148_);
  nor (_37346_, _22027_, _22203_);
  nor (_37347_, _21863_, _22214_);
  and (_37348_, _37347_, _37346_);
  and (_37349_, _37348_, _37345_);
  and (_37350_, _37349_, _37344_);
  nor (_37351_, _37350_, _18609_);
  not (_37352_, _21557_);
  nor (_37353_, _21754_, _37352_);
  nor (_37354_, _37353_, _37351_);
  not (_37355_, _37354_);
  and (_37356_, _37355_, _37342_);
  and (_37357_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_37358_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_37359_, _37358_, _37357_);
  and (_37360_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_37361_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_37362_, _37361_, _37360_);
  and (_37363_, _37362_, _37359_);
  nor (_37364_, _37363_, _37321_);
  and (_37365_, _37321_, ABINPUT[8]);
  nor (_37366_, _37365_, _37364_);
  not (_37367_, _37366_);
  and (_37368_, _37367_, _37339_);
  not (_37369_, _37368_);
  and (_37370_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_37371_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_37372_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_37373_, _37372_, _37371_);
  and (_37374_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_37375_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_37376_, _37375_, _37374_);
  and (_37377_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_37378_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_37379_, _37378_, _37377_);
  and (_37380_, _37379_, _37376_);
  and (_37381_, _37380_, _37373_);
  nor (_37382_, _37381_, _37297_);
  nor (_37383_, _37382_, _37370_);
  not (_37384_, _37383_);
  and (_37385_, _37384_, _37282_);
  not (_37386_, _37385_);
  and (_37387_, _37279_, _21645_);
  and (_37388_, _37387_, _22698_);
  not (_37389_, _22709_);
  and (_37390_, _23864_, _22852_);
  nor (_37391_, _37390_, _37389_);
  nor (_37392_, _37391_, _37388_);
  and (_37393_, _37392_, _37386_);
  and (_37394_, _37393_, _37369_);
  not (_37395_, _37394_);
  and (_37396_, _37395_, _37356_);
  not (_37397_, _23638_);
  and (_37398_, _37397_, _37303_);
  not (_37399_, _37398_);
  and (_37400_, _37280_, _22698_);
  and (_37401_, _37400_, _19318_);
  and (_37402_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_37403_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_37404_, _37403_, _37402_);
  and (_37405_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_37406_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37407_, _37406_, _37405_);
  and (_37408_, _37407_, _37404_);
  nor (_37409_, _37408_, _37321_);
  and (_37410_, _37321_, ABINPUT[5]);
  nor (_37411_, _37410_, _37409_);
  not (_37412_, _37411_);
  and (_37413_, _37412_, _37339_);
  and (_37414_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_37415_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_37416_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_37417_, _37416_, _37415_);
  and (_37418_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_37419_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_37420_, _37419_, _37418_);
  and (_37421_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_37422_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_37423_, _37422_, _37421_);
  and (_37424_, _37423_, _37420_);
  and (_37425_, _37424_, _37417_);
  nor (_37426_, _37425_, _37297_);
  nor (_37427_, _37426_, _37414_);
  not (_37428_, _37427_);
  and (_37429_, _37428_, _37282_);
  or (_37430_, _37429_, _37413_);
  nor (_37431_, _37430_, _37401_);
  and (_37432_, _37431_, _37399_);
  nor (_37433_, _37432_, _37355_);
  nor (_37434_, _37433_, _37396_);
  not (_37435_, _37434_);
  not (_37436_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_37437_, _25337_, _37436_);
  nor (_37438_, _37437_, _25780_);
  not (_37439_, _37438_);
  and (_37440_, _37439_, _37400_);
  not (_37441_, _37440_);
  and (_37442_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_37443_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_37444_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_37445_, _37444_, _37443_);
  and (_37446_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_37447_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_37448_, _37447_, _37446_);
  and (_37449_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_37450_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_37451_, _37450_, _37449_);
  and (_37452_, _37451_, _37448_);
  and (_37453_, _37452_, _37445_);
  nor (_37454_, _37453_, _37297_);
  nor (_37455_, _37454_, _37442_);
  not (_37456_, _37455_);
  and (_37457_, _37456_, _37282_);
  nor (_37458_, _37457_, _37387_);
  and (_37459_, _37458_, _37441_);
  not (_37460_, _23789_);
  and (_37461_, _37460_, _37303_);
  and (_37462_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_37463_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_37464_, _37463_, _37462_);
  and (_37465_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_37466_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_37467_, _37466_, _37465_);
  and (_37468_, _37467_, _37464_);
  nor (_37469_, _37468_, _37321_);
  and (_37470_, _37321_, ABINPUT[7]);
  nor (_37471_, _37470_, _37469_);
  not (_37472_, _37471_);
  and (_37473_, _37472_, _37339_);
  nor (_37474_, _37473_, _37461_);
  and (_37475_, _37474_, _37459_);
  not (_37476_, _37475_);
  and (_37477_, _37476_, _37356_);
  and (_37478_, _37400_, _19606_);
  not (_37479_, _37478_);
  and (_37480_, _37338_, _37279_);
  and (_37481_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_37482_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_37483_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_37484_, _37483_, _37482_);
  and (_37485_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_37486_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_37487_, _37486_, _37485_);
  and (_37488_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_37489_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_37490_, _37489_, _37488_);
  and (_37491_, _37490_, _37487_);
  and (_37492_, _37491_, _37484_);
  nor (_37493_, _37492_, _37297_);
  nor (_37494_, _37493_, _37481_);
  not (_37495_, _37494_);
  and (_37496_, _37495_, _37282_);
  nor (_37497_, _37496_, _37480_);
  and (_37498_, _37497_, _37479_);
  not (_37499_, _23562_);
  and (_37500_, _37499_, _37303_);
  and (_37501_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_37502_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_37503_, _37502_, _37501_);
  and (_37504_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_37505_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_37506_, _37505_, _37504_);
  and (_37507_, _37506_, _37503_);
  nor (_37508_, _37507_, _37321_);
  and (_37509_, _37321_, ABINPUT[4]);
  nor (_37510_, _37509_, _37508_);
  not (_37511_, _37510_);
  and (_37512_, _37511_, _37339_);
  nor (_37513_, _37512_, _37500_);
  and (_37514_, _37513_, _37498_);
  nor (_37515_, _37514_, _37355_);
  nor (_37516_, _37515_, _37477_);
  not (_37517_, _23713_);
  and (_37518_, _37517_, _37303_);
  not (_37519_, _37518_);
  not (_37520_, _37314_);
  and (_37521_, _37400_, _37520_);
  and (_37522_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37523_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_37524_, _37523_, _37522_);
  and (_37525_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_37526_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37527_, _37526_, _37525_);
  and (_37528_, _37527_, _37524_);
  nor (_37529_, _37528_, _37321_);
  and (_37530_, _37321_, ABINPUT[6]);
  nor (_37531_, _37530_, _37529_);
  not (_37532_, _37531_);
  and (_37533_, _37532_, _37339_);
  and (_37534_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_37535_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_37536_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_37537_, _37536_, _37535_);
  and (_37538_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_37539_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_37540_, _37539_, _37538_);
  and (_37541_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_37542_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_37543_, _37542_, _37541_);
  and (_37544_, _37543_, _37540_);
  and (_37545_, _37544_, _37537_);
  nor (_37546_, _37545_, _37297_);
  nor (_37547_, _37546_, _37534_);
  not (_37548_, _37547_);
  and (_37549_, _37548_, _37282_);
  or (_37550_, _37549_, _37533_);
  nor (_37551_, _37550_, _37521_);
  and (_37552_, _37551_, _37519_);
  not (_37553_, _37552_);
  and (_37554_, _37553_, _37356_);
  not (_37555_, _23486_);
  and (_37556_, _37555_, _37303_);
  not (_37557_, _37556_);
  and (_37558_, _37400_, _21111_);
  and (_37559_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  not (_37560_, _37559_);
  and (_37561_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_37562_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_37563_, _37562_, _37561_);
  and (_37564_, _37563_, _37560_);
  and (_37565_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_37566_, _37565_, _37321_);
  and (_37567_, _37566_, _37564_);
  and (_37568_, _37321_, _36463_);
  or (_37569_, _37568_, _37567_);
  not (_37570_, _37569_);
  and (_37571_, _37570_, _37339_);
  and (_37572_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_37573_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_37574_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_37575_, _37574_, _37573_);
  and (_37576_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_37577_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_37578_, _37577_, _37576_);
  and (_37579_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_37580_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_37581_, _37580_, _37579_);
  and (_37582_, _37581_, _37578_);
  and (_37583_, _37582_, _37575_);
  nor (_37584_, _37583_, _37297_);
  nor (_37585_, _37584_, _37572_);
  not (_37586_, _37585_);
  and (_37587_, _37586_, _37282_);
  or (_37588_, _37587_, _37571_);
  nor (_37589_, _37588_, _37558_);
  and (_37590_, _37589_, _37557_);
  nor (_37591_, _37590_, _37355_);
  nor (_37592_, _37591_, _37554_);
  or (_37593_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_37594_, _37592_);
  or (_37595_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_37596_, _37595_, _37593_);
  or (_37597_, _37596_, _37516_);
  and (_37598_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_37599_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_37600_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_37601_, _37600_, _37599_);
  and (_37602_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_37603_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_37604_, _37603_, _37602_);
  and (_37605_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_37606_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_37607_, _37606_, _37605_);
  and (_37608_, _37607_, _37604_);
  and (_37609_, _37608_, _37601_);
  nor (_37610_, _37609_, _37297_);
  nor (_37611_, _37610_, _37598_);
  not (_37612_, _37611_);
  and (_37613_, _37612_, _37282_);
  nor (_37614_, _37338_, _22852_);
  nor (_37615_, _37614_, _37613_);
  and (_37616_, _37322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_37617_, _37324_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_37618_, _37617_, _37616_);
  and (_37619_, _37327_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_37620_, _37329_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_37621_, _37620_, _37619_);
  and (_37622_, _37621_, _37618_);
  nor (_37623_, _37622_, _37321_);
  and (_37624_, _37321_, ABINPUT[9]);
  nor (_37625_, _37624_, _37623_);
  not (_37626_, _37625_);
  and (_37627_, _37626_, _37339_);
  not (_37628_, _23939_);
  and (_37629_, _37628_, _37303_);
  nor (_37630_, _37629_, _37627_);
  and (_37631_, _37630_, _37615_);
  and (_37632_, _37631_, _37356_);
  nor (_37633_, _37553_, _37356_);
  nor (_37634_, _37633_, _37632_);
  not (_37635_, _37516_);
  or (_37636_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_37637_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_37638_, _37637_, _37636_);
  or (_37639_, _37638_, _37635_);
  and (_37640_, _37639_, _37634_);
  and (_37641_, _37640_, _37597_);
  and (_37642_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_37643_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_37644_, _37643_, _37635_);
  or (_37645_, _37644_, _37642_);
  not (_37646_, _37634_);
  and (_37647_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_37648_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_37649_, _37648_, _37516_);
  or (_37650_, _37649_, _37647_);
  and (_37651_, _37650_, _37646_);
  and (_37652_, _37651_, _37645_);
  or (_37653_, _37652_, _37641_);
  and (_37654_, _37653_, _37435_);
  not (_37655_, _37307_);
  and (_37656_, _16372_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_37657_, _37656_, _16557_);
  nor (_37658_, _17004_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_37659_, _37658_, _37657_);
  not (_37660_, _37659_);
  and (_37661_, _37660_, _37592_);
  nor (_37662_, _37661_, _37655_);
  and (_37663_, _37656_, _26126_);
  nor (_37664_, _16873_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_37665_, _37664_, _37663_);
  not (_37666_, _37665_);
  and (_37667_, _37666_, _37434_);
  nor (_37668_, _37660_, _37592_);
  nor (_37669_, _37668_, _37667_);
  and (_37670_, _37669_, _37662_);
  and (_37671_, _37656_, _32583_);
  nor (_37672_, _17123_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_37673_, _37672_, _37671_);
  nand (_37674_, _37673_, _37516_);
  or (_37675_, _37673_, _37516_);
  and (_37676_, _37675_, _37674_);
  not (_37677_, _37676_);
  nor (_37678_, _37666_, _37434_);
  not (_37679_, _37678_);
  nor (_37680_, _37656_, _16557_);
  and (_37681_, _37656_, _16198_);
  nor (_37682_, _37681_, _37680_);
  not (_37683_, _37682_);
  and (_37684_, _37683_, _37634_);
  nor (_37685_, _37683_, _37634_);
  nor (_37686_, _37685_, _37684_);
  and (_37687_, _37686_, _37679_);
  and (_37688_, _37687_, _37677_);
  and (_37689_, _37688_, _37670_);
  or (_37690_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_37691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_37692_, _37592_, _37691_);
  and (_37693_, _37692_, _37690_);
  or (_37694_, _37693_, _37516_);
  and (_37695_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  not (_37696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_37697_, _37592_, _37696_);
  or (_37698_, _37697_, _37695_);
  or (_37699_, _37698_, _37635_);
  and (_37700_, _37699_, _37634_);
  and (_37701_, _37700_, _37694_);
  and (_37702_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_37703_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_37704_, _37703_, _37635_);
  or (_37705_, _37704_, _37702_);
  not (_37706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_37707_, _37592_, _37706_);
  and (_37708_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_37709_, _37708_, _37516_);
  or (_37710_, _37709_, _37707_);
  and (_37711_, _37710_, _37646_);
  and (_37712_, _37711_, _37705_);
  or (_37713_, _37712_, _37701_);
  and (_37714_, _37713_, _37434_);
  or (_37715_, _37714_, _37689_);
  or (_37716_, _37715_, _37654_);
  not (_37717_, _37689_);
  or (_37718_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_37719_, _37718_, _39026_);
  and (_40145_, _37719_, _37716_);
  nor (_37720_, _37659_, _37655_);
  nor (_37721_, _37673_, _37655_);
  and (_37722_, _37721_, _37720_);
  and (_37723_, _37682_, _37307_);
  nor (_37724_, _37665_, _37655_);
  and (_37725_, _37724_, _37723_);
  and (_37726_, _37725_, _37722_);
  or (_37727_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_37728_, _37726_);
  and (_37729_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_37730_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_37731_, _37730_, _37729_);
  and (_37732_, _37731_, ABINPUT[0]);
  not (_37733_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_37734_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_37735_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_37736_, _37735_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_37737_, _37736_, _37734_);
  and (_37738_, _37729_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_37739_, _37738_);
  and (_37740_, _37739_, _37737_);
  or (_37741_, _37740_, _37733_);
  or (_37742_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[10]);
  and (_37743_, _37742_, _37741_);
  or (_37744_, _37743_, _37732_);
  and (_37745_, _37744_, _37307_);
  or (_37746_, _37745_, _37728_);
  and (_40157_, _37746_, _37727_);
  not (_37747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_37748_, _37724_, _37723_);
  nor (_37749_, _37721_, _37720_);
  and (_37750_, _37749_, _37307_);
  and (_37751_, _37750_, _37748_);
  nor (_37752_, _37751_, _37747_);
  not (_37753_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_37754_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _37753_);
  nor (_37755_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_37756_, _37755_, _37754_);
  and (_37757_, _37756_, ABINPUT[0]);
  and (_37758_, _37733_, ABINPUT[3]);
  or (_37759_, _37758_, _37757_);
  and (_37760_, _37755_, _37753_);
  nor (_37761_, _37760_, _37733_);
  nor (_37762_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_37763_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _37735_);
  nor (_37764_, _37763_, _37762_);
  and (_37765_, _37764_, _37761_);
  or (_37766_, _37765_, _37759_);
  and (_37767_, _37766_, _37307_);
  and (_37768_, _37767_, _37751_);
  or (_40438_, _37768_, _37752_);
  not (_37769_, _37751_);
  and (_37770_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37771_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_37772_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _37735_);
  nor (_37773_, _37772_, _37771_);
  not (_37774_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor (_37775_, _37774_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_37776_, _37775_, _37753_);
  nor (_37777_, _37776_, _37733_);
  and (_37778_, _37777_, _37773_);
  and (_37779_, _37775_, _37754_);
  and (_37780_, _37779_, ABINPUT[0]);
  and (_37781_, _37733_, ABINPUT[4]);
  or (_37782_, _37781_, _37780_);
  or (_37783_, _37782_, _37778_);
  and (_37784_, _37783_, _37307_);
  and (_37785_, _37784_, _37751_);
  or (_40441_, _37785_, _37770_);
  not (_37786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_37787_, _37751_, _37786_);
  nor (_37788_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nor (_37789_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _37735_);
  nor (_37790_, _37789_, _37788_);
  and (_37791_, _37774_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_37792_, _37791_, _37753_);
  nor (_37793_, _37792_, _37733_);
  and (_37794_, _37793_, _37790_);
  and (_37795_, _37754_, _37791_);
  and (_37796_, _37795_, ABINPUT[0]);
  and (_37797_, _37733_, ABINPUT[5]);
  or (_37798_, _37797_, _37796_);
  or (_37799_, _37798_, _37794_);
  and (_37800_, _37799_, _37307_);
  and (_37801_, _37800_, _37751_);
  or (_40445_, _37801_, _37787_);
  and (_37802_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_37803_, _37754_, _37729_);
  and (_37804_, _37803_, ABINPUT[0]);
  nor (_37805_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_37806_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _37735_);
  nor (_37807_, _37806_, _37805_);
  and (_37808_, _37729_, _37753_);
  not (_37809_, _37808_);
  and (_37810_, _37809_, _37807_);
  or (_37811_, _37810_, _37733_);
  or (_37812_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[6]);
  and (_37813_, _37812_, _37811_);
  or (_37814_, _37813_, _37804_);
  and (_37815_, _37814_, _37307_);
  and (_37816_, _37815_, _37751_);
  or (_40451_, _37816_, _37802_);
  not (_37817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_37818_, _37751_, _37817_);
  nor (_37819_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_37820_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _37735_);
  nor (_37821_, _37820_, _37819_);
  and (_37822_, _37755_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_37823_, _37822_, _37733_);
  and (_37824_, _37823_, _37821_);
  and (_37825_, _37755_, _37730_);
  and (_37826_, _37825_, ABINPUT[0]);
  and (_37827_, _37733_, ABINPUT[7]);
  or (_37828_, _37827_, _37826_);
  or (_37829_, _37828_, _37824_);
  and (_37830_, _37829_, _37307_);
  and (_37831_, _37830_, _37751_);
  or (_40457_, _37831_, _37818_);
  and (_37832_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_37833_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_37834_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _37735_);
  nor (_37835_, _37834_, _37833_);
  and (_37836_, _37775_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_37837_, _37836_, _37733_);
  and (_37838_, _37837_, _37835_);
  and (_37839_, _37775_, _37730_);
  and (_37840_, _37839_, ABINPUT[0]);
  and (_37841_, _37733_, ABINPUT[8]);
  or (_37842_, _37841_, _37840_);
  or (_37843_, _37842_, _37838_);
  and (_37844_, _37843_, _37307_);
  and (_37845_, _37844_, _37751_);
  or (_40463_, _37845_, _37832_);
  not (_37846_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_37847_, _37751_, _37846_);
  nor (_37848_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_37849_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _37735_);
  nor (_37850_, _37849_, _37848_);
  and (_37851_, _37791_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_37852_, _37851_, _37733_);
  and (_37853_, _37852_, _37850_);
  and (_37854_, _37791_, _37730_);
  and (_37855_, _37854_, ABINPUT[0]);
  and (_37856_, _37733_, ABINPUT[9]);
  or (_37857_, _37856_, _37855_);
  or (_37858_, _37857_, _37853_);
  and (_37859_, _37858_, _37307_);
  and (_37860_, _37859_, _37751_);
  or (_40469_, _37860_, _37847_);
  and (_37861_, _37769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_37862_, _37751_, _37745_);
  or (_40472_, _37862_, _37861_);
  not (_37863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_37864_, _37720_, _37673_);
  and (_37865_, _37864_, _37748_);
  nor (_37866_, _37865_, _37863_);
  and (_37867_, _37865_, _37767_);
  or (_40480_, _37867_, _37866_);
  or (_37868_, _37865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  not (_37869_, _37865_);
  or (_37870_, _37869_, _37784_);
  and (_40484_, _37870_, _37868_);
  not (_37871_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_37872_, _37865_, _37871_);
  and (_37873_, _37865_, _37800_);
  or (_40488_, _37873_, _37872_);
  not (_37874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_37875_, _37865_, _37874_);
  and (_37876_, _37865_, _37815_);
  or (_40492_, _37876_, _37875_);
  not (_37877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_37878_, _37865_, _37877_);
  and (_37879_, _37865_, _37830_);
  or (_40496_, _37879_, _37878_);
  not (_37880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_37881_, _37865_, _37880_);
  and (_37882_, _37865_, _37844_);
  or (_40500_, _37882_, _37881_);
  not (_37883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_37884_, _37865_, _37883_);
  and (_37885_, _37865_, _37859_);
  or (_40504_, _37885_, _37884_);
  or (_37886_, _37865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_37887_, _37869_, _37745_);
  and (_40507_, _37887_, _37886_);
  not (_37888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_37889_, _37721_, _37659_);
  and (_37890_, _37889_, _37748_);
  nor (_37891_, _37890_, _37888_);
  and (_37892_, _37890_, _37767_);
  or (_40515_, _37892_, _37891_);
  or (_37893_, _37890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  not (_37894_, _37890_);
  or (_37895_, _37894_, _37784_);
  and (_40519_, _37895_, _37893_);
  not (_37896_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_37897_, _37890_, _37896_);
  and (_37898_, _37890_, _37800_);
  or (_40523_, _37898_, _37897_);
  or (_37899_, _37890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_37900_, _37894_, _37815_);
  and (_40527_, _37900_, _37899_);
  not (_37901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_37902_, _37890_, _37901_);
  and (_37903_, _37890_, _37830_);
  or (_40531_, _37903_, _37902_);
  or (_37904_, _37890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_37905_, _37894_, _37844_);
  and (_40535_, _37905_, _37904_);
  not (_37906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_37907_, _37890_, _37906_);
  and (_37908_, _37890_, _37859_);
  or (_40539_, _37908_, _37907_);
  or (_37909_, _37890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_37910_, _37894_, _37745_);
  and (_40542_, _37910_, _37909_);
  not (_37911_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_37912_, _37748_, _37722_);
  nor (_37913_, _37912_, _37911_);
  and (_37914_, _37912_, _37767_);
  or (_40548_, _37914_, _37913_);
  or (_37915_, _37912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  not (_37916_, _37912_);
  or (_37917_, _37916_, _37784_);
  and (_40552_, _37917_, _37915_);
  not (_37918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_37919_, _37912_, _37918_);
  and (_37920_, _37912_, _37800_);
  or (_40556_, _37920_, _37919_);
  not (_37921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_37922_, _37912_, _37921_);
  and (_37923_, _37912_, _37815_);
  or (_40560_, _37923_, _37922_);
  not (_37924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_37925_, _37912_, _37924_);
  and (_37926_, _37912_, _37830_);
  or (_40564_, _37926_, _37925_);
  or (_37927_, _37912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_37928_, _37916_, _37844_);
  and (_40568_, _37928_, _37927_);
  not (_37929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_37930_, _37912_, _37929_);
  and (_37931_, _37912_, _37859_);
  or (_40572_, _37931_, _37930_);
  nor (_37932_, _37912_, _37706_);
  and (_37933_, _37912_, _37745_);
  or (_40574_, _37933_, _37932_);
  not (_37934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_37935_, _37724_, _37683_);
  and (_37936_, _37935_, _37749_);
  nor (_37937_, _37936_, _37934_);
  and (_37938_, _37936_, _37767_);
  or (_40580_, _37938_, _37937_);
  or (_37939_, _37936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  not (_37940_, _37936_);
  or (_37941_, _37940_, _37784_);
  and (_40584_, _37941_, _37939_);
  not (_37942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_37943_, _37936_, _37942_);
  and (_37944_, _37936_, _37800_);
  or (_40588_, _37944_, _37943_);
  and (_37945_, _37940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_37946_, _37936_, _37815_);
  or (_40592_, _37946_, _37945_);
  not (_37947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_37948_, _37936_, _37947_);
  and (_37949_, _37936_, _37830_);
  or (_40596_, _37949_, _37948_);
  and (_37950_, _37940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_37951_, _37936_, _37844_);
  or (_40600_, _37951_, _37950_);
  not (_37952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_37953_, _37936_, _37952_);
  and (_37954_, _37936_, _37859_);
  or (_40604_, _37954_, _37953_);
  and (_37955_, _37940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_37956_, _37936_, _37745_);
  or (_40607_, _37956_, _37955_);
  not (_37957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_37958_, _37935_, _37864_);
  nor (_37959_, _37958_, _37957_);
  and (_37960_, _37958_, _37767_);
  or (_40612_, _37960_, _37959_);
  or (_37961_, _37958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  not (_37962_, _37958_);
  or (_37963_, _37962_, _37784_);
  and (_40616_, _37963_, _37961_);
  not (_37964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_37965_, _37958_, _37964_);
  and (_37966_, _37958_, _37800_);
  or (_40620_, _37966_, _37965_);
  or (_37967_, _37958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_37968_, _37962_, _37815_);
  and (_40624_, _37968_, _37967_);
  not (_37969_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_37970_, _37958_, _37969_);
  and (_37971_, _37958_, _37830_);
  or (_40628_, _37971_, _37970_);
  not (_37972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_37973_, _37958_, _37972_);
  and (_37974_, _37958_, _37844_);
  or (_40632_, _37974_, _37973_);
  not (_37975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_37976_, _37958_, _37975_);
  and (_37977_, _37958_, _37859_);
  or (_40636_, _37977_, _37976_);
  or (_37978_, _37958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_37979_, _37962_, _37745_);
  and (_40639_, _37979_, _37978_);
  not (_37980_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_37981_, _37935_, _37889_);
  nor (_37982_, _37981_, _37980_);
  and (_37983_, _37981_, _37767_);
  or (_40644_, _37983_, _37982_);
  or (_37984_, _37981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  not (_37985_, _37981_);
  or (_37986_, _37985_, _37784_);
  and (_40648_, _37986_, _37984_);
  not (_37987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_37988_, _37981_, _37987_);
  and (_37989_, _37981_, _37800_);
  or (_40652_, _37989_, _37988_);
  or (_37990_, _37981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_37991_, _37985_, _37815_);
  and (_40656_, _37991_, _37990_);
  not (_37992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_37993_, _37981_, _37992_);
  and (_37994_, _37981_, _37830_);
  or (_40660_, _37994_, _37993_);
  and (_37995_, _37985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_37996_, _37981_, _37844_);
  or (_40664_, _37996_, _37995_);
  not (_37997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_37998_, _37981_, _37997_);
  and (_37999_, _37981_, _37859_);
  or (_40668_, _37999_, _37998_);
  and (_38000_, _37985_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_38001_, _37981_, _37745_);
  or (_40671_, _38001_, _38000_);
  not (_38002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_38003_, _37935_, _37722_);
  nor (_38004_, _38003_, _38002_);
  and (_38005_, _38003_, _37767_);
  or (_40676_, _38005_, _38004_);
  or (_38006_, _38003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  not (_38007_, _38003_);
  or (_38008_, _38007_, _37784_);
  and (_40680_, _38008_, _38006_);
  not (_38009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_38010_, _38003_, _38009_);
  and (_38011_, _38003_, _37800_);
  or (_40684_, _38011_, _38010_);
  or (_38012_, _38003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_38013_, _38007_, _37815_);
  and (_40688_, _38013_, _38012_);
  not (_38014_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_38015_, _38003_, _38014_);
  and (_38016_, _38003_, _37830_);
  or (_40692_, _38016_, _38015_);
  not (_38017_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_38018_, _38003_, _38017_);
  and (_38019_, _38003_, _37844_);
  or (_40696_, _38019_, _38018_);
  not (_38020_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_38021_, _38003_, _38020_);
  and (_38022_, _38003_, _37859_);
  or (_40700_, _38022_, _38021_);
  or (_38023_, _38003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_38024_, _38007_, _37745_);
  and (_40703_, _38024_, _38023_);
  not (_38025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_38026_, _37723_, _37665_);
  and (_38027_, _38026_, _37749_);
  nor (_38028_, _38027_, _38025_);
  and (_38029_, _38027_, _37767_);
  or (_40711_, _38029_, _38028_);
  or (_38030_, _38027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  not (_38031_, _38027_);
  or (_38032_, _38031_, _37784_);
  and (_40715_, _38032_, _38030_);
  not (_38033_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_38034_, _38027_, _38033_);
  and (_38035_, _38027_, _37800_);
  or (_40719_, _38035_, _38034_);
  not (_38036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_38037_, _38027_, _38036_);
  and (_38038_, _38027_, _37815_);
  or (_40723_, _38038_, _38037_);
  not (_38039_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_38040_, _38027_, _38039_);
  and (_38041_, _38027_, _37830_);
  or (_40727_, _38041_, _38040_);
  not (_38042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_38043_, _38027_, _38042_);
  and (_38044_, _38027_, _37844_);
  or (_40731_, _38044_, _38043_);
  not (_38045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_38046_, _38027_, _38045_);
  and (_38047_, _38027_, _37859_);
  or (_40735_, _38047_, _38046_);
  or (_38048_, _38027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_38049_, _38031_, _37745_);
  and (_40738_, _38049_, _38048_);
  not (_38050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_38051_, _38026_, _37864_);
  nor (_38052_, _38051_, _38050_);
  and (_38053_, _38051_, _37767_);
  or (_40743_, _38053_, _38052_);
  or (_38054_, _38051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  not (_38055_, _38051_);
  or (_38056_, _38055_, _37784_);
  and (_40747_, _38056_, _38054_);
  not (_38057_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_38058_, _38051_, _38057_);
  and (_38059_, _38051_, _37800_);
  or (_40751_, _38059_, _38058_);
  or (_38060_, _38051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_38061_, _38055_, _37815_);
  and (_40755_, _38061_, _38060_);
  not (_38062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_38063_, _38051_, _38062_);
  and (_38064_, _38051_, _37830_);
  or (_40759_, _38064_, _38063_);
  or (_38065_, _38051_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_38066_, _38055_, _37844_);
  and (_40763_, _38066_, _38065_);
  not (_38067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_38068_, _38051_, _38067_);
  and (_38069_, _38051_, _37859_);
  or (_40767_, _38069_, _38068_);
  nor (_38070_, _38051_, _37696_);
  and (_38071_, _38051_, _37745_);
  or (_40770_, _38071_, _38070_);
  not (_38072_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_38073_, _38026_, _37889_);
  nor (_38074_, _38073_, _38072_);
  and (_38075_, _38073_, _37767_);
  or (_40775_, _38075_, _38074_);
  not (_38076_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_38078_, _38073_, _38076_);
  and (_38079_, _38073_, _37784_);
  or (_40779_, _38079_, _38078_);
  not (_38080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_38081_, _38073_, _38080_);
  and (_38082_, _38073_, _37800_);
  or (_40783_, _38082_, _38081_);
  not (_38083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_38084_, _38073_, _38083_);
  and (_38085_, _38073_, _37815_);
  or (_40787_, _38085_, _38084_);
  not (_38087_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_38088_, _38073_, _38087_);
  and (_38089_, _38073_, _37830_);
  or (_40791_, _38089_, _38088_);
  or (_38090_, _38073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  not (_38091_, _38073_);
  or (_38092_, _38091_, _37844_);
  and (_40795_, _38092_, _38090_);
  not (_38093_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_38095_, _38073_, _38093_);
  and (_38096_, _38073_, _37859_);
  or (_40799_, _38096_, _38095_);
  nor (_38097_, _38073_, _37691_);
  and (_38098_, _38073_, _37745_);
  or (_40801_, _38098_, _38097_);
  not (_38099_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_38100_, _38026_, _37722_);
  nor (_38101_, _38100_, _38099_);
  and (_38102_, _38100_, _37767_);
  or (_40806_, _38102_, _38101_);
  not (_38104_, _38100_);
  and (_38105_, _38104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_38106_, _38100_, _37784_);
  or (_40810_, _38106_, _38105_);
  not (_38107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_38108_, _38100_, _38107_);
  and (_38109_, _38100_, _37800_);
  or (_40814_, _38109_, _38108_);
  and (_38110_, _38104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_38112_, _38100_, _37815_);
  or (_40818_, _38112_, _38110_);
  not (_38113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_38114_, _38100_, _38113_);
  and (_38115_, _38100_, _37830_);
  or (_40822_, _38115_, _38114_);
  or (_38116_, _38100_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_38117_, _38104_, _37844_);
  and (_40826_, _38117_, _38116_);
  not (_38118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_38120_, _38100_, _38118_);
  and (_38121_, _38100_, _37859_);
  or (_40830_, _38121_, _38120_);
  and (_38122_, _38104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_38123_, _38100_, _37745_);
  or (_40833_, _38123_, _38122_);
  not (_38124_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_38125_, _37749_, _37725_);
  nor (_38126_, _38125_, _38124_);
  and (_38127_, _38125_, _37767_);
  or (_40839_, _38127_, _38126_);
  not (_38129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_38130_, _38125_, _38129_);
  and (_38131_, _38125_, _37784_);
  or (_40843_, _38131_, _38130_);
  not (_38132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_38133_, _38125_, _38132_);
  and (_38134_, _38125_, _37800_);
  or (_40847_, _38134_, _38133_);
  not (_38135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_38136_, _38125_, _38135_);
  and (_38137_, _38125_, _37815_);
  or (_40851_, _38137_, _38136_);
  not (_38138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_38139_, _38125_, _38138_);
  and (_38140_, _38125_, _37830_);
  or (_40855_, _38140_, _38139_);
  not (_38141_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_38142_, _38125_, _38141_);
  and (_38143_, _38125_, _37844_);
  or (_40859_, _38143_, _38142_);
  not (_38144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_38145_, _38125_, _38144_);
  and (_38146_, _38125_, _37859_);
  or (_40863_, _38146_, _38145_);
  or (_38147_, _38125_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  not (_38148_, _38125_);
  or (_38149_, _38148_, _37745_);
  and (_40866_, _38149_, _38147_);
  not (_38150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_38151_, _37864_, _37725_);
  nor (_38152_, _38151_, _38150_);
  and (_38153_, _38151_, _37767_);
  or (_40871_, _38153_, _38152_);
  or (_38154_, _38151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  not (_38155_, _38151_);
  or (_38156_, _38155_, _37784_);
  and (_40875_, _38156_, _38154_);
  not (_38157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_38158_, _38151_, _38157_);
  and (_38159_, _38151_, _37800_);
  or (_40879_, _38159_, _38158_);
  or (_38160_, _38151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_38161_, _38155_, _37815_);
  and (_40883_, _38161_, _38160_);
  not (_38162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_38163_, _38151_, _38162_);
  and (_38164_, _38151_, _37830_);
  or (_40887_, _38164_, _38163_);
  or (_38165_, _38151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_38166_, _38155_, _37844_);
  and (_40891_, _38166_, _38165_);
  not (_38167_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_38168_, _38151_, _38167_);
  and (_38169_, _38151_, _37859_);
  or (_40895_, _38169_, _38168_);
  or (_38170_, _38151_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_38171_, _38155_, _37745_);
  and (_40898_, _38171_, _38170_);
  not (_38172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_38173_, _37889_, _37725_);
  nor (_38174_, _38173_, _38172_);
  and (_38175_, _38173_, _37767_);
  or (_40903_, _38175_, _38174_);
  or (_38176_, _38173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  not (_38177_, _38173_);
  or (_38178_, _38177_, _37784_);
  and (_40907_, _38178_, _38176_);
  not (_38179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_38180_, _38173_, _38179_);
  and (_38181_, _38173_, _37800_);
  or (_40911_, _38181_, _38180_);
  or (_38182_, _38173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_38183_, _38177_, _37815_);
  and (_40915_, _38183_, _38182_);
  not (_38184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_38185_, _38173_, _38184_);
  and (_38186_, _38173_, _37830_);
  or (_40919_, _38186_, _38185_);
  or (_38187_, _38173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_38188_, _38177_, _37844_);
  and (_40923_, _38188_, _38187_);
  not (_38189_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_38190_, _38173_, _38189_);
  and (_38191_, _38173_, _37859_);
  or (_40927_, _38191_, _38190_);
  or (_38192_, _38173_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_38193_, _38177_, _37745_);
  and (_40930_, _38193_, _38192_);
  not (_38194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_38195_, _37726_, _38194_);
  and (_38196_, _37767_, _37726_);
  or (_40935_, _38196_, _38195_);
  or (_38197_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_38198_, _37784_, _37728_);
  and (_40939_, _38198_, _38197_);
  not (_38199_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_38200_, _37726_, _38199_);
  and (_38201_, _37800_, _37726_);
  or (_40943_, _38201_, _38200_);
  or (_38202_, _37726_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_38203_, _37815_, _37728_);
  and (_40947_, _38203_, _38202_);
  not (_38204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_38205_, _37726_, _38204_);
  and (_38206_, _37830_, _37726_);
  or (_40951_, _38206_, _38205_);
  not (_38207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_38208_, _37726_, _38207_);
  and (_38209_, _37844_, _37726_);
  or (_40955_, _38209_, _38208_);
  not (_38210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_38211_, _37726_, _38210_);
  and (_38212_, _37859_, _37726_);
  or (_40959_, _38212_, _38211_);
  and (_38213_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_38214_, _37592_, _37863_);
  or (_38215_, _38214_, _38213_);
  and (_38216_, _38215_, _37516_);
  nor (_38217_, _37592_, _37911_);
  and (_38218_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_38219_, _38218_, _38217_);
  and (_38220_, _38219_, _37635_);
  or (_38221_, _38220_, _38216_);
  or (_38222_, _38221_, _37435_);
  and (_38223_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_38224_, _37592_, _37957_);
  or (_38225_, _38224_, _38223_);
  and (_38226_, _38225_, _37516_);
  nor (_38227_, _37592_, _38002_);
  and (_38228_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_38229_, _38228_, _38227_);
  and (_38230_, _38229_, _37635_);
  or (_38231_, _38230_, _38226_);
  or (_38232_, _38231_, _37434_);
  and (_38233_, _38232_, _37646_);
  and (_38234_, _38233_, _38222_);
  nand (_38235_, _37592_, _38025_);
  or (_38236_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_38237_, _38236_, _38235_);
  and (_38238_, _38237_, _37516_);
  or (_38239_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_38240_, _37592_, _38072_);
  and (_38241_, _38240_, _38239_);
  and (_38242_, _38241_, _37635_);
  or (_38243_, _38242_, _38238_);
  or (_38244_, _38243_, _37435_);
  nand (_38245_, _37592_, _38124_);
  or (_38246_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_38247_, _38246_, _38245_);
  and (_38248_, _38247_, _37516_);
  or (_38249_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_38250_, _37592_, _38172_);
  and (_38251_, _38250_, _38249_);
  and (_38252_, _38251_, _37635_);
  or (_38253_, _38252_, _38248_);
  or (_38254_, _38253_, _37434_);
  and (_38255_, _38254_, _37634_);
  and (_38256_, _38255_, _38244_);
  or (_38257_, _38256_, _38234_);
  or (_38258_, _38257_, _37689_);
  or (_38259_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_38260_, _38259_, _39026_);
  and (_00048_, _38260_, _38258_);
  and (_38261_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_38262_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_38263_, _38262_, _38261_);
  and (_38264_, _38263_, _37516_);
  and (_38265_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_38266_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_38267_, _38266_, _38265_);
  and (_38268_, _38267_, _37635_);
  or (_38269_, _38268_, _38264_);
  or (_38270_, _38269_, _37435_);
  and (_38271_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_38272_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_38273_, _38272_, _38271_);
  and (_38274_, _38273_, _37516_);
  and (_38275_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_38276_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_38277_, _38276_, _38275_);
  and (_38278_, _38277_, _37635_);
  or (_38279_, _38278_, _38274_);
  or (_38280_, _38279_, _37434_);
  and (_38281_, _38280_, _37646_);
  and (_38282_, _38281_, _38270_);
  or (_38283_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_38284_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_38285_, _38284_, _38283_);
  and (_38286_, _38285_, _37516_);
  or (_38287_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand (_38288_, _37592_, _38076_);
  and (_38289_, _38288_, _38287_);
  and (_38291_, _38289_, _37635_);
  or (_38293_, _38291_, _38286_);
  or (_38295_, _38293_, _37435_);
  nand (_38297_, _37592_, _38129_);
  or (_38299_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_38301_, _38299_, _38297_);
  and (_38303_, _38301_, _37516_);
  or (_38305_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_38307_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_38309_, _38307_, _38305_);
  and (_38311_, _38309_, _37635_);
  or (_38313_, _38311_, _38303_);
  or (_38315_, _38313_, _37434_);
  and (_38317_, _38315_, _37634_);
  and (_38319_, _38317_, _38295_);
  or (_38321_, _38319_, _38282_);
  or (_38323_, _38321_, _37689_);
  or (_38325_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_38327_, _38325_, _39026_);
  and (_00050_, _38327_, _38323_);
  and (_38330_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_38332_, _37592_, _37871_);
  or (_38334_, _38332_, _38330_);
  and (_38336_, _38334_, _37516_);
  nor (_38338_, _37592_, _37918_);
  and (_38340_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_38342_, _38340_, _38338_);
  and (_38344_, _38342_, _37635_);
  or (_38345_, _38344_, _38336_);
  or (_38346_, _38345_, _37435_);
  and (_38347_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_38348_, _37592_, _37964_);
  or (_38349_, _38348_, _38347_);
  and (_38350_, _38349_, _37516_);
  nor (_38351_, _37592_, _38009_);
  and (_38352_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_38353_, _38352_, _38351_);
  and (_38354_, _38353_, _37635_);
  or (_38355_, _38354_, _38350_);
  or (_38356_, _38355_, _37434_);
  and (_38357_, _38356_, _37646_);
  and (_38358_, _38357_, _38346_);
  nand (_38359_, _37592_, _38033_);
  or (_38360_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_38361_, _38360_, _38359_);
  and (_38362_, _38361_, _37516_);
  or (_38363_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_38364_, _37592_, _38080_);
  and (_38365_, _38364_, _38363_);
  and (_38366_, _38365_, _37635_);
  or (_38367_, _38366_, _38362_);
  or (_38368_, _38367_, _37435_);
  nand (_38369_, _37592_, _38132_);
  or (_38370_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_38371_, _38370_, _38369_);
  and (_38372_, _38371_, _37516_);
  or (_38373_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_38374_, _37592_, _38179_);
  and (_38375_, _38374_, _38373_);
  and (_38376_, _38375_, _37635_);
  or (_38377_, _38376_, _38372_);
  or (_38378_, _38377_, _37434_);
  and (_38379_, _38378_, _37634_);
  and (_38380_, _38379_, _38368_);
  or (_38381_, _38380_, _38358_);
  or (_38382_, _38381_, _37689_);
  or (_38383_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_38384_, _38383_, _39026_);
  and (_00052_, _38384_, _38382_);
  or (_38385_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_38386_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_38387_, _38386_, _38385_);
  or (_38388_, _38387_, _37516_);
  nand (_38389_, _37592_, _38135_);
  or (_38390_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_38391_, _38390_, _38389_);
  or (_38392_, _38391_, _37635_);
  and (_38393_, _38392_, _37634_);
  and (_38394_, _38393_, _38388_);
  and (_38395_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_38396_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_38397_, _38396_, _37635_);
  or (_38398_, _38397_, _38395_);
  and (_38399_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_38400_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_38401_, _38400_, _37516_);
  or (_38402_, _38401_, _38399_);
  and (_38403_, _38402_, _37646_);
  and (_38404_, _38403_, _38398_);
  or (_38405_, _38404_, _38394_);
  and (_38406_, _38405_, _37435_);
  or (_38407_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand (_38408_, _37592_, _38083_);
  and (_38409_, _38408_, _38407_);
  or (_38410_, _38409_, _37516_);
  nand (_38411_, _37592_, _38036_);
  or (_38412_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_38413_, _38412_, _38411_);
  or (_38414_, _38413_, _37635_);
  and (_38415_, _38414_, _37634_);
  and (_38416_, _38415_, _38410_);
  and (_38417_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_38418_, _37592_, _37874_);
  or (_38419_, _38418_, _37635_);
  or (_38420_, _38419_, _38417_);
  nor (_38421_, _37592_, _37921_);
  and (_38422_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_38423_, _38422_, _37516_);
  or (_38424_, _38423_, _38421_);
  and (_38425_, _38424_, _37646_);
  and (_38426_, _38425_, _38420_);
  or (_38427_, _38426_, _38416_);
  and (_38428_, _38427_, _37434_);
  or (_38429_, _38428_, _37689_);
  or (_38430_, _38429_, _38406_);
  or (_38431_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_38432_, _38431_, _39026_);
  and (_00053_, _38432_, _38430_);
  and (_38433_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_38434_, _37592_, _37877_);
  or (_38435_, _38434_, _38433_);
  and (_38436_, _38435_, _37516_);
  nor (_38437_, _37592_, _37924_);
  and (_38438_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_38439_, _38438_, _38437_);
  and (_38440_, _38439_, _37635_);
  or (_38441_, _38440_, _38436_);
  or (_38442_, _38441_, _37435_);
  and (_38443_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_38444_, _37592_, _37969_);
  or (_38445_, _38444_, _38443_);
  and (_38446_, _38445_, _37516_);
  nor (_38447_, _37592_, _38014_);
  and (_38448_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_38449_, _38448_, _38447_);
  and (_38450_, _38449_, _37635_);
  or (_38451_, _38450_, _38446_);
  or (_38452_, _38451_, _37434_);
  and (_38453_, _38452_, _37646_);
  and (_38454_, _38453_, _38442_);
  nand (_38455_, _37592_, _38039_);
  or (_38456_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_38457_, _38456_, _38455_);
  and (_38458_, _38457_, _37516_);
  or (_38459_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_38460_, _37592_, _38087_);
  and (_38461_, _38460_, _38459_);
  and (_38462_, _38461_, _37635_);
  or (_38463_, _38462_, _38458_);
  or (_38464_, _38463_, _37435_);
  nand (_38465_, _37592_, _38138_);
  or (_38466_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_38467_, _38466_, _38465_);
  and (_38468_, _38467_, _37516_);
  or (_38469_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_38470_, _37592_, _38184_);
  and (_38471_, _38470_, _38469_);
  and (_38472_, _38471_, _37635_);
  or (_38473_, _38472_, _38468_);
  or (_38474_, _38473_, _37434_);
  and (_38475_, _38474_, _37634_);
  and (_38476_, _38475_, _38464_);
  or (_38477_, _38476_, _38454_);
  or (_38478_, _38477_, _37689_);
  or (_38479_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_38480_, _38479_, _39026_);
  and (_00055_, _38480_, _38478_);
  and (_38481_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_38482_, _37592_, _37880_);
  or (_38483_, _38482_, _38481_);
  and (_38484_, _38483_, _37516_);
  and (_38485_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_38486_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_38487_, _38486_, _38485_);
  and (_38488_, _38487_, _37635_);
  or (_38489_, _38488_, _38484_);
  or (_38490_, _38489_, _37435_);
  and (_38491_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_38492_, _37592_, _37972_);
  or (_38493_, _38492_, _38491_);
  and (_38494_, _38493_, _37516_);
  nor (_38495_, _37592_, _38017_);
  and (_38496_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_38497_, _38496_, _38495_);
  and (_38498_, _38497_, _37635_);
  or (_38499_, _38498_, _38494_);
  or (_38500_, _38499_, _37434_);
  and (_38501_, _38500_, _37646_);
  and (_38502_, _38501_, _38490_);
  nand (_38503_, _37592_, _38042_);
  or (_38504_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_38505_, _38504_, _38503_);
  and (_38506_, _38505_, _37516_);
  or (_38507_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_38508_, _37594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_38509_, _38508_, _38507_);
  and (_38510_, _38509_, _37635_);
  or (_38511_, _38510_, _38506_);
  or (_38512_, _38511_, _37435_);
  nand (_38513_, _37592_, _38141_);
  or (_38514_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_38515_, _38514_, _38513_);
  and (_38516_, _38515_, _37516_);
  and (_38517_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_38518_, _37592_, _38207_);
  or (_38519_, _38518_, _38517_);
  and (_38520_, _38519_, _37635_);
  or (_38521_, _38520_, _38516_);
  or (_38522_, _38521_, _37434_);
  and (_38523_, _38522_, _37634_);
  and (_38524_, _38523_, _38512_);
  or (_38525_, _38524_, _38502_);
  or (_38526_, _38525_, _37689_);
  or (_38527_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_38528_, _38527_, _39026_);
  and (_00057_, _38528_, _38526_);
  and (_38529_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_38530_, _37592_, _37883_);
  or (_38531_, _38530_, _38529_);
  and (_38532_, _38531_, _37516_);
  nor (_38533_, _37592_, _37929_);
  and (_38534_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_38535_, _38534_, _38533_);
  and (_38536_, _38535_, _37635_);
  or (_38537_, _38536_, _38532_);
  or (_38538_, _38537_, _37435_);
  and (_38539_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_38540_, _37592_, _37975_);
  or (_38541_, _38540_, _38539_);
  and (_38542_, _38541_, _37516_);
  nor (_38543_, _37592_, _38020_);
  and (_38544_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_38545_, _38544_, _38543_);
  and (_38546_, _38545_, _37635_);
  or (_38547_, _38546_, _38542_);
  or (_38548_, _38547_, _37434_);
  and (_38549_, _38548_, _37646_);
  and (_38550_, _38549_, _38538_);
  nand (_38551_, _37592_, _38045_);
  or (_38552_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_38553_, _38552_, _38551_);
  and (_38554_, _38553_, _37516_);
  or (_38555_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_38556_, _37592_, _38093_);
  and (_38557_, _38556_, _38555_);
  and (_38558_, _38557_, _37635_);
  or (_38559_, _38558_, _38554_);
  or (_38560_, _38559_, _37435_);
  nand (_38561_, _37592_, _38144_);
  or (_38562_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_38563_, _38562_, _38561_);
  and (_38564_, _38563_, _37516_);
  or (_38565_, _37592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_38566_, _37592_, _38189_);
  and (_38567_, _38566_, _38565_);
  and (_38568_, _38567_, _37635_);
  or (_38569_, _38568_, _38564_);
  or (_38570_, _38569_, _37434_);
  and (_38571_, _38570_, _37634_);
  and (_38572_, _38571_, _38560_);
  or (_38573_, _38572_, _38550_);
  or (_38574_, _38573_, _37689_);
  or (_38575_, _37717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_38576_, _38575_, _39026_);
  and (_00059_, _38576_, _38574_);
  or (_38577_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_38578_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_38579_, _38578_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_38580_, _38579_, _38577_);
  nand (_38585_, _38580_, _39026_);
  or (_38591_, \oc8051_gm_cxrom_1.cell0.data [7], _39026_);
  and (_00067_, _38591_, _38585_);
  or (_38602_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38608_, \oc8051_gm_cxrom_1.cell0.data [0], _38578_);
  nand (_38612_, _38608_, _38602_);
  nand (_38613_, _38612_, _39026_);
  or (_38614_, \oc8051_gm_cxrom_1.cell0.data [0], _39026_);
  and (_00098_, _38614_, _38613_);
  or (_38615_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38616_, \oc8051_gm_cxrom_1.cell0.data [1], _38578_);
  nand (_38617_, _38616_, _38615_);
  nand (_38618_, _38617_, _39026_);
  or (_38619_, \oc8051_gm_cxrom_1.cell0.data [1], _39026_);
  and (_00100_, _38619_, _38618_);
  or (_38620_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38621_, \oc8051_gm_cxrom_1.cell0.data [2], _38578_);
  nand (_38622_, _38621_, _38620_);
  nand (_38623_, _38622_, _39026_);
  or (_38624_, \oc8051_gm_cxrom_1.cell0.data [2], _39026_);
  and (_00102_, _38624_, _38623_);
  or (_38625_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38626_, \oc8051_gm_cxrom_1.cell0.data [3], _38578_);
  nand (_38627_, _38626_, _38625_);
  nand (_38628_, _38627_, _39026_);
  or (_38629_, \oc8051_gm_cxrom_1.cell0.data [3], _39026_);
  and (_00104_, _38629_, _38628_);
  or (_38630_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38631_, \oc8051_gm_cxrom_1.cell0.data [4], _38578_);
  nand (_38632_, _38631_, _38630_);
  nand (_38633_, _38632_, _39026_);
  or (_38634_, \oc8051_gm_cxrom_1.cell0.data [4], _39026_);
  and (_00106_, _38634_, _38633_);
  or (_38635_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38636_, \oc8051_gm_cxrom_1.cell0.data [5], _38578_);
  nand (_38637_, _38636_, _38635_);
  nand (_38638_, _38637_, _39026_);
  or (_38639_, \oc8051_gm_cxrom_1.cell0.data [5], _39026_);
  and (_00108_, _38639_, _38638_);
  or (_38640_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_38641_, \oc8051_gm_cxrom_1.cell0.data [6], _38578_);
  nand (_38642_, _38641_, _38640_);
  nand (_38645_, _38642_, _39026_);
  or (_38648_, \oc8051_gm_cxrom_1.cell0.data [6], _39026_);
  and (_00110_, _38648_, _38645_);
  or (_38653_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_38654_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_38655_, _38654_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_38659_, _38655_, _38653_);
  nand (_38665_, _38659_, _39026_);
  or (_38666_, \oc8051_gm_cxrom_1.cell1.data [7], _39026_);
  and (_00117_, _38666_, _38665_);
  or (_38667_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38673_, \oc8051_gm_cxrom_1.cell1.data [0], _38654_);
  nand (_38677_, _38673_, _38667_);
  nand (_38678_, _38677_, _39026_);
  or (_38679_, \oc8051_gm_cxrom_1.cell1.data [0], _39026_);
  and (_00150_, _38679_, _38678_);
  or (_38688_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38689_, \oc8051_gm_cxrom_1.cell1.data [1], _38654_);
  nand (_38690_, _38689_, _38688_);
  nand (_38691_, _38690_, _39026_);
  or (_38697_, \oc8051_gm_cxrom_1.cell1.data [1], _39026_);
  and (_00152_, _38697_, _38691_);
  or (_38701_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38702_, \oc8051_gm_cxrom_1.cell1.data [2], _38654_);
  nand (_38707_, _38702_, _38701_);
  nand (_38712_, _38707_, _39026_);
  or (_38713_, \oc8051_gm_cxrom_1.cell1.data [2], _39026_);
  and (_00154_, _38713_, _38712_);
  or (_38718_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38723_, \oc8051_gm_cxrom_1.cell1.data [3], _38654_);
  nand (_38724_, _38723_, _38718_);
  nand (_38725_, _38724_, _39026_);
  or (_38729_, \oc8051_gm_cxrom_1.cell1.data [3], _39026_);
  and (_00156_, _38729_, _38725_);
  or (_38735_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38736_, \oc8051_gm_cxrom_1.cell1.data [4], _38654_);
  nand (_38737_, _38736_, _38735_);
  nand (_38743_, _38737_, _39026_);
  or (_38747_, \oc8051_gm_cxrom_1.cell1.data [4], _39026_);
  and (_00158_, _38747_, _38743_);
  or (_38748_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38753_, \oc8051_gm_cxrom_1.cell1.data [5], _38654_);
  nand (_38758_, _38753_, _38748_);
  nand (_38759_, _38758_, _39026_);
  or (_38760_, \oc8051_gm_cxrom_1.cell1.data [5], _39026_);
  and (_00160_, _38760_, _38759_);
  or (_38769_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_38770_, \oc8051_gm_cxrom_1.cell1.data [6], _38654_);
  nand (_38771_, _38770_, _38769_);
  nand (_38775_, _38771_, _39026_);
  or (_38781_, \oc8051_gm_cxrom_1.cell1.data [6], _39026_);
  and (_00162_, _38781_, _38775_);
  or (_38782_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_38785_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_38791_, _38785_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_38793_, _38791_, _38782_);
  nand (_38794_, _38793_, _39026_);
  or (_38796_, \oc8051_gm_cxrom_1.cell2.data [7], _39026_);
  and (_00170_, _38796_, _38794_);
  or (_38804_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38805_, \oc8051_gm_cxrom_1.cell2.data [0], _38785_);
  nand (_38807_, _38805_, _38804_);
  nand (_38813_, _38807_, _39026_);
  or (_38816_, \oc8051_gm_cxrom_1.cell2.data [0], _39026_);
  and (_00203_, _38816_, _38813_);
  or (_38818_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38824_, \oc8051_gm_cxrom_1.cell2.data [1], _38785_);
  nand (_38826_, _38824_, _38818_);
  nand (_38827_, _38826_, _39026_);
  or (_38828_, \oc8051_gm_cxrom_1.cell2.data [1], _39026_);
  and (_00205_, _38828_, _38827_);
  or (_38829_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38830_, \oc8051_gm_cxrom_1.cell2.data [2], _38785_);
  nand (_38831_, _38830_, _38829_);
  nand (_38832_, _38831_, _39026_);
  or (_38833_, \oc8051_gm_cxrom_1.cell2.data [2], _39026_);
  and (_00207_, _38833_, _38832_);
  or (_38834_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38835_, \oc8051_gm_cxrom_1.cell2.data [3], _38785_);
  nand (_38836_, _38835_, _38834_);
  nand (_38837_, _38836_, _39026_);
  or (_38838_, \oc8051_gm_cxrom_1.cell2.data [3], _39026_);
  and (_00209_, _38838_, _38837_);
  or (_38839_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38840_, \oc8051_gm_cxrom_1.cell2.data [4], _38785_);
  nand (_38841_, _38840_, _38839_);
  nand (_38842_, _38841_, _39026_);
  or (_38843_, \oc8051_gm_cxrom_1.cell2.data [4], _39026_);
  and (_00211_, _38843_, _38842_);
  or (_38844_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38845_, \oc8051_gm_cxrom_1.cell2.data [5], _38785_);
  nand (_38846_, _38845_, _38844_);
  nand (_38847_, _38846_, _39026_);
  or (_38848_, \oc8051_gm_cxrom_1.cell2.data [5], _39026_);
  and (_00213_, _38848_, _38847_);
  or (_38849_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_38850_, \oc8051_gm_cxrom_1.cell2.data [6], _38785_);
  nand (_38851_, _38850_, _38849_);
  nand (_38852_, _38851_, _39026_);
  or (_38853_, \oc8051_gm_cxrom_1.cell2.data [6], _39026_);
  and (_00215_, _38853_, _38852_);
  or (_38854_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_38855_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_38856_, _38855_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_38857_, _38856_, _38854_);
  nand (_38858_, _38857_, _39026_);
  or (_38859_, \oc8051_gm_cxrom_1.cell3.data [7], _39026_);
  and (_00223_, _38859_, _38858_);
  or (_38860_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38861_, \oc8051_gm_cxrom_1.cell3.data [0], _38855_);
  nand (_38862_, _38861_, _38860_);
  nand (_38863_, _38862_, _39026_);
  or (_38864_, \oc8051_gm_cxrom_1.cell3.data [0], _39026_);
  and (_00255_, _38864_, _38863_);
  or (_38865_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38866_, \oc8051_gm_cxrom_1.cell3.data [1], _38855_);
  nand (_38867_, _38866_, _38865_);
  nand (_38868_, _38867_, _39026_);
  or (_38869_, \oc8051_gm_cxrom_1.cell3.data [1], _39026_);
  and (_00257_, _38869_, _38868_);
  or (_38870_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38871_, \oc8051_gm_cxrom_1.cell3.data [2], _38855_);
  nand (_38872_, _38871_, _38870_);
  nand (_38873_, _38872_, _39026_);
  or (_38874_, \oc8051_gm_cxrom_1.cell3.data [2], _39026_);
  and (_00258_, _38874_, _38873_);
  or (_38875_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38876_, \oc8051_gm_cxrom_1.cell3.data [3], _38855_);
  nand (_38877_, _38876_, _38875_);
  nand (_38878_, _38877_, _39026_);
  or (_38879_, \oc8051_gm_cxrom_1.cell3.data [3], _39026_);
  and (_00260_, _38879_, _38878_);
  or (_38880_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38881_, \oc8051_gm_cxrom_1.cell3.data [4], _38855_);
  nand (_38882_, _38881_, _38880_);
  nand (_38883_, _38882_, _39026_);
  or (_38884_, \oc8051_gm_cxrom_1.cell3.data [4], _39026_);
  and (_00262_, _38884_, _38883_);
  or (_38885_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38886_, \oc8051_gm_cxrom_1.cell3.data [5], _38855_);
  nand (_38887_, _38886_, _38885_);
  nand (_38888_, _38887_, _39026_);
  or (_38889_, \oc8051_gm_cxrom_1.cell3.data [5], _39026_);
  and (_00264_, _38889_, _38888_);
  or (_38890_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_38891_, \oc8051_gm_cxrom_1.cell3.data [6], _38855_);
  nand (_38892_, _38891_, _38890_);
  nand (_38893_, _38892_, _39026_);
  or (_38894_, \oc8051_gm_cxrom_1.cell3.data [6], _39026_);
  and (_00266_, _38894_, _38893_);
  or (_38895_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_38896_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_38897_, _38896_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_38898_, _38897_, _38895_);
  nand (_38899_, _38898_, _39026_);
  or (_38900_, \oc8051_gm_cxrom_1.cell4.data [7], _39026_);
  and (_00274_, _38900_, _38899_);
  or (_38901_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38902_, \oc8051_gm_cxrom_1.cell4.data [0], _38896_);
  nand (_38903_, _38902_, _38901_);
  nand (_38904_, _38903_, _39026_);
  or (_38905_, \oc8051_gm_cxrom_1.cell4.data [0], _39026_);
  and (_00306_, _38905_, _38904_);
  or (_38906_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38907_, \oc8051_gm_cxrom_1.cell4.data [1], _38896_);
  nand (_38908_, _38907_, _38906_);
  nand (_38909_, _38908_, _39026_);
  or (_38910_, \oc8051_gm_cxrom_1.cell4.data [1], _39026_);
  and (_00308_, _38910_, _38909_);
  or (_38911_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38912_, \oc8051_gm_cxrom_1.cell4.data [2], _38896_);
  nand (_38913_, _38912_, _38911_);
  nand (_38914_, _38913_, _39026_);
  or (_38915_, \oc8051_gm_cxrom_1.cell4.data [2], _39026_);
  and (_00310_, _38915_, _38914_);
  or (_38916_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38917_, \oc8051_gm_cxrom_1.cell4.data [3], _38896_);
  nand (_38918_, _38917_, _38916_);
  nand (_38919_, _38918_, _39026_);
  or (_38920_, \oc8051_gm_cxrom_1.cell4.data [3], _39026_);
  and (_00312_, _38920_, _38919_);
  or (_38921_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38922_, \oc8051_gm_cxrom_1.cell4.data [4], _38896_);
  nand (_38923_, _38922_, _38921_);
  nand (_38924_, _38923_, _39026_);
  or (_38925_, \oc8051_gm_cxrom_1.cell4.data [4], _39026_);
  and (_00314_, _38925_, _38924_);
  or (_38926_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38927_, \oc8051_gm_cxrom_1.cell4.data [5], _38896_);
  nand (_38928_, _38927_, _38926_);
  nand (_38929_, _38928_, _39026_);
  or (_38930_, \oc8051_gm_cxrom_1.cell4.data [5], _39026_);
  and (_00316_, _38930_, _38929_);
  or (_38931_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_38932_, \oc8051_gm_cxrom_1.cell4.data [6], _38896_);
  nand (_38933_, _38932_, _38931_);
  nand (_38934_, _38933_, _39026_);
  or (_38935_, \oc8051_gm_cxrom_1.cell4.data [6], _39026_);
  and (_00318_, _38935_, _38934_);
  or (_38936_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_38938_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_38939_, _38938_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_38940_, _38939_, _38936_);
  nand (_38941_, _38940_, _39026_);
  or (_38942_, \oc8051_gm_cxrom_1.cell5.data [7], _39026_);
  and (_00326_, _38942_, _38941_);
  or (_38943_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38944_, \oc8051_gm_cxrom_1.cell5.data [0], _38938_);
  nand (_38945_, _38944_, _38943_);
  nand (_38946_, _38945_, _39026_);
  or (_38947_, \oc8051_gm_cxrom_1.cell5.data [0], _39026_);
  and (_00358_, _38947_, _38946_);
  or (_38948_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38949_, \oc8051_gm_cxrom_1.cell5.data [1], _38938_);
  nand (_38950_, _38949_, _38948_);
  nand (_38951_, _38950_, _39026_);
  or (_38952_, \oc8051_gm_cxrom_1.cell5.data [1], _39026_);
  and (_00360_, _38952_, _38951_);
  or (_38953_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38954_, \oc8051_gm_cxrom_1.cell5.data [2], _38938_);
  nand (_38955_, _38954_, _38953_);
  nand (_38956_, _38955_, _39026_);
  or (_38957_, \oc8051_gm_cxrom_1.cell5.data [2], _39026_);
  and (_00362_, _38957_, _38956_);
  or (_38958_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38959_, \oc8051_gm_cxrom_1.cell5.data [3], _38938_);
  nand (_38960_, _38959_, _38958_);
  nand (_38961_, _38960_, _39026_);
  or (_38962_, \oc8051_gm_cxrom_1.cell5.data [3], _39026_);
  and (_00364_, _38962_, _38961_);
  or (_38963_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38964_, \oc8051_gm_cxrom_1.cell5.data [4], _38938_);
  nand (_38965_, _38964_, _38963_);
  nand (_38966_, _38965_, _39026_);
  or (_38967_, \oc8051_gm_cxrom_1.cell5.data [4], _39026_);
  and (_00366_, _38967_, _38966_);
  or (_38968_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38969_, \oc8051_gm_cxrom_1.cell5.data [5], _38938_);
  nand (_38970_, _38969_, _38968_);
  nand (_38971_, _38970_, _39026_);
  or (_38972_, \oc8051_gm_cxrom_1.cell5.data [5], _39026_);
  and (_00368_, _38972_, _38971_);
  or (_38974_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_38975_, \oc8051_gm_cxrom_1.cell5.data [6], _38938_);
  nand (_38976_, _38975_, _38974_);
  nand (_38977_, _38976_, _39026_);
  or (_38978_, \oc8051_gm_cxrom_1.cell5.data [6], _39026_);
  and (_00370_, _38978_, _38977_);
  or (_38979_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_38980_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_38981_, _38980_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_38982_, _38981_, _38979_);
  nand (_38983_, _38982_, _39026_);
  or (_38984_, \oc8051_gm_cxrom_1.cell6.data [7], _39026_);
  and (_00378_, _38984_, _38983_);
  or (_38985_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_38986_, \oc8051_gm_cxrom_1.cell6.data [0], _38980_);
  nand (_38987_, _38986_, _38985_);
  nand (_38988_, _38987_, _39026_);
  or (_38989_, \oc8051_gm_cxrom_1.cell6.data [0], _39026_);
  and (_00410_, _38989_, _38988_);
  or (_38990_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_38991_, \oc8051_gm_cxrom_1.cell6.data [1], _38980_);
  nand (_38992_, _38991_, _38990_);
  nand (_38994_, _38992_, _39026_);
  or (_38996_, \oc8051_gm_cxrom_1.cell6.data [1], _39026_);
  and (_00412_, _38996_, _38994_);
  or (_38998_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_38999_, \oc8051_gm_cxrom_1.cell6.data [2], _38980_);
  nand (_39000_, _38999_, _38998_);
  nand (_39001_, _39000_, _39026_);
  or (_39002_, \oc8051_gm_cxrom_1.cell6.data [2], _39026_);
  and (_00414_, _39002_, _39001_);
  or (_39003_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_39004_, \oc8051_gm_cxrom_1.cell6.data [3], _38980_);
  nand (_39005_, _39004_, _39003_);
  nand (_39006_, _39005_, _39026_);
  or (_39007_, \oc8051_gm_cxrom_1.cell6.data [3], _39026_);
  and (_00416_, _39007_, _39006_);
  or (_39008_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_39009_, \oc8051_gm_cxrom_1.cell6.data [4], _38980_);
  nand (_39010_, _39009_, _39008_);
  nand (_39011_, _39010_, _39026_);
  or (_39012_, \oc8051_gm_cxrom_1.cell6.data [4], _39026_);
  and (_00418_, _39012_, _39011_);
  or (_39013_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_39014_, \oc8051_gm_cxrom_1.cell6.data [5], _38980_);
  nand (_39015_, _39014_, _39013_);
  nand (_39016_, _39015_, _39026_);
  or (_39018_, \oc8051_gm_cxrom_1.cell6.data [5], _39026_);
  and (_00420_, _39018_, _39016_);
  or (_39021_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_39023_, \oc8051_gm_cxrom_1.cell6.data [6], _38980_);
  nand (_39025_, _39023_, _39021_);
  nand (_39027_, _39025_, _39026_);
  or (_39029_, \oc8051_gm_cxrom_1.cell6.data [6], _39026_);
  and (_00422_, _39029_, _39027_);
  or (_39032_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_39034_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_39035_, _39034_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_39036_, _39035_, _39032_);
  nand (_39037_, _39036_, _39026_);
  or (_39038_, \oc8051_gm_cxrom_1.cell7.data [7], _39026_);
  and (_00430_, _39038_, _39037_);
  or (_39039_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39040_, \oc8051_gm_cxrom_1.cell7.data [0], _39034_);
  nand (_39041_, _39040_, _39039_);
  nand (_39042_, _39041_, _39026_);
  or (_39043_, \oc8051_gm_cxrom_1.cell7.data [0], _39026_);
  and (_00462_, _39043_, _39042_);
  or (_39044_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39045_, \oc8051_gm_cxrom_1.cell7.data [1], _39034_);
  nand (_39046_, _39045_, _39044_);
  nand (_39047_, _39046_, _39026_);
  or (_39048_, \oc8051_gm_cxrom_1.cell7.data [1], _39026_);
  and (_00464_, _39048_, _39047_);
  or (_39049_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39050_, \oc8051_gm_cxrom_1.cell7.data [2], _39034_);
  nand (_39051_, _39050_, _39049_);
  nand (_39052_, _39051_, _39026_);
  or (_39053_, \oc8051_gm_cxrom_1.cell7.data [2], _39026_);
  and (_00466_, _39053_, _39052_);
  or (_39054_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39055_, \oc8051_gm_cxrom_1.cell7.data [3], _39034_);
  nand (_39056_, _39055_, _39054_);
  nand (_39057_, _39056_, _39026_);
  or (_39058_, \oc8051_gm_cxrom_1.cell7.data [3], _39026_);
  and (_00468_, _39058_, _39057_);
  or (_39059_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39060_, \oc8051_gm_cxrom_1.cell7.data [4], _39034_);
  nand (_39061_, _39060_, _39059_);
  nand (_39062_, _39061_, _39026_);
  or (_39063_, \oc8051_gm_cxrom_1.cell7.data [4], _39026_);
  and (_00470_, _39063_, _39062_);
  or (_39064_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39065_, \oc8051_gm_cxrom_1.cell7.data [5], _39034_);
  nand (_39066_, _39065_, _39064_);
  nand (_39067_, _39066_, _39026_);
  or (_39068_, \oc8051_gm_cxrom_1.cell7.data [5], _39026_);
  and (_00472_, _39068_, _39067_);
  or (_39069_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_39070_, \oc8051_gm_cxrom_1.cell7.data [6], _39034_);
  nand (_39071_, _39070_, _39069_);
  nand (_39072_, _39071_, _39026_);
  or (_39073_, \oc8051_gm_cxrom_1.cell7.data [6], _39026_);
  and (_00474_, _39073_, _39072_);
  or (_39074_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_39075_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_39076_, _39075_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_39077_, _39076_, _39074_);
  nand (_39078_, _39077_, _39026_);
  or (_39079_, \oc8051_gm_cxrom_1.cell8.data [7], _39026_);
  and (_00482_, _39079_, _39078_);
  or (_39080_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39081_, \oc8051_gm_cxrom_1.cell8.data [0], _39075_);
  nand (_39082_, _39081_, _39080_);
  nand (_39083_, _39082_, _39026_);
  or (_39084_, \oc8051_gm_cxrom_1.cell8.data [0], _39026_);
  and (_00514_, _39084_, _39083_);
  or (_39085_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39086_, \oc8051_gm_cxrom_1.cell8.data [1], _39075_);
  nand (_39087_, _39086_, _39085_);
  nand (_39088_, _39087_, _39026_);
  or (_39089_, \oc8051_gm_cxrom_1.cell8.data [1], _39026_);
  and (_00516_, _39089_, _39088_);
  or (_39090_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39091_, \oc8051_gm_cxrom_1.cell8.data [2], _39075_);
  nand (_39092_, _39091_, _39090_);
  nand (_39093_, _39092_, _39026_);
  or (_39094_, \oc8051_gm_cxrom_1.cell8.data [2], _39026_);
  and (_00518_, _39094_, _39093_);
  or (_39095_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39096_, \oc8051_gm_cxrom_1.cell8.data [3], _39075_);
  nand (_39097_, _39096_, _39095_);
  nand (_39098_, _39097_, _39026_);
  or (_39099_, \oc8051_gm_cxrom_1.cell8.data [3], _39026_);
  and (_00520_, _39099_, _39098_);
  or (_39100_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39101_, \oc8051_gm_cxrom_1.cell8.data [4], _39075_);
  nand (_39102_, _39101_, _39100_);
  nand (_39103_, _39102_, _39026_);
  or (_39104_, \oc8051_gm_cxrom_1.cell8.data [4], _39026_);
  and (_00522_, _39104_, _39103_);
  or (_39105_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39106_, \oc8051_gm_cxrom_1.cell8.data [5], _39075_);
  nand (_39107_, _39106_, _39105_);
  nand (_39108_, _39107_, _39026_);
  or (_39109_, \oc8051_gm_cxrom_1.cell8.data [5], _39026_);
  and (_00524_, _39109_, _39108_);
  or (_39110_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_39111_, \oc8051_gm_cxrom_1.cell8.data [6], _39075_);
  nand (_39112_, _39111_, _39110_);
  nand (_39113_, _39112_, _39026_);
  or (_39114_, \oc8051_gm_cxrom_1.cell8.data [6], _39026_);
  and (_00526_, _39114_, _39113_);
  or (_39115_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_39116_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_39117_, _39116_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_39118_, _39117_, _39115_);
  nand (_39119_, _39118_, _39026_);
  or (_39120_, \oc8051_gm_cxrom_1.cell9.data [7], _39026_);
  and (_00534_, _39120_, _39119_);
  or (_39121_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39122_, \oc8051_gm_cxrom_1.cell9.data [0], _39116_);
  nand (_39123_, _39122_, _39121_);
  nand (_39124_, _39123_, _39026_);
  or (_39125_, \oc8051_gm_cxrom_1.cell9.data [0], _39026_);
  and (_00566_, _39125_, _39124_);
  or (_39126_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39127_, \oc8051_gm_cxrom_1.cell9.data [1], _39116_);
  nand (_39128_, _39127_, _39126_);
  nand (_39129_, _39128_, _39026_);
  or (_39130_, \oc8051_gm_cxrom_1.cell9.data [1], _39026_);
  and (_00568_, _39130_, _39129_);
  or (_39131_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39132_, \oc8051_gm_cxrom_1.cell9.data [2], _39116_);
  nand (_39133_, _39132_, _39131_);
  nand (_39134_, _39133_, _39026_);
  or (_39135_, \oc8051_gm_cxrom_1.cell9.data [2], _39026_);
  and (_00570_, _39135_, _39134_);
  or (_39136_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39137_, \oc8051_gm_cxrom_1.cell9.data [3], _39116_);
  nand (_39138_, _39137_, _39136_);
  nand (_39139_, _39138_, _39026_);
  or (_39140_, \oc8051_gm_cxrom_1.cell9.data [3], _39026_);
  and (_00572_, _39140_, _39139_);
  or (_39141_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39142_, \oc8051_gm_cxrom_1.cell9.data [4], _39116_);
  nand (_39143_, _39142_, _39141_);
  nand (_39144_, _39143_, _39026_);
  or (_39145_, \oc8051_gm_cxrom_1.cell9.data [4], _39026_);
  and (_00574_, _39145_, _39144_);
  or (_39146_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39147_, \oc8051_gm_cxrom_1.cell9.data [5], _39116_);
  nand (_39148_, _39147_, _39146_);
  nand (_39149_, _39148_, _39026_);
  or (_39150_, \oc8051_gm_cxrom_1.cell9.data [5], _39026_);
  and (_00576_, _39150_, _39149_);
  or (_39151_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_39152_, \oc8051_gm_cxrom_1.cell9.data [6], _39116_);
  nand (_39153_, _39152_, _39151_);
  nand (_39154_, _39153_, _39026_);
  or (_39155_, \oc8051_gm_cxrom_1.cell9.data [6], _39026_);
  and (_00578_, _39155_, _39154_);
  or (_39156_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_39157_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_39158_, _39157_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_39159_, _39158_, _39156_);
  nand (_39160_, _39159_, _39026_);
  or (_39161_, \oc8051_gm_cxrom_1.cell10.data [7], _39026_);
  and (_00586_, _39161_, _39160_);
  or (_39162_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39163_, \oc8051_gm_cxrom_1.cell10.data [0], _39157_);
  nand (_39164_, _39163_, _39162_);
  nand (_39165_, _39164_, _39026_);
  or (_39166_, \oc8051_gm_cxrom_1.cell10.data [0], _39026_);
  and (_00618_, _39166_, _39165_);
  or (_39167_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39168_, \oc8051_gm_cxrom_1.cell10.data [1], _39157_);
  nand (_39169_, _39168_, _39167_);
  nand (_39170_, _39169_, _39026_);
  or (_39171_, \oc8051_gm_cxrom_1.cell10.data [1], _39026_);
  and (_00620_, _39171_, _39170_);
  or (_39172_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39173_, \oc8051_gm_cxrom_1.cell10.data [2], _39157_);
  nand (_39174_, _39173_, _39172_);
  nand (_39175_, _39174_, _39026_);
  or (_39176_, \oc8051_gm_cxrom_1.cell10.data [2], _39026_);
  and (_00622_, _39176_, _39175_);
  or (_39177_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39178_, \oc8051_gm_cxrom_1.cell10.data [3], _39157_);
  nand (_39179_, _39178_, _39177_);
  nand (_39180_, _39179_, _39026_);
  or (_39181_, \oc8051_gm_cxrom_1.cell10.data [3], _39026_);
  and (_00624_, _39181_, _39180_);
  or (_39182_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39183_, \oc8051_gm_cxrom_1.cell10.data [4], _39157_);
  nand (_39184_, _39183_, _39182_);
  nand (_39185_, _39184_, _39026_);
  or (_39186_, \oc8051_gm_cxrom_1.cell10.data [4], _39026_);
  and (_00626_, _39186_, _39185_);
  or (_39187_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39188_, \oc8051_gm_cxrom_1.cell10.data [5], _39157_);
  nand (_39189_, _39188_, _39187_);
  nand (_39190_, _39189_, _39026_);
  or (_39191_, \oc8051_gm_cxrom_1.cell10.data [5], _39026_);
  and (_00628_, _39191_, _39190_);
  or (_39192_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_39193_, \oc8051_gm_cxrom_1.cell10.data [6], _39157_);
  nand (_39194_, _39193_, _39192_);
  nand (_39195_, _39194_, _39026_);
  or (_39196_, \oc8051_gm_cxrom_1.cell10.data [6], _39026_);
  and (_00630_, _39196_, _39195_);
  or (_39197_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_39198_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_39199_, _39198_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_39200_, _39199_, _39197_);
  nand (_39201_, _39200_, _39026_);
  or (_39202_, \oc8051_gm_cxrom_1.cell11.data [7], _39026_);
  and (_00638_, _39202_, _39201_);
  or (_39203_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39204_, \oc8051_gm_cxrom_1.cell11.data [0], _39198_);
  nand (_39205_, _39204_, _39203_);
  nand (_39206_, _39205_, _39026_);
  or (_39207_, \oc8051_gm_cxrom_1.cell11.data [0], _39026_);
  and (_00670_, _39207_, _39206_);
  or (_39208_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39209_, \oc8051_gm_cxrom_1.cell11.data [1], _39198_);
  nand (_39210_, _39209_, _39208_);
  nand (_39211_, _39210_, _39026_);
  or (_39212_, \oc8051_gm_cxrom_1.cell11.data [1], _39026_);
  and (_00672_, _39212_, _39211_);
  or (_39213_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39214_, \oc8051_gm_cxrom_1.cell11.data [2], _39198_);
  nand (_39215_, _39214_, _39213_);
  nand (_39216_, _39215_, _39026_);
  or (_39217_, \oc8051_gm_cxrom_1.cell11.data [2], _39026_);
  and (_00674_, _39217_, _39216_);
  or (_39218_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39219_, \oc8051_gm_cxrom_1.cell11.data [3], _39198_);
  nand (_39220_, _39219_, _39218_);
  nand (_39221_, _39220_, _39026_);
  or (_39222_, \oc8051_gm_cxrom_1.cell11.data [3], _39026_);
  and (_00676_, _39222_, _39221_);
  or (_39223_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39224_, \oc8051_gm_cxrom_1.cell11.data [4], _39198_);
  nand (_39225_, _39224_, _39223_);
  nand (_39226_, _39225_, _39026_);
  or (_39227_, \oc8051_gm_cxrom_1.cell11.data [4], _39026_);
  and (_00678_, _39227_, _39226_);
  or (_39228_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39229_, \oc8051_gm_cxrom_1.cell11.data [5], _39198_);
  nand (_39230_, _39229_, _39228_);
  nand (_39231_, _39230_, _39026_);
  or (_39232_, \oc8051_gm_cxrom_1.cell11.data [5], _39026_);
  and (_00680_, _39232_, _39231_);
  or (_39233_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_39234_, \oc8051_gm_cxrom_1.cell11.data [6], _39198_);
  nand (_39235_, _39234_, _39233_);
  nand (_39236_, _39235_, _39026_);
  or (_39237_, \oc8051_gm_cxrom_1.cell11.data [6], _39026_);
  and (_00682_, _39237_, _39236_);
  or (_39238_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_39239_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_39240_, _39239_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_39241_, _39240_, _39238_);
  nand (_39242_, _39241_, _39026_);
  or (_39243_, \oc8051_gm_cxrom_1.cell12.data [7], _39026_);
  and (_00690_, _39243_, _39242_);
  or (_39244_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39245_, \oc8051_gm_cxrom_1.cell12.data [0], _39239_);
  nand (_39246_, _39245_, _39244_);
  nand (_39247_, _39246_, _39026_);
  or (_39248_, \oc8051_gm_cxrom_1.cell12.data [0], _39026_);
  and (_00722_, _39248_, _39247_);
  or (_39249_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39250_, \oc8051_gm_cxrom_1.cell12.data [1], _39239_);
  nand (_39251_, _39250_, _39249_);
  nand (_39252_, _39251_, _39026_);
  or (_39253_, \oc8051_gm_cxrom_1.cell12.data [1], _39026_);
  and (_00724_, _39253_, _39252_);
  or (_39254_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39255_, \oc8051_gm_cxrom_1.cell12.data [2], _39239_);
  nand (_39256_, _39255_, _39254_);
  nand (_39257_, _39256_, _39026_);
  or (_39258_, \oc8051_gm_cxrom_1.cell12.data [2], _39026_);
  and (_00726_, _39258_, _39257_);
  or (_39259_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39260_, \oc8051_gm_cxrom_1.cell12.data [3], _39239_);
  nand (_39261_, _39260_, _39259_);
  nand (_39262_, _39261_, _39026_);
  or (_39263_, \oc8051_gm_cxrom_1.cell12.data [3], _39026_);
  and (_00728_, _39263_, _39262_);
  or (_39264_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39265_, \oc8051_gm_cxrom_1.cell12.data [4], _39239_);
  nand (_39266_, _39265_, _39264_);
  nand (_39267_, _39266_, _39026_);
  or (_39268_, \oc8051_gm_cxrom_1.cell12.data [4], _39026_);
  and (_00730_, _39268_, _39267_);
  or (_39269_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39270_, \oc8051_gm_cxrom_1.cell12.data [5], _39239_);
  nand (_39271_, _39270_, _39269_);
  nand (_39272_, _39271_, _39026_);
  or (_39273_, \oc8051_gm_cxrom_1.cell12.data [5], _39026_);
  and (_00732_, _39273_, _39272_);
  or (_39274_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_39275_, \oc8051_gm_cxrom_1.cell12.data [6], _39239_);
  nand (_39276_, _39275_, _39274_);
  nand (_39277_, _39276_, _39026_);
  or (_39278_, \oc8051_gm_cxrom_1.cell12.data [6], _39026_);
  and (_00734_, _39278_, _39277_);
  or (_39279_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_39280_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_39281_, _39280_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_39282_, _39281_, _39279_);
  nand (_39283_, _39282_, _39026_);
  or (_39284_, \oc8051_gm_cxrom_1.cell13.data [7], _39026_);
  and (_00742_, _39284_, _39283_);
  or (_39285_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39286_, \oc8051_gm_cxrom_1.cell13.data [0], _39280_);
  nand (_39287_, _39286_, _39285_);
  nand (_39288_, _39287_, _39026_);
  or (_39289_, \oc8051_gm_cxrom_1.cell13.data [0], _39026_);
  and (_00774_, _39289_, _39288_);
  or (_39290_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39291_, \oc8051_gm_cxrom_1.cell13.data [1], _39280_);
  nand (_39292_, _39291_, _39290_);
  nand (_39293_, _39292_, _39026_);
  or (_39294_, \oc8051_gm_cxrom_1.cell13.data [1], _39026_);
  and (_00776_, _39294_, _39293_);
  or (_39295_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39296_, \oc8051_gm_cxrom_1.cell13.data [2], _39280_);
  nand (_39297_, _39296_, _39295_);
  nand (_39298_, _39297_, _39026_);
  or (_39299_, \oc8051_gm_cxrom_1.cell13.data [2], _39026_);
  and (_00778_, _39299_, _39298_);
  or (_39300_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39301_, \oc8051_gm_cxrom_1.cell13.data [3], _39280_);
  nand (_39302_, _39301_, _39300_);
  nand (_39303_, _39302_, _39026_);
  or (_39304_, \oc8051_gm_cxrom_1.cell13.data [3], _39026_);
  and (_00780_, _39304_, _39303_);
  or (_39305_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39306_, \oc8051_gm_cxrom_1.cell13.data [4], _39280_);
  nand (_39307_, _39306_, _39305_);
  nand (_39308_, _39307_, _39026_);
  or (_39309_, \oc8051_gm_cxrom_1.cell13.data [4], _39026_);
  and (_00782_, _39309_, _39308_);
  or (_39310_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39311_, \oc8051_gm_cxrom_1.cell13.data [5], _39280_);
  nand (_39312_, _39311_, _39310_);
  nand (_39313_, _39312_, _39026_);
  or (_39314_, \oc8051_gm_cxrom_1.cell13.data [5], _39026_);
  and (_00784_, _39314_, _39313_);
  or (_39315_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_39316_, \oc8051_gm_cxrom_1.cell13.data [6], _39280_);
  nand (_39317_, _39316_, _39315_);
  nand (_39318_, _39317_, _39026_);
  or (_39319_, \oc8051_gm_cxrom_1.cell13.data [6], _39026_);
  and (_00786_, _39319_, _39318_);
  or (_39320_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_39321_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_39322_, _39321_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_39323_, _39322_, _39320_);
  nand (_39324_, _39323_, _39026_);
  or (_39325_, \oc8051_gm_cxrom_1.cell14.data [7], _39026_);
  and (_00794_, _39325_, _39324_);
  or (_39326_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39327_, \oc8051_gm_cxrom_1.cell14.data [0], _39321_);
  nand (_39328_, _39327_, _39326_);
  nand (_39329_, _39328_, _39026_);
  or (_39330_, \oc8051_gm_cxrom_1.cell14.data [0], _39026_);
  and (_00826_, _39330_, _39329_);
  or (_39331_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39332_, \oc8051_gm_cxrom_1.cell14.data [1], _39321_);
  nand (_39333_, _39332_, _39331_);
  nand (_39334_, _39333_, _39026_);
  or (_39335_, \oc8051_gm_cxrom_1.cell14.data [1], _39026_);
  and (_00828_, _39335_, _39334_);
  or (_39336_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39337_, \oc8051_gm_cxrom_1.cell14.data [2], _39321_);
  nand (_39338_, _39337_, _39336_);
  nand (_39339_, _39338_, _39026_);
  or (_39340_, \oc8051_gm_cxrom_1.cell14.data [2], _39026_);
  and (_00829_, _39340_, _39339_);
  or (_39341_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39342_, \oc8051_gm_cxrom_1.cell14.data [3], _39321_);
  nand (_39343_, _39342_, _39341_);
  nand (_39344_, _39343_, _39026_);
  or (_39345_, \oc8051_gm_cxrom_1.cell14.data [3], _39026_);
  and (_00831_, _39345_, _39344_);
  or (_39346_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39347_, \oc8051_gm_cxrom_1.cell14.data [4], _39321_);
  nand (_39348_, _39347_, _39346_);
  nand (_39349_, _39348_, _39026_);
  or (_39350_, \oc8051_gm_cxrom_1.cell14.data [4], _39026_);
  and (_00833_, _39350_, _39349_);
  or (_39351_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39352_, \oc8051_gm_cxrom_1.cell14.data [5], _39321_);
  nand (_39353_, _39352_, _39351_);
  nand (_39354_, _39353_, _39026_);
  or (_39355_, \oc8051_gm_cxrom_1.cell14.data [5], _39026_);
  and (_00835_, _39355_, _39354_);
  or (_39356_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_39357_, \oc8051_gm_cxrom_1.cell14.data [6], _39321_);
  nand (_39358_, _39357_, _39356_);
  nand (_39359_, _39358_, _39026_);
  or (_39360_, \oc8051_gm_cxrom_1.cell14.data [6], _39026_);
  and (_00837_, _39360_, _39359_);
  or (_39361_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_39362_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_39363_, _39362_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_39364_, _39363_, _39361_);
  nand (_39365_, _39364_, _39026_);
  or (_39366_, \oc8051_gm_cxrom_1.cell15.data [7], _39026_);
  and (_00845_, _39366_, _39365_);
  or (_39367_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39368_, \oc8051_gm_cxrom_1.cell15.data [0], _39362_);
  nand (_39369_, _39368_, _39367_);
  nand (_39370_, _39369_, _39026_);
  or (_39371_, \oc8051_gm_cxrom_1.cell15.data [0], _39026_);
  and (_00877_, _39371_, _39370_);
  or (_39372_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39373_, \oc8051_gm_cxrom_1.cell15.data [1], _39362_);
  nand (_39374_, _39373_, _39372_);
  nand (_39375_, _39374_, _39026_);
  or (_39376_, \oc8051_gm_cxrom_1.cell15.data [1], _39026_);
  and (_00879_, _39376_, _39375_);
  or (_39377_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39378_, \oc8051_gm_cxrom_1.cell15.data [2], _39362_);
  nand (_39379_, _39378_, _39377_);
  nand (_39380_, _39379_, _39026_);
  or (_39381_, \oc8051_gm_cxrom_1.cell15.data [2], _39026_);
  and (_00881_, _39381_, _39380_);
  or (_39382_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39383_, \oc8051_gm_cxrom_1.cell15.data [3], _39362_);
  nand (_39384_, _39383_, _39382_);
  nand (_39385_, _39384_, _39026_);
  or (_39386_, \oc8051_gm_cxrom_1.cell15.data [3], _39026_);
  and (_00883_, _39386_, _39385_);
  or (_39387_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39388_, \oc8051_gm_cxrom_1.cell15.data [4], _39362_);
  nand (_39389_, _39388_, _39387_);
  nand (_39390_, _39389_, _39026_);
  or (_39391_, \oc8051_gm_cxrom_1.cell15.data [4], _39026_);
  and (_00885_, _39391_, _39390_);
  or (_39392_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39393_, \oc8051_gm_cxrom_1.cell15.data [5], _39362_);
  nand (_39394_, _39393_, _39392_);
  nand (_39395_, _39394_, _39026_);
  or (_39396_, \oc8051_gm_cxrom_1.cell15.data [5], _39026_);
  and (_00887_, _39396_, _39395_);
  or (_39397_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_39398_, \oc8051_gm_cxrom_1.cell15.data [6], _39362_);
  nand (_39399_, _39398_, _39397_);
  nand (_39400_, _39399_, _39026_);
  or (_39401_, \oc8051_gm_cxrom_1.cell15.data [6], _39026_);
  and (_00889_, _39401_, _39400_);
  nor (_00920_, _20304_, rst);
  nor (_00924_, _37299_, rst);
  and (_39402_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_39403_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_39404_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_39405_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_39406_, _39405_, _39404_);
  and (_39407_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_39408_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_39409_, _39408_, _39407_);
  and (_39410_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_39411_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_39412_, _39411_, _39410_);
  and (_39413_, _39412_, _39409_);
  and (_39414_, _39413_, _39406_);
  nor (_39415_, _39414_, _18729_);
  nor (_39416_, _39415_, _39403_);
  nor (_39417_, _39416_, _37283_);
  nor (_39418_, _39417_, _39402_);
  nor (_00928_, _39418_, rst);
  nor (_01049_, _21089_, rst);
  and (_01052_, _19584_, _39026_);
  nor (_01055_, _19286_, rst);
  nor (_01058_, _19046_, rst);
  and (_01060_, _20598_, _39026_);
  nor (_01063_, _19835_, rst);
  nor (_01066_, _20075_, rst);
  nor (_01069_, _37585_, rst);
  nor (_01072_, _37494_, rst);
  nor (_01075_, _37427_, rst);
  nor (_01078_, _37547_, rst);
  nor (_01081_, _37455_, rst);
  nor (_01084_, _37383_, rst);
  nor (_01087_, _37611_, rst);
  and (_39419_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_39420_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_39421_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_39422_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_39423_, _39422_, _39421_);
  and (_39424_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_39425_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_39426_, _39425_, _39424_);
  and (_39427_, _39426_, _39423_);
  and (_39428_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_39429_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_39430_, _39429_, _39428_);
  and (_39431_, _39430_, _39427_);
  nor (_39432_, _39431_, _18729_);
  nor (_39433_, _39432_, _39420_);
  nor (_39434_, _39433_, _37283_);
  nor (_39435_, _39434_, _39419_);
  nor (_01090_, _39435_, rst);
  and (_39436_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_39437_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_39438_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_39439_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_39440_, _39439_, _39438_);
  and (_39441_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_39442_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_39443_, _39442_, _39441_);
  and (_39444_, _39443_, _39440_);
  and (_39445_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_39446_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_39447_, _39446_, _39445_);
  and (_39448_, _39447_, _39444_);
  nor (_39449_, _39448_, _18729_);
  nor (_39450_, _39449_, _39437_);
  nor (_39451_, _39450_, _37283_);
  nor (_39452_, _39451_, _39436_);
  nor (_01093_, _39452_, rst);
  and (_39453_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_39454_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_39455_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_39456_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_39457_, _39456_, _39455_);
  and (_39458_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_39459_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_39460_, _39459_, _39458_);
  and (_39461_, _39460_, _39457_);
  and (_39462_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_39463_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_39464_, _39463_, _39462_);
  and (_39465_, _39464_, _39461_);
  nor (_39466_, _39465_, _18729_);
  nor (_39467_, _39466_, _39454_);
  nor (_39468_, _39467_, _37283_);
  nor (_39469_, _39468_, _39453_);
  nor (_01096_, _39469_, rst);
  and (_39470_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_39471_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_39472_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_39473_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_39474_, _39473_, _39472_);
  and (_39475_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_39476_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_39477_, _39476_, _39475_);
  and (_39478_, _39477_, _39474_);
  and (_39479_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_39480_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_39481_, _39480_, _39479_);
  and (_39482_, _39481_, _39478_);
  nor (_39483_, _39482_, _18729_);
  nor (_39484_, _39483_, _39471_);
  nor (_39485_, _39484_, _37283_);
  nor (_39486_, _39485_, _39470_);
  nor (_01099_, _39486_, rst);
  and (_39487_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_39488_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_39489_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_39490_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_39491_, _39490_, _39489_);
  and (_39492_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_39493_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_39494_, _39493_, _39492_);
  and (_39495_, _39494_, _39491_);
  and (_39496_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_39497_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_39498_, _39497_, _39496_);
  and (_39499_, _39498_, _39495_);
  nor (_39500_, _39499_, _18729_);
  nor (_39501_, _39500_, _39488_);
  nor (_39502_, _39501_, _37283_);
  nor (_39503_, _39502_, _39487_);
  nor (_01102_, _39503_, rst);
  and (_39504_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_39505_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_39506_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_39507_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_39508_, _39507_, _39506_);
  and (_39509_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_39510_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_39511_, _39510_, _39509_);
  and (_39512_, _39511_, _39508_);
  and (_39513_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_39514_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_39515_, _39514_, _39513_);
  and (_39516_, _39515_, _39512_);
  nor (_39517_, _39516_, _18729_);
  nor (_39518_, _39517_, _39505_);
  nor (_39519_, _39518_, _37283_);
  nor (_39520_, _39519_, _39504_);
  nor (_01105_, _39520_, rst);
  and (_39521_, _37283_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_39522_, _18729_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_39523_, _18795_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_39524_, _18893_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_39525_, _39524_, _39523_);
  and (_39526_, _18947_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_39527_, _18849_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_39528_, _39527_, _39526_);
  and (_39529_, _39528_, _39525_);
  and (_39530_, _18926_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_39531_, _18762_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_39532_, _39531_, _39530_);
  and (_39533_, _39532_, _39529_);
  nor (_39534_, _39533_, _18729_);
  nor (_39535_, _39534_, _39522_);
  nor (_39536_, _39535_, _37283_);
  nor (_39537_, _39536_, _39521_);
  nor (_01107_, _39537_, rst);
  not (_39538_, _37631_);
  nor (_39539_, _39538_, _37342_);
  nor (_39540_, _37476_, _37394_);
  and (_39541_, _39540_, _39539_);
  and (_39542_, _39541_, _37552_);
  nor (_39543_, _37475_, _37394_);
  and (_39544_, _39543_, _39539_);
  and (_39545_, _39544_, _37552_);
  nor (_39546_, _39545_, _39542_);
  and (_39547_, _37476_, _37394_);
  and (_39548_, _39547_, _39539_);
  and (_39549_, _39548_, _37552_);
  nor (_39550_, _37476_, _37342_);
  and (_39551_, _37631_, _37394_);
  and (_39552_, _39551_, _39550_);
  and (_39553_, _39552_, _37552_);
  nor (_39554_, _39553_, _39549_);
  and (_39555_, _39554_, _39546_);
  and (_39556_, _39550_, _37553_);
  and (_39557_, _39556_, _37631_);
  and (_39558_, _37552_, _37476_);
  nor (_39559_, _37631_, _37342_);
  and (_39560_, _39559_, _39558_);
  nor (_39561_, _39560_, _39557_);
  and (_39562_, _39548_, _37553_);
  not (_39563_, _39562_);
  and (_39564_, _39559_, _39540_);
  and (_39565_, _39564_, _37552_);
  and (_39566_, _39544_, _37553_);
  nor (_39567_, _39566_, _39565_);
  and (_39568_, _39567_, _39563_);
  and (_39569_, _39568_, _39561_);
  and (_39570_, _39569_, _39555_);
  not (_39571_, _39570_);
  nor (_39572_, _37342_, _16372_);
  and (_39573_, _37342_, _16372_);
  nor (_39574_, _39573_, _39572_);
  nor (_39575_, _37394_, _16057_);
  and (_39576_, _37394_, _16057_);
  nor (_39577_, _39576_, _39575_);
  nor (_39578_, _37631_, _16198_);
  and (_39579_, _37631_, _16198_);
  nor (_39580_, _39579_, _39578_);
  nor (_39581_, _39580_, _39577_);
  nor (_39582_, _37552_, _16547_);
  and (_39583_, _37552_, _16547_);
  nor (_39584_, _39583_, _39582_);
  nor (_39585_, _37475_, _16721_);
  and (_39586_, _37475_, _16721_);
  nor (_39587_, _39586_, _39585_);
  nor (_39588_, _39587_, _39584_);
  nand (_39589_, _39588_, _39581_);
  nor (_39590_, _39589_, _39574_);
  nor (_39591_, _37514_, _17123_);
  and (_39592_, _37514_, _17123_);
  nor (_39593_, _39592_, _39591_);
  not (_39594_, _39593_);
  nor (_39595_, _37590_, _17004_);
  and (_39596_, _37590_, _17004_);
  nor (_39597_, _39596_, _39595_);
  nor (_39598_, _37432_, _16873_);
  and (_39599_, _37432_, _16873_);
  nor (_39600_, _39599_, _39598_);
  nor (_39601_, _39600_, _39597_);
  and (_39602_, _39601_, _39594_);
  and (_39603_, _39602_, _39590_);
  and (_39604_, _39603_, _15752_);
  and (_39605_, _39604_, _39571_);
  not (_39606_, _37514_);
  nor (_39607_, _37590_, _39606_);
  and (_39608_, _22621_, _21372_);
  not (_39609_, _39608_);
  nor (_39610_, _21972_, _22335_);
  and (_39611_, _39610_, _39609_);
  and (_39612_, _20620_, _19067_);
  and (_39613_, _39612_, _20816_);
  or (_39614_, _39613_, _20827_);
  and (_39615_, _22368_, _22621_);
  or (_39616_, _39615_, _22478_);
  nor (_39617_, _39616_, _39614_);
  and (_39618_, _39617_, _39611_);
  and (_39619_, _21776_, _21874_);
  nor (_39620_, _39619_, _21906_);
  not (_39621_, _20358_);
  and (_39622_, _22313_, _39621_);
  nor (_39623_, _21143_, _20347_);
  not (_39624_, _39623_);
  and (_39625_, _39624_, _19067_);
  not (_39626_, _39625_);
  and (_39627_, _39626_, _39622_);
  and (_39628_, _39627_, _39620_);
  and (_39629_, _39628_, _39618_);
  and (_39630_, _39629_, _22247_);
  nor (_39631_, _39630_, _18609_);
  and (_39632_, _18664_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_39633_, _39632_);
  and (_39634_, _39633_, p1in_reg[1]);
  and (_39635_, _39632_, p1_in[1]);
  or (_39636_, _39635_, _39634_);
  or (_39637_, _39636_, _39631_);
  not (_39638_, _39631_);
  or (_39639_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_39640_, _39639_, _39637_);
  and (_39641_, _39640_, _39607_);
  and (_39642_, _37590_, _37514_);
  and (_39643_, _39633_, p1in_reg[0]);
  and (_39644_, _39632_, p1_in[0]);
  or (_39645_, _39644_, _39643_);
  or (_39646_, _39645_, _39631_);
  nand (_39647_, _39631_, _29181_);
  and (_39648_, _39647_, _39646_);
  and (_39649_, _39648_, _39642_);
  or (_39650_, _39649_, _39641_);
  and (_39651_, _37590_, _39606_);
  and (_39652_, _39633_, p1in_reg[2]);
  and (_39653_, _39632_, p1_in[2]);
  or (_39654_, _39653_, _39652_);
  or (_39655_, _39654_, _39631_);
  nand (_39656_, _39631_, _29464_);
  and (_39657_, _39656_, _39655_);
  and (_39658_, _39657_, _39651_);
  nor (_39659_, _37590_, _37514_);
  and (_39660_, _39633_, p1in_reg[3]);
  and (_39661_, _39632_, p1_in[3]);
  or (_39662_, _39661_, _39660_);
  or (_39663_, _39662_, _39631_);
  or (_39664_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_39665_, _39664_, _39663_);
  and (_39666_, _39665_, _39659_);
  or (_39667_, _39666_, _39658_);
  or (_39668_, _39667_, _39650_);
  and (_39669_, _39668_, _37432_);
  not (_39670_, _37432_);
  and (_39671_, _39633_, p1in_reg[5]);
  and (_39672_, _39632_, p1_in[5]);
  or (_39673_, _39672_, _39671_);
  or (_39674_, _39673_, _39631_);
  nand (_39675_, _39631_, _29910_);
  and (_39676_, _39675_, _39674_);
  and (_39677_, _39676_, _39607_);
  and (_39678_, _39633_, p1in_reg[4]);
  and (_39679_, _39632_, p1_in[4]);
  or (_39680_, _39679_, _39678_);
  or (_39681_, _39680_, _39631_);
  nand (_39682_, _39631_, _29758_);
  and (_39683_, _39682_, _39681_);
  and (_39684_, _39683_, _39642_);
  or (_39685_, _39684_, _39677_);
  and (_39686_, _39633_, p1in_reg[6]);
  and (_39687_, _39632_, p1_in[6]);
  or (_39688_, _39687_, _39686_);
  or (_39689_, _39688_, _39631_);
  nand (_39690_, _39631_, _30061_);
  and (_39691_, _39690_, _39689_);
  and (_39692_, _39691_, _39651_);
  and (_39693_, _39633_, p1in_reg[7]);
  and (_39694_, _39632_, p1_in[7]);
  or (_39695_, _39694_, _39693_);
  or (_39696_, _39695_, _39631_);
  nand (_39697_, _39631_, _27644_);
  and (_39698_, _39697_, _39696_);
  and (_39699_, _39698_, _39659_);
  or (_39700_, _39699_, _39692_);
  or (_39701_, _39700_, _39685_);
  and (_39702_, _39701_, _39670_);
  or (_39703_, _39702_, _39669_);
  and (_39704_, _39703_, _39548_);
  and (_39705_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_39706_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_39707_, _39706_, _39705_);
  and (_39708_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_39709_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_39710_, _39709_, _39708_);
  or (_39711_, _39710_, _39707_);
  and (_39712_, _39711_, _37432_);
  and (_39713_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_39714_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_39715_, _39714_, _39713_);
  and (_39716_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_39717_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_39718_, _39717_, _39716_);
  or (_39719_, _39718_, _39715_);
  and (_39720_, _39719_, _39670_);
  or (_39721_, _39720_, _39712_);
  and (_39722_, _39559_, _39543_);
  and (_39723_, _39722_, _39721_);
  or (_39724_, _39723_, _39704_);
  and (_39725_, _39724_, _37552_);
  and (_39726_, _39633_, p3in_reg[0]);
  and (_39727_, _39632_, p3_in[0]);
  or (_39728_, _39727_, _39726_);
  or (_39729_, _39728_, _39631_);
  nand (_39730_, _39631_, _31307_);
  and (_39731_, _39730_, _39729_);
  or (_39732_, _39731_, _39670_);
  and (_39733_, _39633_, p3in_reg[4]);
  and (_39734_, _39632_, p3_in[4]);
  or (_39735_, _39734_, _39733_);
  or (_39736_, _39735_, _39631_);
  nand (_39737_, _39631_, _31961_);
  and (_39738_, _39737_, _39736_);
  or (_39739_, _39738_, _37432_);
  and (_39740_, _39739_, _39642_);
  and (_39741_, _39740_, _39732_);
  and (_39742_, _39633_, p3in_reg[3]);
  and (_39743_, _39632_, p3_in[3]);
  or (_39744_, _39743_, _39742_);
  or (_39745_, _39744_, _39631_);
  nand (_39746_, _39631_, _31798_);
  and (_39747_, _39746_, _39745_);
  or (_39748_, _39747_, _39670_);
  and (_39749_, _39633_, p3in_reg[7]);
  and (_39750_, _39632_, p3_in[7]);
  or (_39751_, _39750_, _39749_);
  or (_39752_, _39751_, _39631_);
  nand (_39753_, _39631_, _27969_);
  and (_39754_, _39753_, _39752_);
  or (_39755_, _39754_, _37432_);
  and (_39756_, _39755_, _39659_);
  and (_39757_, _39756_, _39748_);
  or (_39758_, _39757_, _39741_);
  and (_39759_, _39633_, p3in_reg[2]);
  and (_39760_, _39632_, p3_in[2]);
  or (_39761_, _39760_, _39759_);
  or (_39762_, _39761_, _39631_);
  nand (_39763_, _39631_, _31634_);
  and (_39764_, _39763_, _39762_);
  or (_39765_, _39764_, _39670_);
  and (_39766_, _39633_, p3in_reg[6]);
  and (_39767_, _39632_, p3_in[6]);
  or (_39768_, _39767_, _39766_);
  or (_39769_, _39768_, _39631_);
  nand (_39770_, _39631_, _32288_);
  and (_39771_, _39770_, _39769_);
  or (_39772_, _39771_, _37432_);
  and (_39773_, _39772_, _39651_);
  and (_39774_, _39773_, _39765_);
  and (_39775_, _39633_, p3in_reg[1]);
  and (_39776_, _39632_, p3_in[1]);
  or (_39777_, _39776_, _39775_);
  or (_39778_, _39777_, _39631_);
  nand (_39779_, _39631_, _31471_);
  and (_39780_, _39779_, _39778_);
  or (_39781_, _39780_, _39670_);
  and (_39782_, _39633_, p3in_reg[5]);
  and (_39783_, _39632_, p3_in[5]);
  or (_39784_, _39783_, _39782_);
  or (_39785_, _39784_, _39631_);
  nand (_39786_, _39631_, _32125_);
  and (_39787_, _39786_, _39785_);
  or (_39788_, _39787_, _37432_);
  and (_39789_, _39788_, _39607_);
  and (_39790_, _39789_, _39781_);
  or (_39791_, _39790_, _39774_);
  or (_39792_, _39791_, _39758_);
  and (_39793_, _39792_, _39545_);
  and (_39794_, _39633_, p2in_reg[0]);
  and (_39795_, _39632_, p2_in[0]);
  or (_39796_, _39795_, _39794_);
  or (_39797_, _39796_, _39631_);
  nand (_39798_, _39631_, _30169_);
  and (_39799_, _39798_, _39797_);
  or (_39800_, _39799_, _39670_);
  and (_39801_, _39633_, p2in_reg[4]);
  and (_39802_, _39632_, p2_in[4]);
  or (_39803_, _39802_, _39801_);
  or (_39804_, _39803_, _39631_);
  nand (_39805_, _39631_, _30817_);
  and (_39806_, _39805_, _39804_);
  or (_39807_, _39806_, _37432_);
  and (_39808_, _39807_, _39642_);
  and (_39809_, _39808_, _39800_);
  and (_39810_, _39633_, p2in_reg[3]);
  and (_39811_, _39632_, p2_in[3]);
  or (_39812_, _39811_, _39810_);
  or (_39813_, _39812_, _39631_);
  nand (_39814_, _39631_, _30655_);
  and (_39815_, _39814_, _39813_);
  or (_39816_, _39815_, _39670_);
  and (_39817_, _39633_, p2in_reg[7]);
  and (_39818_, _39632_, p2_in[7]);
  or (_39819_, _39818_, _39817_);
  or (_39820_, _39819_, _39631_);
  nand (_39821_, _39631_, _27763_);
  and (_39822_, _39821_, _39820_);
  or (_39823_, _39822_, _37432_);
  and (_39824_, _39823_, _39659_);
  and (_39825_, _39824_, _39816_);
  or (_39826_, _39825_, _39809_);
  and (_39827_, _39633_, p2in_reg[2]);
  and (_39828_, _39632_, p2_in[2]);
  or (_39829_, _39828_, _39827_);
  or (_39830_, _39829_, _39631_);
  nand (_39831_, _39631_, _30493_);
  and (_39832_, _39831_, _39830_);
  or (_39833_, _39832_, _39670_);
  and (_39834_, _39633_, p2in_reg[6]);
  and (_39835_, _39632_, p2_in[6]);
  or (_39836_, _39835_, _39834_);
  or (_39837_, _39836_, _39631_);
  nand (_39838_, _39631_, _31143_);
  and (_39839_, _39838_, _39837_);
  or (_39840_, _39839_, _37432_);
  and (_39841_, _39840_, _39651_);
  and (_39842_, _39841_, _39833_);
  and (_39843_, _39633_, p2in_reg[1]);
  and (_39844_, _39632_, p2_in[1]);
  or (_39845_, _39844_, _39843_);
  or (_39846_, _39845_, _39631_);
  nand (_39847_, _39631_, _30331_);
  and (_39848_, _39847_, _39846_);
  or (_39849_, _39848_, _39670_);
  and (_39850_, _39633_, p2in_reg[5]);
  and (_39851_, _39632_, p2_in[5]);
  or (_39852_, _39851_, _39850_);
  or (_39853_, _39852_, _39631_);
  nand (_39854_, _39631_, _30980_);
  and (_39855_, _39854_, _39853_);
  or (_39856_, _39855_, _37432_);
  and (_39857_, _39856_, _39607_);
  and (_39858_, _39857_, _39849_);
  or (_39859_, _39858_, _39842_);
  or (_39860_, _39859_, _39826_);
  and (_39861_, _39860_, _39542_);
  or (_39862_, _39861_, _39793_);
  and (_39863_, _39556_, _39551_);
  or (_39864_, _39670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_39865_, _37432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_39866_, _39865_, _39659_);
  and (_39867_, _39866_, _39864_);
  or (_39868_, _39670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_39869_, _37432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_39870_, _39869_, _39651_);
  and (_39871_, _39870_, _39868_);
  or (_39872_, _39871_, _39867_);
  nand (_39873_, _37432_, _33793_);
  or (_39874_, _37432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_39875_, _39874_, _39642_);
  and (_39876_, _39875_, _39873_);
  or (_39877_, _39670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_39878_, _37432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_39879_, _39878_, _39607_);
  and (_39880_, _39879_, _39877_);
  or (_39881_, _39880_, _39876_);
  or (_39882_, _39881_, _39872_);
  and (_39883_, _39882_, _39863_);
  and (_39884_, _39559_, _39547_);
  and (_39885_, _39884_, _37552_);
  or (_39886_, _39670_, _25478_);
  or (_39887_, _37432_, _25888_);
  and (_39888_, _39887_, _39607_);
  and (_39889_, _39888_, _39886_);
  not (_39890_, _27363_);
  and (_39891_, _39890_, _27222_);
  nor (_39892_, _39890_, _27222_);
  nor (_39893_, _39892_, _39891_);
  not (_39894_, _26366_);
  nor (_39895_, _27070_, _39894_);
  and (_39896_, _27070_, _39894_);
  nor (_39897_, _39896_, _39895_);
  nor (_39898_, _39897_, _39893_);
  and (_39899_, _39897_, _39893_);
  nor (_39900_, _39899_, _39898_);
  not (_39901_, _26539_);
  nor (_39902_, _26658_, _39901_);
  and (_39903_, _26658_, _39901_);
  nor (_39904_, _39903_, _39902_);
  nor (_39905_, _26929_, _26788_);
  and (_39906_, _26929_, _26788_);
  nor (_39907_, _39906_, _39905_);
  nor (_39908_, _39907_, _39904_);
  and (_39909_, _39907_, _39904_);
  or (_39910_, _39909_, _39908_);
  or (_39911_, _39910_, _39900_);
  nand (_39912_, _39910_, _39900_);
  and (_39913_, _39912_, _39911_);
  or (_39914_, _39913_, _39670_);
  or (_39915_, _37432_, _25791_);
  and (_39916_, _39915_, _39642_);
  and (_39917_, _39916_, _39914_);
  or (_39918_, _39917_, _39889_);
  or (_39919_, _39670_, _25619_);
  or (_39920_, _37432_, _26040_);
  and (_39921_, _39920_, _39651_);
  and (_39922_, _39921_, _39919_);
  or (_39923_, _39670_, _25705_);
  or (_39924_, _37432_, _25381_);
  and (_39925_, _39924_, _39659_);
  and (_39926_, _39925_, _39923_);
  or (_39927_, _39926_, _39922_);
  or (_39928_, _39927_, _39918_);
  and (_39929_, _39928_, _39885_);
  or (_39930_, _39929_, _39883_);
  or (_39931_, _39930_, _39862_);
  and (_39932_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_39933_, _39932_, _39670_);
  and (_39934_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_39935_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_39936_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_39937_, _39936_, _39935_);
  or (_39938_, _39937_, _39934_);
  or (_39939_, _39938_, _39933_);
  and (_39940_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_39941_, _39940_, _37432_);
  and (_39942_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_39943_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_39944_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_39945_, _39944_, _39943_);
  or (_39946_, _39945_, _39942_);
  or (_39947_, _39946_, _39941_);
  and (_39948_, _39947_, _39566_);
  and (_39949_, _39948_, _39939_);
  and (_39950_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_39951_, _39950_, _39670_);
  and (_39952_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_39953_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_39954_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_39955_, _39954_, _39953_);
  or (_39956_, _39955_, _39952_);
  or (_39957_, _39956_, _39951_);
  and (_39958_, _39557_, _37395_);
  and (_39959_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_39960_, _39959_, _37432_);
  and (_39961_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_39962_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_39963_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_39964_, _39963_, _39962_);
  or (_39965_, _39964_, _39961_);
  or (_39966_, _39965_, _39960_);
  and (_39967_, _39966_, _39958_);
  and (_39968_, _39967_, _39957_);
  or (_39969_, _39968_, _39949_);
  and (_39970_, _39633_, p0in_reg[2]);
  and (_39971_, _39632_, p0_in[2]);
  or (_39972_, _39971_, _39970_);
  or (_39973_, _39972_, _39631_);
  nand (_39974_, _39631_, _28401_);
  and (_39975_, _39974_, _39973_);
  and (_39976_, _39975_, _39651_);
  and (_39977_, _39633_, p0in_reg[1]);
  and (_39978_, _39632_, p0_in[1]);
  or (_39979_, _39978_, _39977_);
  or (_39980_, _39979_, _39631_);
  or (_39981_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_39982_, _39981_, _39980_);
  and (_39983_, _39982_, _39607_);
  or (_39984_, _39983_, _39976_);
  and (_39985_, _39633_, p0in_reg[3]);
  and (_39986_, _39632_, p0_in[3]);
  or (_39987_, _39986_, _39985_);
  or (_39988_, _39987_, _39631_);
  or (_39989_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_39990_, _39989_, _39988_);
  and (_39991_, _39990_, _39659_);
  and (_39992_, _39633_, p0in_reg[0]);
  and (_39993_, _39632_, p0_in[0]);
  or (_39994_, _39993_, _39992_);
  or (_39995_, _39994_, _39631_);
  nand (_39996_, _39631_, _28142_);
  and (_39997_, _39996_, _39995_);
  and (_39998_, _39997_, _39642_);
  or (_39999_, _39998_, _39991_);
  or (_40000_, _39999_, _39984_);
  and (_40002_, _40000_, _37432_);
  and (_40004_, _39633_, p0in_reg[6]);
  and (_40006_, _39632_, p0_in[6]);
  or (_40008_, _40006_, _40004_);
  or (_40010_, _40008_, _39631_);
  nand (_40012_, _39631_, _29039_);
  and (_40014_, _40012_, _40010_);
  and (_40016_, _40014_, _39651_);
  and (_40018_, _39633_, p0in_reg[5]);
  and (_40020_, _39632_, p0_in[5]);
  or (_40022_, _40020_, _40018_);
  or (_40024_, _40022_, _39631_);
  nand (_40026_, _39631_, _28887_);
  and (_40028_, _40026_, _40024_);
  and (_40030_, _40028_, _39607_);
  or (_40032_, _40030_, _40016_);
  and (_40034_, _39633_, p0in_reg[7]);
  and (_40036_, _39632_, p0_in[7]);
  or (_40038_, _40036_, _40034_);
  or (_40040_, _40038_, _39631_);
  or (_40042_, _39638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_40044_, _40042_, _40040_);
  and (_40046_, _40044_, _39659_);
  and (_40048_, _39633_, p0in_reg[4]);
  and (_40050_, _39632_, p0_in[4]);
  or (_40052_, _40050_, _40048_);
  or (_40054_, _40052_, _39631_);
  nand (_40056_, _39631_, _28736_);
  and (_40058_, _40056_, _40054_);
  and (_40060_, _40058_, _39642_);
  or (_40062_, _40060_, _40046_);
  or (_40063_, _40062_, _40032_);
  and (_40064_, _40063_, _39670_);
  or (_40065_, _40064_, _40002_);
  and (_40066_, _40065_, _39553_);
  and (_40067_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_40068_, _40067_, _39670_);
  and (_40069_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_40070_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_40071_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_40072_, _40071_, _40070_);
  or (_40073_, _40072_, _40069_);
  or (_40074_, _40073_, _40068_);
  and (_40075_, _39607_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_40076_, _40075_, _37432_);
  and (_40077_, _39659_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_40078_, _39642_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_40079_, _39651_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_40080_, _40079_, _40078_);
  or (_40081_, _40080_, _40077_);
  or (_40082_, _40081_, _40076_);
  and (_40083_, _40082_, _39565_);
  and (_40084_, _40083_, _40074_);
  or (_40085_, _40084_, _40066_);
  or (_40086_, _40085_, _39969_);
  or (_40087_, _40086_, _39931_);
  nor (_40088_, _40087_, _39725_);
  nor (_40089_, _40088_, _39605_);
  and (_40090_, _39565_, _26104_);
  and (_40091_, _39605_, ABINPUT[0]);
  or (_40092_, _40091_, _40090_);
  or (_40093_, _40092_, _40089_);
  nor (_40094_, _39631_, _39555_);
  nand (_40095_, _39590_, _25326_);
  or (_40096_, _40095_, _40094_);
  nor (_40097_, _40096_, _39570_);
  nand (_40098_, _39659_, _39894_);
  nand (_40099_, _39642_, _27070_);
  and (_40100_, _40099_, _40098_);
  nand (_40101_, _39651_, _27363_);
  nand (_40102_, _39607_, _27222_);
  and (_40103_, _40102_, _40101_);
  and (_40104_, _40103_, _40100_);
  or (_40105_, _40104_, _37432_);
  nand (_40106_, _39659_, _26929_);
  nand (_40107_, _39642_, _39901_);
  and (_40108_, _40107_, _40106_);
  not (_40109_, _26788_);
  nand (_40110_, _39651_, _40109_);
  not (_40111_, _26658_);
  nand (_40112_, _39607_, _40111_);
  and (_40113_, _40112_, _40110_);
  and (_40114_, _40113_, _40108_);
  or (_40115_, _40114_, _39670_);
  and (_40116_, _40115_, _40090_);
  and (_40117_, _40116_, _40105_);
  nor (_40118_, _40117_, _40097_);
  and (_40119_, _40118_, _40093_);
  and (_40120_, _39607_, ABINPUT[4]);
  and (_40121_, _39659_, ABINPUT[6]);
  or (_40122_, _40121_, _40120_);
  and (_40123_, _39642_, ABINPUT[3]);
  and (_40124_, _39651_, ABINPUT[5]);
  or (_40125_, _40124_, _40123_);
  or (_40126_, _40125_, _40122_);
  and (_40127_, _40126_, _37432_);
  and (_40128_, _39607_, ABINPUT[8]);
  and (_40129_, _39659_, ABINPUT[10]);
  or (_40130_, _40129_, _40128_);
  and (_40131_, _39642_, ABINPUT[7]);
  and (_40132_, _39651_, ABINPUT[9]);
  or (_40133_, _40132_, _40131_);
  or (_40134_, _40133_, _40130_);
  and (_40135_, _40134_, _39670_);
  or (_40136_, _40135_, _40127_);
  and (_40137_, _40136_, _40097_);
  or (_40138_, _40137_, _40119_);
  and (_01522_, _40138_, _39026_);
  and (_40139_, _37552_, _37432_);
  and (_40140_, _40139_, _39642_);
  and (_40141_, _40140_, _39564_);
  and (_40142_, _40141_, _26072_);
  not (_40143_, _25261_);
  and (_40144_, _40140_, _39884_);
  and (_40146_, _40144_, _40143_);
  nor (_40147_, _40146_, _40142_);
  and (_40148_, _40139_, _39659_);
  and (_40149_, _40148_, _39552_);
  nand (_40150_, _40149_, _23971_);
  and (_40151_, _40150_, _40147_);
  nor (_40152_, _40151_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_40153_, _40152_);
  nor (_40154_, _22884_, _16372_);
  and (_40155_, _40154_, _39603_);
  not (_40156_, _40155_);
  and (_40158_, _39642_, _37432_);
  and (_40159_, _40158_, _40090_);
  not (_40160_, _26235_);
  and (_40161_, _39659_, _39670_);
  nor (_40162_, _40161_, _40160_);
  and (_40163_, _40162_, _39590_);
  nor (_40164_, _40163_, _40159_);
  and (_40165_, _40164_, _40156_);
  and (_40166_, _40165_, _40153_);
  and (_40167_, _40139_, _39651_);
  and (_40168_, _40167_, _39552_);
  and (_40169_, _40168_, _23971_);
  or (_40170_, _40169_, rst);
  nor (_01524_, _40170_, _40166_);
  or (_40171_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_40172_, _40158_, _39566_);
  and (_40173_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_40174_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_40175_, _40174_, _40173_);
  and (_40176_, _40158_, _37553_);
  and (_40177_, _40176_, _39552_);
  and (_40178_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_40179_, _40176_, _39541_);
  and (_40180_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_40181_, _40180_, _40178_);
  or (_40182_, _40181_, _40175_);
  and (_40183_, _40140_, _39722_);
  and (_40184_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_40185_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_40186_, _40185_, _40184_);
  and (_40188_, _40139_, _39607_);
  and (_40189_, _40188_, _39552_);
  and (_40190_, _40189_, _37304_);
  and (_40191_, _40140_, _39544_);
  and (_40192_, _40191_, _39754_);
  or (_40193_, _40192_, _40190_);
  or (_40194_, _40193_, _40186_);
  or (_40195_, _40194_, _40182_);
  and (_40196_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_40197_, _40140_, _39541_);
  and (_40198_, _40197_, _39822_);
  and (_40199_, _40140_, _39548_);
  and (_40200_, _40199_, _39698_);
  or (_40201_, _40200_, _40198_);
  and (_40202_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_40203_, _40140_, _39552_);
  and (_40204_, _40203_, _40044_);
  or (_40205_, _40204_, _40202_);
  or (_40206_, _40205_, _40201_);
  or (_40207_, _40206_, _40196_);
  nor (_40209_, _40207_, _40195_);
  nand (_40210_, _40209_, _40166_);
  and (_40211_, _40210_, _40171_);
  or (_40212_, _40211_, _40169_);
  nand (_40213_, _40169_, _24026_);
  and (_40214_, _40213_, _39026_);
  and (_01526_, _40214_, _40212_);
  nor (_01529_, _37354_, rst);
  or (_40215_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_40216_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_40217_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_40218_, _40217_, _40216_);
  and (_40219_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_40220_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_40221_, _40220_, _40219_);
  or (_40222_, _40221_, _40218_);
  and (_40223_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_40224_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_40225_, _40224_, _40223_);
  and (_40226_, _40189_, _37555_);
  and (_40227_, _40191_, _39731_);
  or (_40228_, _40227_, _40226_);
  or (_40229_, _40228_, _40225_);
  or (_40230_, _40229_, _40222_);
  and (_40231_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_40232_, _40197_, _39799_);
  and (_40233_, _40199_, _39648_);
  or (_40234_, _40233_, _40232_);
  and (_40235_, _40203_, _39997_);
  and (_40236_, _40144_, _39913_);
  or (_40237_, _40236_, _40235_);
  or (_40238_, _40237_, _40234_);
  or (_40239_, _40238_, _40231_);
  nor (_40240_, _40239_, _40230_);
  nand (_40241_, _40240_, _40166_);
  and (_40242_, _40241_, _40215_);
  or (_40243_, _40242_, _40169_);
  nand (_40244_, _40169_, _24199_);
  and (_40245_, _40244_, _39026_);
  and (_02205_, _40245_, _40243_);
  or (_40246_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_40247_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_40248_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_40249_, _40248_, _40247_);
  and (_40250_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_40251_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_40252_, _40251_, _40250_);
  or (_40253_, _40252_, _40249_);
  and (_40254_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_40255_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_40256_, _40255_, _40254_);
  and (_40257_, _40189_, _37499_);
  and (_40258_, _40191_, _39780_);
  or (_40259_, _40258_, _40257_);
  or (_40260_, _40259_, _40256_);
  or (_40261_, _40260_, _40253_);
  and (_40262_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_40263_, _40197_, _39848_);
  and (_40264_, _40199_, _39640_);
  or (_40265_, _40264_, _40263_);
  and (_40266_, _40203_, _39982_);
  and (_40267_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_40268_, _40267_, _40266_);
  or (_40269_, _40268_, _40265_);
  or (_40270_, _40269_, _40262_);
  nor (_40271_, _40270_, _40261_);
  nand (_40272_, _40271_, _40166_);
  and (_40273_, _40272_, _40246_);
  or (_40274_, _40273_, _40169_);
  nand (_40275_, _40169_, _24295_);
  and (_40276_, _40275_, _39026_);
  and (_02207_, _40276_, _40274_);
  or (_40277_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_40278_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_40279_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_40280_, _40279_, _40278_);
  and (_40281_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_40282_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_40283_, _40282_, _40281_);
  or (_40284_, _40283_, _40280_);
  and (_40285_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_40286_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_40287_, _40286_, _40285_);
  and (_40288_, _40189_, _37397_);
  and (_40289_, _40191_, _39764_);
  or (_40290_, _40289_, _40288_);
  or (_40291_, _40290_, _40287_);
  or (_40292_, _40291_, _40284_);
  and (_40293_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_40294_, _40197_, _39832_);
  and (_40295_, _40199_, _39657_);
  or (_40296_, _40295_, _40294_);
  and (_40297_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_40298_, _40203_, _39975_);
  or (_40299_, _40298_, _40297_);
  or (_40300_, _40299_, _40296_);
  or (_40301_, _40300_, _40293_);
  nor (_40302_, _40301_, _40292_);
  nand (_40303_, _40302_, _40166_);
  and (_40304_, _40303_, _40277_);
  or (_40305_, _40304_, _40169_);
  nand (_40306_, _40169_, _24392_);
  and (_40307_, _40306_, _39026_);
  and (_02209_, _40307_, _40305_);
  or (_40308_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_40309_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_40310_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_40311_, _40310_, _40309_);
  and (_40312_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_40313_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_40314_, _40313_, _40312_);
  or (_40315_, _40314_, _40311_);
  and (_40316_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_40317_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_40318_, _40317_, _40316_);
  and (_40319_, _40189_, _37517_);
  and (_40320_, _40191_, _39747_);
  or (_40321_, _40320_, _40319_);
  or (_40322_, _40321_, _40318_);
  or (_40323_, _40322_, _40315_);
  and (_40324_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_40325_, _40197_, _39815_);
  and (_40326_, _40199_, _39665_);
  or (_40327_, _40326_, _40325_);
  and (_40328_, _40203_, _39990_);
  and (_40329_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_40330_, _40329_, _40328_);
  or (_40331_, _40330_, _40327_);
  or (_40332_, _40331_, _40324_);
  nor (_40333_, _40332_, _40323_);
  nand (_40334_, _40333_, _40166_);
  and (_40335_, _40334_, _40308_);
  or (_40336_, _40335_, _40169_);
  nand (_40337_, _40169_, _24489_);
  and (_40338_, _40337_, _39026_);
  and (_02211_, _40338_, _40336_);
  or (_40339_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_40340_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_40341_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_40342_, _40341_, _40340_);
  and (_40343_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_40344_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_40345_, _40344_, _40343_);
  or (_40346_, _40345_, _40342_);
  and (_40347_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_40348_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_40349_, _40348_, _40347_);
  and (_40350_, _40189_, _37460_);
  and (_40351_, _40191_, _39738_);
  or (_40352_, _40351_, _40350_);
  or (_40353_, _40352_, _40349_);
  or (_40354_, _40353_, _40346_);
  and (_40355_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_40356_, _40197_, _39806_);
  and (_40357_, _40199_, _39683_);
  or (_40358_, _40357_, _40356_);
  and (_40359_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_40360_, _40203_, _40058_);
  or (_40361_, _40360_, _40359_);
  or (_40362_, _40361_, _40358_);
  or (_40363_, _40362_, _40355_);
  nor (_40364_, _40363_, _40354_);
  nand (_40365_, _40364_, _40166_);
  and (_40366_, _40365_, _40339_);
  or (_40367_, _40366_, _40169_);
  nand (_40368_, _40169_, _24586_);
  and (_40369_, _40368_, _39026_);
  and (_02213_, _40369_, _40367_);
  or (_40370_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_40371_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_40372_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_40373_, _40372_, _40371_);
  and (_40374_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_40375_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_40376_, _40375_, _40374_);
  or (_40377_, _40376_, _40373_);
  and (_40378_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_40379_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_40380_, _40379_, _40378_);
  not (_40381_, _23864_);
  and (_40382_, _40189_, _40381_);
  and (_40383_, _40191_, _39787_);
  or (_40384_, _40383_, _40382_);
  or (_40385_, _40384_, _40380_);
  or (_40386_, _40385_, _40377_);
  and (_40387_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_40388_, _40197_, _39855_);
  and (_40389_, _40199_, _39676_);
  or (_40390_, _40389_, _40388_);
  and (_40391_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_40392_, _40203_, _40028_);
  or (_40393_, _40392_, _40391_);
  or (_40394_, _40393_, _40390_);
  or (_40395_, _40394_, _40387_);
  nor (_40396_, _40395_, _40386_);
  nand (_40397_, _40396_, _40166_);
  and (_40398_, _40397_, _40370_);
  or (_40399_, _40398_, _40169_);
  nand (_40400_, _40169_, _24683_);
  and (_40401_, _40400_, _39026_);
  and (_02215_, _40401_, _40399_);
  or (_40402_, _40166_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_40403_, _40172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_40404_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_40405_, _40404_, _40403_);
  and (_40406_, _40177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_40407_, _40179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_40408_, _40407_, _40406_);
  or (_40409_, _40408_, _40405_);
  and (_40410_, _40183_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_40411_, _40149_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_40412_, _40411_, _40410_);
  and (_40413_, _40189_, _37628_);
  and (_40414_, _40191_, _39771_);
  or (_40415_, _40414_, _40413_);
  or (_40416_, _40415_, _40412_);
  or (_40417_, _40416_, _40409_);
  and (_40418_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_40419_, _40197_, _39839_);
  and (_40420_, _40199_, _39691_);
  or (_40421_, _40420_, _40419_);
  and (_40422_, _40203_, _40014_);
  and (_40423_, _40144_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_40424_, _40423_, _40422_);
  or (_40425_, _40424_, _40421_);
  or (_40426_, _40425_, _40418_);
  nor (_40427_, _40426_, _40417_);
  nand (_40428_, _40427_, _40166_);
  and (_40429_, _40428_, _40402_);
  or (_40430_, _40429_, _40169_);
  nand (_40431_, _40169_, _24780_);
  and (_40432_, _40431_, _39026_);
  and (_02217_, _40432_, _40430_);
  or (_40433_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_40434_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_40435_, _39632_, _40434_);
  and (_40436_, _40435_, _39026_);
  and (_02773_, _40436_, _40433_);
  and (_40437_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_40439_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or (_40440_, _40439_, _40437_);
  and (_02777_, _40440_, _39026_);
  nor (_03155_, _37342_, rst);
  nor (_03162_, _37438_, rst);
  nor (_03166_, _37335_, rst);
  nor (_40442_, ABINPUT[28], ABINPUT[27]);
  nor (_40443_, ABINPUT[30], ABINPUT[29]);
  and (_40444_, _40443_, _40442_);
  nor (_40446_, ABINPUT[32], ABINPUT[31]);
  nor (_40447_, ABINPUT[33], ABINPUT[34]);
  and (_40448_, _40447_, _40446_);
  and (_40449_, _40448_, _40444_);
  not (_40450_, _22643_);
  or (_40452_, _21732_, _21710_);
  and (_40453_, _40452_, _21132_);
  nor (_40454_, _40453_, _22588_);
  nor (_40455_, _40454_, _18609_);
  nor (_40456_, _40454_, _37352_);
  nor (_40458_, _40456_, _40455_);
  and (_40459_, _40458_, _40450_);
  and (_40460_, _40459_, _40449_);
  nor (_40461_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_40462_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_40464_, _40462_, _40461_);
  nor (_40465_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_40466_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_40467_, _40466_, _40465_);
  and (_40468_, _40467_, _40464_);
  and (_40470_, _40468_, _21579_);
  nor (_40471_, _40470_, _40460_);
  and (_40473_, _40458_, _19857_);
  nor (_40474_, _40473_, _40450_);
  nand (_40475_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_40476_, _40475_, _40471_);
  not (_40477_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_40478_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _40477_);
  and (_40479_, _37822_, _37821_);
  and (_40481_, _37792_, _37790_);
  nor (_40482_, _40481_, _40479_);
  and (_40483_, _37764_, _37760_);
  and (_40485_, _37808_, _37807_);
  nor (_40486_, _40485_, _40483_);
  and (_40487_, _40486_, _40482_);
  and (_40489_, _37836_, _37835_);
  and (_40490_, _37776_, _37773_);
  nor (_40491_, _40490_, _40489_);
  and (_40493_, _37738_, _37737_);
  and (_40494_, _37851_, _37850_);
  nor (_40495_, _40494_, _40493_);
  and (_40497_, _40495_, _40491_);
  and (_40498_, _40497_, _40487_);
  nor (_40499_, _40498_, _40478_);
  and (_40501_, _40478_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_40502_, _40501_, _40499_);
  nor (_40503_, _40502_, _40458_);
  not (_40505_, _40503_);
  and (_40506_, _40505_, _40476_);
  and (_40508_, _22632_, _20631_);
  nor (_40509_, _40508_, _22599_);
  or (_40510_, _40509_, _40506_);
  and (_40511_, _21165_, _21132_);
  nor (_40512_, _40511_, _21339_);
  not (_40513_, _40512_);
  and (_40514_, _39612_, _20729_);
  not (_40516_, _40514_);
  and (_40517_, _21776_, _21819_);
  nor (_40518_, _40517_, _22159_);
  and (_40520_, _40518_, _40516_);
  and (_40521_, _39612_, _20685_);
  nor (_40522_, _40521_, _20696_);
  and (_40524_, _40522_, _40520_);
  or (_40525_, _21710_, _21329_);
  or (_40526_, _40525_, _21874_);
  and (_40528_, _40526_, _21132_);
  not (_40529_, _40528_);
  and (_40530_, _40529_, _40524_);
  not (_40532_, _40530_);
  and (_40533_, _40532_, _40506_);
  nor (_40534_, _40533_, _40513_);
  and (_40536_, _40534_, _40510_);
  nor (_40537_, _40536_, _37352_);
  or (_40538_, _21438_, _19606_);
  nor (_40540_, _40538_, _20871_);
  and (_40541_, _21448_, _20347_);
  nor (_40543_, _40541_, _40540_);
  nor (_40544_, _40543_, _18609_);
  nor (_40545_, _40544_, _21590_);
  not (_40546_, _40545_);
  nor (_40547_, _40546_, _40537_);
  not (_40549_, _25196_);
  nor (_40550_, _25337_, _40143_);
  and (_40551_, _40550_, _40549_);
  not (_40553_, _40551_);
  and (_40554_, _40553_, _40474_);
  not (_40555_, _21579_);
  and (_40557_, _26441_, _27167_);
  nor (_40558_, _40557_, _40555_);
  nor (_40559_, _40558_, _40554_);
  not (_40561_, _40559_);
  nor (_40562_, _40561_, _40547_);
  not (_40563_, _40562_);
  nor (_40565_, _22884_, _17145_);
  not (_40566_, _40565_);
  nor (_40567_, _40566_, _40458_);
  and (_40569_, _40567_, _39590_);
  nor (_40570_, _40569_, _40563_);
  and (_40571_, _40570_, _40156_);
  nor (_40573_, _21601_, rst);
  and (_03175_, _40573_, _40571_);
  and (_03179_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39026_);
  and (_03182_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39026_);
  not (_40575_, _39418_);
  not (_40576_, _40456_);
  and (_40577_, _40522_, _40518_);
  nor (_40578_, _40577_, _37352_);
  not (_40579_, _40578_);
  and (_40581_, _21132_, _22731_);
  and (_40582_, _40581_, _20838_);
  not (_40583_, _40582_);
  and (_40585_, _21547_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_40586_, _40585_, _21459_);
  and (_40587_, _40541_, _22731_);
  nor (_40589_, _40587_, _40586_);
  and (_40590_, _40589_, _40583_);
  and (_40591_, _40590_, _40579_);
  and (_40593_, _40591_, _40576_);
  nor (_40594_, _40593_, _40575_);
  and (_40595_, _40593_, _37299_);
  nor (_40597_, _40595_, _40594_);
  and (_40598_, _40597_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_40599_, _40597_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_40601_, _39537_);
  nor (_40602_, _40593_, _40601_);
  and (_40603_, _40593_, _37611_);
  nor (_40605_, _40603_, _40602_);
  and (_40606_, _40605_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_40608_, _40605_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_40609_, _40608_, _40606_);
  not (_40610_, _39520_);
  nor (_40611_, _40593_, _40610_);
  and (_40613_, _40593_, _37383_);
  nor (_40614_, _40613_, _40611_);
  and (_40615_, _40614_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_40617_, _40614_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_40618_, _39503_);
  nor (_40619_, _40593_, _40618_);
  and (_40621_, _40593_, _37455_);
  nor (_40622_, _40621_, _40619_);
  nand (_40623_, _40622_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_40625_, _39486_);
  nor (_40626_, _40593_, _40625_);
  and (_40627_, _40593_, _37547_);
  nor (_40629_, _40627_, _40626_);
  and (_40630_, _40629_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_40631_, _40629_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_40633_, _39469_);
  nor (_40634_, _40593_, _40633_);
  and (_40635_, _40593_, _37427_);
  nor (_40637_, _40635_, _40634_);
  and (_40638_, _40637_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_40640_, _39452_);
  nor (_40641_, _40593_, _40640_);
  and (_40642_, _40593_, _37494_);
  nor (_40643_, _40642_, _40641_);
  and (_40645_, _40643_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_40646_, _39435_);
  nor (_40647_, _40593_, _40646_);
  and (_40649_, _40593_, _37585_);
  nor (_40650_, _40649_, _40647_);
  and (_40651_, _40650_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_40653_, _40643_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_40654_, _40653_, _40645_);
  and (_40655_, _40654_, _40651_);
  nor (_40657_, _40655_, _40645_);
  not (_40658_, _40657_);
  nor (_40659_, _40637_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_40661_, _40659_, _40638_);
  and (_40662_, _40661_, _40658_);
  nor (_40663_, _40662_, _40638_);
  nor (_40665_, _40663_, _40631_);
  or (_40666_, _40665_, _40630_);
  or (_40667_, _40622_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_40669_, _40667_, _40623_);
  nand (_40670_, _40669_, _40666_);
  and (_40672_, _40670_, _40623_);
  nor (_40673_, _40672_, _40617_);
  or (_40674_, _40673_, _40615_);
  and (_40675_, _40674_, _40609_);
  nor (_40677_, _40675_, _40606_);
  nor (_40678_, _40677_, _40599_);
  or (_40679_, _40678_, _40598_);
  and (_40681_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_40682_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_40683_, _40682_, _40681_);
  and (_40685_, _40683_, _40679_);
  and (_40686_, _40685_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_40687_, _40686_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_40689_, _40687_, _40597_);
  not (_40690_, _40597_);
  not (_40691_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_40693_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_40694_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_40695_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_40697_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_40698_, _40679_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_40699_, _40698_, _40697_);
  and (_40701_, _40699_, _40695_);
  and (_40702_, _40701_, _40694_);
  and (_40704_, _40702_, _40693_);
  and (_40705_, _40704_, _40691_);
  nor (_40706_, _40705_, _40690_);
  nor (_40707_, _40706_, _40689_);
  or (_40708_, _40597_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_40709_, _40597_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_40710_, _40709_, _40708_);
  and (_40712_, _40710_, _40707_);
  or (_40713_, _40712_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_40714_, _40712_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_40716_, _40524_, _40512_);
  and (_40717_, _40716_, _21557_);
  and (_40718_, _22577_, _22731_);
  nor (_40720_, _40718_, _22643_);
  and (_40721_, _40720_, _40576_);
  not (_40722_, _40721_);
  nor (_40724_, _40722_, _40717_);
  and (_40725_, _21557_, _21339_);
  nor (_40726_, _40725_, _40544_);
  not (_40728_, _40726_);
  and (_40729_, _40728_, _40593_);
  nor (_40730_, _40729_, _40724_);
  and (_40732_, _40730_, _40714_);
  and (_40733_, _40732_, _40713_);
  and (_40734_, _40724_, _40591_);
  and (_40736_, _40734_, _40726_);
  and (_40737_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_40739_, _40725_, ABINPUT[18]);
  and (_40740_, _21601_, ABINPUT[26]);
  or (_40741_, _40740_, _40739_);
  or (_40742_, _40741_, _40737_);
  and (_40744_, _40587_, _37300_);
  and (_40745_, _40734_, _40728_);
  and (_40746_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_40748_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_40749_, _40748_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_40750_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_40752_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_40753_, _40752_, _40750_);
  and (_40754_, _40753_, _40749_);
  and (_40756_, _40754_, _40683_);
  and (_40757_, _40756_, _40746_);
  and (_40758_, _40757_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_40760_, _40758_, _40434_);
  and (_40761_, _40758_, _40434_);
  or (_40762_, _40761_, _40760_);
  and (_40764_, _40762_, _40745_);
  or (_40765_, _40764_, _40744_);
  nor (_40766_, _40765_, _40742_);
  nand (_40768_, _40766_, _40571_);
  or (_40769_, _40768_, _40733_);
  nor (_40771_, _18784_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_40772_, _40771_, _37283_);
  nor (_40773_, _40772_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_40774_, _40773_);
  and (_40776_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_40777_, _40776_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_40778_, _40777_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_40780_, _40778_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_40781_, _40780_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_40782_, _40781_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_40784_, _40782_, _40774_);
  and (_40785_, _40784_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_40786_, _40785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_40788_, _40786_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_40789_, _40788_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_40790_, _40789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_40792_, _40790_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_40793_, _40792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_40794_, _40792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_40796_, _40794_, _40793_);
  or (_40797_, _40796_, _40571_);
  and (_40798_, _40797_, _39026_);
  and (_03185_, _40798_, _40769_);
  and (_40800_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39026_);
  and (_40802_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_40803_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_40804_, _18653_, _40803_);
  not (_40805_, _40804_);
  not (_40807_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_40808_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_40809_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_40811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_40812_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_40813_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_40815_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_40816_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_40817_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_40819_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_40820_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_40821_, _40820_, _40819_);
  and (_40823_, _40821_, _40817_);
  and (_40824_, _40823_, _40816_);
  and (_40825_, _40824_, _40815_);
  and (_40827_, _40825_, _40813_);
  and (_40828_, _40827_, _40812_);
  and (_40829_, _40828_, _40811_);
  and (_40831_, _40829_, _40809_);
  and (_40832_, _40831_, _40808_);
  nor (_40834_, _40832_, _40807_);
  and (_40835_, _40832_, _40807_);
  nor (_40836_, _40835_, _40834_);
  nor (_40837_, _40831_, _40808_);
  or (_40838_, _40837_, _40832_);
  and (_40840_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_40841_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_40842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_40844_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_40845_, _40844_, _40841_);
  and (_40846_, _40845_, _40842_);
  nor (_40848_, _40846_, _40841_);
  nor (_40849_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_40850_, _40849_, _40840_);
  not (_40852_, _40850_);
  nor (_40853_, _40852_, _40848_);
  nor (_40854_, _40853_, _40840_);
  not (_40856_, _40854_);
  and (_40857_, _40856_, _40828_);
  and (_40858_, _40857_, _40811_);
  and (_40860_, _40858_, _40809_);
  and (_40861_, _40860_, _40838_);
  nor (_40862_, _40860_, _40838_);
  or (_40864_, _40862_, _40861_);
  not (_40865_, _40864_);
  and (_40867_, _40854_, _40831_);
  and (_40868_, _40854_, _40829_);
  nor (_40869_, _40868_, _40809_);
  nor (_40870_, _40869_, _40867_);
  not (_40872_, _40870_);
  and (_40873_, _40854_, _40828_);
  and (_40874_, _40854_, _40825_);
  and (_40876_, _40874_, _40813_);
  nor (_40877_, _40876_, _40812_);
  nor (_40878_, _40877_, _40873_);
  not (_40880_, _40878_);
  nor (_40881_, _40874_, _40813_);
  or (_40882_, _40881_, _40876_);
  not (_40884_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_40885_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_40886_, _40854_, _40824_);
  and (_40888_, _40886_, _40885_);
  nor (_40889_, _40888_, _40884_);
  nor (_40890_, _40889_, _40874_);
  not (_40892_, _40890_);
  and (_40893_, _40854_, _40821_);
  and (_40894_, _40893_, _40817_);
  nor (_40896_, _40894_, _40816_);
  nor (_40897_, _40896_, _40886_);
  not (_40899_, _40897_);
  nor (_40900_, _40893_, _40817_);
  nor (_40901_, _40900_, _40894_);
  not (_40902_, _40901_);
  and (_40904_, _40854_, _40820_);
  nor (_40905_, _40904_, _40819_);
  nor (_40906_, _40905_, _40893_);
  not (_40908_, _40906_);
  not (_40909_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_40910_, _40854_, _40909_);
  nor (_40912_, _40854_, _40909_);
  nor (_40913_, _40912_, _40910_);
  not (_40914_, _40913_);
  not (_40916_, _21089_);
  and (_40917_, _19286_, _19046_);
  and (_40918_, _40917_, _19584_);
  and (_40920_, _40918_, _40916_);
  not (_40921_, _20075_);
  and (_40922_, _20304_, _40921_);
  not (_40924_, _20598_);
  and (_40925_, _40924_, _19835_);
  and (_40926_, _40925_, _40922_);
  and (_40928_, _40926_, _40920_);
  nor (_40929_, _40916_, _19584_);
  and (_40931_, _40929_, _40917_);
  not (_40932_, _20304_);
  and (_40933_, _40932_, _20075_);
  and (_40934_, _20598_, _19835_);
  and (_40936_, _40934_, _40933_);
  and (_40937_, _40936_, _40931_);
  nor (_40938_, _40937_, _40928_);
  and (_40940_, _40925_, _40933_);
  and (_40941_, _40940_, _40931_);
  not (_40942_, _19835_);
  and (_40944_, _20598_, _40942_);
  and (_40945_, _40944_, _40922_);
  nor (_40946_, _19584_, _19286_);
  and (_40948_, _40946_, _19046_);
  and (_40949_, _40948_, _21089_);
  and (_40950_, _40949_, _40945_);
  nor (_40952_, _40950_, _40941_);
  and (_40953_, _40952_, _40938_);
  and (_40954_, _40948_, _40916_);
  not (_40956_, _40954_);
  nor (_40957_, _20304_, _20075_);
  and (_40958_, _40925_, _40957_);
  nor (_40960_, _40958_, _40936_);
  nor (_40961_, _40960_, _40956_);
  not (_40962_, _40961_);
  nor (_40963_, _21089_, _19584_);
  and (_40964_, _40963_, _40917_);
  and (_40965_, _40936_, _40949_);
  nor (_40966_, _40965_, _40964_);
  and (_40967_, _40966_, _40962_);
  and (_40968_, _40967_, _40953_);
  nor (_40969_, _40940_, _40945_);
  nor (_40970_, _40969_, _40956_);
  and (_40971_, _40918_, _21089_);
  and (_40972_, _20304_, _20075_);
  and (_40973_, _40972_, _19835_);
  and (_40974_, _40973_, _40971_);
  nor (_40975_, _40974_, _40970_);
  not (_40976_, _40971_);
  and (_40977_, _40944_, _40933_);
  nor (_40978_, _40958_, _40977_);
  nor (_40979_, _40978_, _40976_);
  and (_40980_, _40972_, _40942_);
  and (_40981_, _40980_, _40954_);
  nor (_40982_, _40981_, _40979_);
  and (_40983_, _40982_, _40975_);
  and (_40984_, _40983_, _40968_);
  and (_40985_, _40977_, _40949_);
  and (_40986_, _40957_, _40934_);
  and (_40987_, _40954_, _40986_);
  nor (_40988_, _40925_, _40944_);
  and (_40989_, _40972_, _40931_);
  and (_40990_, _40989_, _40988_);
  or (_40991_, _40990_, _40987_);
  nor (_40992_, _40991_, _40985_);
  not (_40993_, _40931_);
  nor (_40994_, _20598_, _19835_);
  and (_40995_, _40933_, _40994_);
  nor (_40996_, _20075_, _40942_);
  and (_40997_, _40996_, _40932_);
  nor (_40998_, _40997_, _40995_);
  nor (_40999_, _40998_, _40993_);
  nor (_41000_, _40971_, _40948_);
  and (_41001_, _40934_, _40922_);
  not (_41002_, _41001_);
  nor (_41003_, _41002_, _41000_);
  nor (_41004_, _41003_, _40999_);
  and (_41005_, _41004_, _40992_);
  nor (_41006_, _40945_, _40995_);
  nor (_41007_, _41006_, _19046_);
  not (_41008_, _19046_);
  and (_41009_, _40986_, _41008_);
  nor (_41010_, _41009_, _41007_);
  and (_41011_, _40980_, _40949_);
  not (_41012_, _41011_);
  and (_41013_, _40957_, _40994_);
  and (_41014_, _41013_, _40954_);
  and (_41015_, _40926_, _40931_);
  nor (_41016_, _41015_, _41014_);
  and (_41017_, _41016_, _41012_);
  and (_41018_, _41017_, _41010_);
  and (_41019_, _41018_, _41005_);
  and (_41020_, _41019_, _40984_);
  and (_41021_, _40922_, _40942_);
  and (_41022_, _40931_, _41021_);
  not (_41023_, _41022_);
  and (_41024_, _40971_, _40940_);
  and (_41025_, _40977_, _40931_);
  nor (_41026_, _41025_, _41024_);
  and (_41027_, _41026_, _41023_);
  and (_41028_, _40940_, _41008_);
  or (_41029_, _40922_, _40933_);
  not (_41030_, _19286_);
  and (_41031_, _19584_, _41030_);
  and (_41032_, _41031_, _19046_);
  and (_41033_, _41032_, _40944_);
  and (_41034_, _41033_, _41029_);
  nor (_41035_, _41034_, _41028_);
  and (_41036_, _40977_, _41008_);
  and (_41037_, _40933_, _40924_);
  and (_41038_, _41032_, _41037_);
  nor (_41039_, _41038_, _41036_);
  and (_41040_, _41039_, _41035_);
  and (_41041_, _41040_, _41027_);
  and (_41042_, _40957_, _40944_);
  and (_41043_, _41042_, _40954_);
  nor (_41044_, _41043_, _40926_);
  nor (_41045_, _41044_, _41000_);
  not (_41046_, _41045_);
  and (_41047_, _40922_, _40994_);
  not (_41048_, _41047_);
  nor (_41049_, _40948_, _40918_);
  nor (_41050_, _41049_, _41048_);
  nor (_41051_, _40986_, _40945_);
  nor (_41052_, _41051_, _40976_);
  nor (_41053_, _41052_, _41050_);
  and (_41054_, _41053_, _41046_);
  and (_41055_, _40977_, _40954_);
  and (_41056_, _41001_, _40920_);
  or (_41057_, _41056_, _41055_);
  and (_41058_, _40973_, _40954_);
  nor (_41059_, _41058_, _41057_);
  nor (_41060_, _40936_, _40995_);
  nor (_41061_, _41060_, _40976_);
  and (_41062_, _40972_, _40944_);
  nor (_41063_, _41062_, _41001_);
  nor (_41064_, _41063_, _40993_);
  nor (_41065_, _41064_, _41061_);
  and (_41066_, _41065_, _41059_);
  and (_41067_, _41066_, _41054_);
  and (_41068_, _41067_, _41041_);
  and (_41069_, _41068_, _41020_);
  nor (_41070_, _40845_, _40842_);
  nor (_41071_, _41070_, _40846_);
  not (_41072_, _41071_);
  nor (_41073_, _41072_, _41069_);
  not (_41074_, _41057_);
  and (_41075_, _40975_, _41074_);
  and (_41076_, _40920_, _41047_);
  not (_41077_, _41076_);
  and (_41078_, _41062_, _40931_);
  or (_41079_, _41031_, _41008_);
  and (_41080_, _41079_, _40977_);
  nor (_41081_, _41080_, _41078_);
  and (_41082_, _41081_, _41077_);
  and (_41083_, _41082_, _40938_);
  and (_41084_, _41083_, _41075_);
  and (_41085_, _41084_, _40992_);
  not (_41086_, _41085_);
  nor (_41087_, _41086_, _41069_);
  not (_41088_, _41087_);
  nor (_41089_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_41090_, _41089_, _40842_);
  and (_41091_, _41090_, _41088_);
  and (_41092_, _41072_, _41069_);
  nor (_41093_, _41092_, _41073_);
  and (_41094_, _41093_, _41091_);
  nor (_41095_, _41094_, _41073_);
  not (_41096_, _41095_);
  and (_41097_, _40852_, _40848_);
  nor (_41098_, _41097_, _40853_);
  and (_41099_, _41098_, _41096_);
  and (_41100_, _41099_, _40914_);
  not (_41101_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_41102_, _40910_, _41101_);
  or (_41103_, _41102_, _40904_);
  and (_41104_, _41103_, _41100_);
  and (_41105_, _41104_, _40908_);
  and (_41106_, _41105_, _40902_);
  and (_41107_, _41106_, _40899_);
  nor (_41108_, _40886_, _40885_);
  or (_41109_, _41108_, _40888_);
  and (_41110_, _41109_, _41107_);
  and (_41111_, _41110_, _40892_);
  and (_41112_, _41111_, _40882_);
  and (_41113_, _41112_, _40880_);
  nor (_41114_, _40873_, _40811_);
  or (_41115_, _41114_, _40868_);
  and (_41116_, _41115_, _41113_);
  and (_41117_, _41116_, _40872_);
  and (_41118_, _41117_, _40865_);
  or (_41119_, _41118_, _40861_);
  nor (_41120_, _41119_, _40836_);
  and (_41121_, _41119_, _40836_);
  or (_41122_, _41121_, _41120_);
  or (_41123_, _41122_, _40805_);
  or (_41124_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_41125_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_41126_, _41125_, _41124_);
  and (_41127_, _41126_, _41123_);
  or (_03188_, _41127_, _40802_);
  nor (_41128_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_03193_, _41128_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_03196_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39026_);
  not (_41129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  not (_41130_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_41131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_41132_, _41131_, _41130_);
  nor (_41133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_41134_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_41135_, _41134_, _41133_);
  and (_41136_, _41135_, _41132_);
  and (_41137_, _41136_, _41129_);
  and (_41138_, \oc8051_top_1.oc8051_rom1.ea_int , _18620_);
  nand (_41139_, _41138_, _18653_);
  nand (_41140_, _41139_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_41141_, _41140_, _41137_);
  and (_03199_, _41141_, _39026_);
  and (_41142_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_41143_, _41142_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_03202_, _41143_, _39026_);
  nor (_41144_, _40773_, _37283_);
  nor (_41145_, _41069_, _18871_);
  nor (_41146_, _41087_, _18827_);
  and (_41147_, _41069_, _18871_);
  nor (_41148_, _41147_, _41145_);
  and (_41149_, _41148_, _41146_);
  nor (_41150_, _41149_, _41145_);
  nor (_41151_, _41150_, _37283_);
  and (_41152_, _41151_, _18740_);
  nor (_41153_, _41151_, _18740_);
  nor (_41154_, _41153_, _41152_);
  nor (_41155_, _41154_, _41144_);
  and (_41156_, _18882_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_41157_, _41156_, _41144_);
  nor (_41158_, _41157_, _41085_);
  or (_41159_, _41158_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_41160_, _41159_, _41155_);
  and (_03204_, _41160_, _39026_);
  not (_41161_, _19508_);
  and (_41162_, _20031_, _41161_);
  not (_41163_, _20533_);
  and (_41164_, _41163_, _20260_);
  and (_41165_, _41164_, _41162_);
  and (_41166_, _18653_, _39026_);
  and (_41167_, _41166_, _18642_);
  nand (_41168_, _41167_, _19242_);
  nor (_41169_, _41168_, _19002_);
  not (_41170_, _21045_);
  and (_41171_, _41170_, _19792_);
  and (_41172_, _41171_, _41169_);
  and (_03212_, _41172_, _41165_);
  not (_41173_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_41174_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_41175_, _41174_, _41173_);
  or (_41176_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_41177_, _41176_, _39026_);
  and (_03214_, _41177_, _41175_);
  and (_03217_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _39026_);
  not (_41178_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_41179_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_41180_, _41179_, _41178_);
  and (_41181_, _41179_, _41178_);
  nor (_41182_, _41181_, _41180_);
  not (_41183_, _41182_);
  and (_41184_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_41185_, _41184_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_41186_, _41184_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_41187_, _41186_, _41185_);
  or (_41188_, _41187_, _41179_);
  and (_41189_, _41188_, _41183_);
  nor (_41190_, _41180_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_41191_, _41180_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_41192_, _41191_, _41190_);
  or (_41193_, _41185_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03223_, _41193_, _39026_);
  and (_41194_, _03223_, _41192_);
  and (_03220_, _41194_, _41189_);
  not (_41195_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_41196_, _40773_, _41195_);
  and (_41197_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_41198_, _41196_);
  and (_41199_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_41200_, _41199_, _41197_);
  and (_03226_, _41200_, _39026_);
  and (_41201_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_41202_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_41203_, _41202_, _41201_);
  and (_03228_, _41203_, _39026_);
  and (_41204_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_41205_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_41206_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _41205_);
  and (_41207_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_41208_, _41207_, _41204_);
  and (_03230_, _41208_, _39026_);
  and (_41209_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_41210_, _41209_, _41206_);
  and (_03232_, _41210_, _39026_);
  or (_41211_, _41205_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_03234_, _41211_, _39026_);
  not (_41212_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_41213_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_41214_, _41213_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_41215_, _41205_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_41216_, _41215_, _39026_);
  and (_03236_, _41216_, _41214_);
  or (_41217_, _41205_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_03238_, _41217_, _39026_);
  nor (_41218_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_41220_, _41218_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_41221_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_41222_, _41221_, _41220_);
  and (_03240_, _41222_, _39026_);
  and (_41223_, _41195_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_41224_, _41223_, _41220_);
  and (_03242_, _41224_, _39026_);
  or (_41225_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  nand (_41226_, _41220_, _24069_);
  and (_41227_, _41226_, _39026_);
  and (_03244_, _41227_, _41225_);
  and (_03246_, _22863_, _37337_);
  or (_41229_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_41230_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_41231_, _39632_, _41230_);
  and (_41232_, _41231_, _39026_);
  and (_03627_, _41232_, _41229_);
  or (_41233_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_41234_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_41235_, _39632_, _41234_);
  and (_41237_, _41235_, _39026_);
  and (_03629_, _41237_, _41233_);
  or (_41238_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_41239_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_41240_, _39632_, _41239_);
  and (_41241_, _41240_, _39026_);
  and (_03631_, _41241_, _41238_);
  or (_41242_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_41243_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_41244_, _39632_, _41243_);
  and (_41246_, _41244_, _39026_);
  and (_03633_, _41246_, _41242_);
  or (_41247_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_41248_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_41249_, _39632_, _41248_);
  and (_41250_, _41249_, _39026_);
  and (_03635_, _41250_, _41247_);
  or (_41251_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_41252_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_41253_, _39632_, _41252_);
  and (_41255_, _41253_, _39026_);
  and (_03637_, _41255_, _41251_);
  or (_41256_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_41257_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_41258_, _39632_, _41257_);
  and (_41259_, _41258_, _39026_);
  and (_03639_, _41259_, _41256_);
  or (_41260_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_41261_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_41262_, _39632_, _41261_);
  and (_41264_, _41262_, _39026_);
  and (_03641_, _41264_, _41260_);
  or (_41265_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_41266_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_41267_, _39632_, _41266_);
  and (_41268_, _41267_, _39026_);
  and (_03643_, _41268_, _41265_);
  or (_41269_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_41270_, _39632_, _40697_);
  and (_41271_, _41270_, _39026_);
  and (_03645_, _41271_, _41269_);
  or (_41273_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_41274_, _39632_, _40695_);
  and (_41275_, _41274_, _39026_);
  and (_03647_, _41275_, _41273_);
  or (_41276_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_41277_, _39632_, _40694_);
  and (_41278_, _41277_, _39026_);
  and (_03649_, _41278_, _41276_);
  or (_41279_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_41281_, _39632_, _40693_);
  and (_41282_, _41281_, _39026_);
  and (_03651_, _41282_, _41279_);
  or (_41283_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_41284_, _39632_, _40691_);
  and (_41285_, _41284_, _39026_);
  and (_03653_, _41285_, _41283_);
  or (_41286_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  not (_41287_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_41288_, _39632_, _41287_);
  and (_41290_, _41288_, _39026_);
  and (_03655_, _41290_, _41286_);
  and (_41291_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_41292_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_41293_, _41292_, _41291_);
  and (_03687_, _41293_, _39026_);
  and (_41294_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_41295_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_41296_, _41295_, _41294_);
  and (_03689_, _41296_, _39026_);
  and (_41298_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_41299_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_41300_, _41299_, _41298_);
  and (_03691_, _41300_, _39026_);
  and (_41301_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_41302_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_41303_, _41302_, _41301_);
  and (_03693_, _41303_, _39026_);
  and (_41304_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_41305_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_41307_, _41305_, _41304_);
  and (_03695_, _41307_, _39026_);
  and (_41308_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_41309_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_41310_, _41309_, _41308_);
  and (_03697_, _41310_, _39026_);
  and (_41311_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_41312_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_41313_, _41312_, _41311_);
  and (_03699_, _41313_, _39026_);
  and (_41315_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_41316_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_41317_, _41316_, _41315_);
  and (_03701_, _41317_, _39026_);
  and (_41318_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_41319_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_41320_, _41319_, _41318_);
  and (_03703_, _41320_, _39026_);
  and (_41321_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_41322_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_41324_, _41322_, _41321_);
  and (_03705_, _41324_, _39026_);
  and (_41325_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_41326_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_41327_, _41326_, _41325_);
  and (_03707_, _41327_, _39026_);
  and (_41328_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_41329_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_41330_, _41329_, _41328_);
  and (_03709_, _41330_, _39026_);
  and (_41332_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_41333_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_41334_, _41333_, _41332_);
  and (_03711_, _41334_, _39026_);
  and (_41335_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_41336_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_41337_, _41336_, _41335_);
  and (_03713_, _41337_, _39026_);
  and (_41338_, _39633_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_41339_, _39632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_41340_, _41339_, _41338_);
  and (_03715_, _41340_, _39026_);
  and (_41341_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_41342_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_41343_, _41342_, _41341_);
  and (_05587_, _41343_, _39026_);
  and (_41344_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_41345_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_41346_, _41345_, _41196_);
  or (_41347_, _41346_, _41344_);
  and (_05589_, _41347_, _39026_);
  and (_41348_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_41349_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_41350_, _41349_, _41196_);
  or (_41351_, _41350_, _41348_);
  and (_05591_, _41351_, _39026_);
  and (_41352_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_41353_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_41354_, _41353_, _41352_);
  and (_05593_, _41354_, _39026_);
  and (_41355_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_41356_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_41357_, _41356_, _41196_);
  or (_41358_, _41357_, _41355_);
  and (_05595_, _41358_, _39026_);
  and (_41359_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_41360_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_41361_, _41360_, _41196_);
  or (_41362_, _41361_, _41359_);
  and (_05597_, _41362_, _39026_);
  and (_41363_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_41364_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_41365_, _41364_, _41196_);
  or (_41366_, _41365_, _41363_);
  and (_05599_, _41366_, _39026_);
  and (_41367_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_41368_, _41196_, _41174_);
  or (_41369_, _41368_, _41367_);
  and (_05601_, _41369_, _39026_);
  and (_41370_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_41371_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_41372_, _41371_, _41370_);
  and (_05603_, _41372_, _39026_);
  and (_41373_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_41374_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_41375_, _41374_, _41373_);
  and (_05605_, _41375_, _39026_);
  and (_41376_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_41377_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_41378_, _41377_, _41376_);
  and (_05607_, _41378_, _39026_);
  and (_41379_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_41380_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_41381_, _41380_, _41379_);
  and (_05609_, _41381_, _39026_);
  and (_41382_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_41383_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_41384_, _41383_, _41382_);
  and (_05611_, _41384_, _39026_);
  and (_41385_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_41386_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_41387_, _41386_, _41385_);
  and (_05613_, _41387_, _39026_);
  and (_41388_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_41389_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_41390_, _41389_, _41388_);
  and (_05615_, _41390_, _39026_);
  and (_41391_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_41392_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_41393_, _41392_, _41391_);
  and (_05617_, _41393_, _39026_);
  and (_41394_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_41395_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_41396_, _41395_, _41394_);
  and (_05619_, _41396_, _39026_);
  and (_41397_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_41398_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_41399_, _41398_, _41397_);
  and (_05621_, _41399_, _39026_);
  and (_41400_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_41401_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_41402_, _41401_, _41400_);
  and (_05623_, _41402_, _39026_);
  and (_41403_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_41404_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_41405_, _41404_, _41403_);
  and (_05625_, _41405_, _39026_);
  and (_41406_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_41407_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_41408_, _41407_, _41406_);
  and (_05627_, _41408_, _39026_);
  and (_41409_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_41410_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_41411_, _41410_, _41409_);
  and (_05629_, _41411_, _39026_);
  and (_41412_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_41413_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_41414_, _41413_, _41412_);
  and (_05631_, _41414_, _39026_);
  and (_41415_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_41416_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_41417_, _41416_, _41415_);
  and (_05633_, _41417_, _39026_);
  and (_41418_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_41419_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_41420_, _41419_, _41418_);
  and (_05635_, _41420_, _39026_);
  and (_41421_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_41422_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_41423_, _41422_, _41421_);
  and (_05637_, _41423_, _39026_);
  and (_41424_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_41425_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_41426_, _41425_, _41424_);
  and (_05639_, _41426_, _39026_);
  and (_41427_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_41428_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_41429_, _41428_, _41427_);
  and (_05641_, _41429_, _39026_);
  and (_41430_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_41431_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_41432_, _41431_, _41430_);
  and (_05643_, _41432_, _39026_);
  and (_41433_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_41434_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_41435_, _41434_, _41433_);
  and (_05645_, _41435_, _39026_);
  and (_41436_, _41196_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_41437_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_41438_, _41437_, _41436_);
  and (_05647_, _41438_, _39026_);
  and (_05650_, _21111_, _39026_);
  and (_05653_, _19606_, _39026_);
  and (_05656_, _19318_, _39026_);
  nor (_05658_, _37314_, rst);
  nor (_05661_, _37569_, rst);
  nor (_05664_, _37510_, rst);
  nor (_05667_, _37411_, rst);
  nor (_05670_, _37531_, rst);
  nor (_05673_, _37471_, rst);
  nor (_05676_, _37366_, rst);
  nor (_05679_, _37625_, rst);
  and (_05709_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39026_);
  and (_05711_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39026_);
  and (_05713_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39026_);
  and (_05715_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39026_);
  and (_05717_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39026_);
  and (_05719_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39026_);
  and (_05721_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39026_);
  or (_41439_, _40736_, _40725_);
  and (_41440_, _41439_, ABINPUT[19]);
  and (_41441_, _40745_, _37586_);
  and (_41442_, _40587_, _40646_);
  and (_41443_, _21601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_41444_, _41443_, _41442_);
  or (_41445_, _41444_, _41441_);
  or (_41446_, _41445_, _41440_);
  nor (_41447_, _21765_, _37352_);
  not (_41448_, _40522_);
  nor (_41449_, _41448_, _22632_);
  and (_41450_, _41449_, _40512_);
  and (_41451_, _41450_, _40520_);
  nor (_41452_, _41451_, _37352_);
  nor (_41453_, _41452_, _41447_);
  and (_41454_, _41453_, _40583_);
  nor (_41455_, _41454_, _40729_);
  nor (_41456_, _40650_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_41457_, _41456_, _40651_);
  and (_41458_, _41457_, _41455_);
  nor (_41459_, _41458_, _41446_);
  nand (_41460_, _41459_, _40571_);
  or (_41461_, _40571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_41462_, _41461_, _39026_);
  and (_05723_, _41462_, _41460_);
  and (_41463_, _41439_, ABINPUT[20]);
  and (_41464_, _40745_, _37495_);
  and (_41465_, _40587_, _40640_);
  and (_41466_, _21601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_41467_, _41466_, _41465_);
  or (_41468_, _41467_, _41464_);
  or (_41469_, _41468_, _41463_);
  nor (_41470_, _40654_, _40651_);
  nor (_41471_, _41470_, _40655_);
  and (_41472_, _41471_, _41455_);
  nor (_41473_, _41472_, _41469_);
  nand (_41474_, _41473_, _40571_);
  or (_41475_, _40571_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_41476_, _41475_, _39026_);
  and (_05725_, _41476_, _41474_);
  and (_41477_, _40586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_41478_, _41439_, ABINPUT[21]);
  and (_41479_, _40745_, _37428_);
  and (_41480_, _40587_, _40633_);
  or (_41481_, _41480_, _41479_);
  or (_41482_, _41481_, _41478_);
  nor (_41483_, _40661_, _40658_);
  nor (_41484_, _41483_, _40662_);
  and (_41485_, _41484_, _41455_);
  or (_41486_, _41485_, _41482_);
  or (_41487_, _41486_, _41477_);
  and (_41488_, _41487_, _40571_);
  not (_41489_, _40571_);
  not (_41490_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_41491_, _40773_, _41490_);
  and (_41492_, _40773_, _41490_);
  nor (_41493_, _41492_, _41491_);
  and (_41494_, _41493_, _41489_);
  or (_41495_, _41494_, _41488_);
  and (_05727_, _41495_, _39026_);
  and (_41496_, _40586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_41497_, _41439_, ABINPUT[22]);
  and (_41498_, _40587_, _40625_);
  and (_41499_, _40745_, _37548_);
  or (_41500_, _41499_, _41498_);
  or (_41501_, _41500_, _41497_);
  or (_41502_, _41501_, _41496_);
  or (_41503_, _40631_, _40630_);
  or (_41504_, _41503_, _40663_);
  nand (_41505_, _41503_, _40663_);
  and (_41506_, _41505_, _41504_);
  and (_41507_, _41506_, _41455_);
  or (_41508_, _41507_, _41502_);
  and (_41509_, _41508_, _40571_);
  and (_41510_, _41491_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_41511_, _41491_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_41512_, _41511_, _41510_);
  and (_41513_, _41512_, _41489_);
  or (_41514_, _41513_, _41509_);
  and (_05729_, _41514_, _39026_);
  or (_41515_, _40669_, _40666_);
  and (_41516_, _40730_, _40670_);
  and (_41517_, _41516_, _41515_);
  and (_41518_, _41439_, ABINPUT[23]);
  and (_41519_, _40587_, _40618_);
  and (_41520_, _40745_, _37456_);
  and (_41521_, _21601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_41522_, _41521_, _41520_);
  or (_41523_, _41522_, _41519_);
  or (_41524_, _41523_, _41518_);
  or (_41525_, _41524_, _41517_);
  and (_41526_, _41525_, _40571_);
  and (_41527_, _41491_, _40776_);
  nor (_41528_, _41510_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_41529_, _41528_, _41527_);
  nor (_41530_, _41529_, _40571_);
  or (_41531_, _41530_, _41526_);
  and (_05731_, _41531_, _39026_);
  and (_41532_, _40586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_41533_, _41439_, ABINPUT[24]);
  and (_41534_, _40587_, _40610_);
  and (_41535_, _40745_, _37384_);
  or (_41536_, _41535_, _41534_);
  or (_41537_, _41536_, _41533_);
  or (_41538_, _41537_, _41532_);
  or (_41539_, _40617_, _40615_);
  or (_41540_, _41539_, _40672_);
  nand (_41541_, _41539_, _40672_);
  and (_41542_, _41541_, _40730_);
  and (_41543_, _41542_, _41540_);
  or (_41544_, _41543_, _41538_);
  and (_41545_, _41544_, _40571_);
  and (_41546_, _41527_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_41547_, _41527_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_41548_, _41547_, _41546_);
  nor (_41549_, _41548_, _40571_);
  or (_41550_, _41549_, _41545_);
  and (_05733_, _41550_, _39026_);
  and (_41551_, _40586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_41552_, _41439_, ABINPUT[25]);
  and (_41553_, _40745_, _37612_);
  and (_41554_, _40587_, _40601_);
  or (_41555_, _41554_, _41553_);
  or (_41556_, _41555_, _41552_);
  nor (_41557_, _40674_, _40609_);
  nor (_41558_, _41557_, _40675_);
  and (_41559_, _41558_, _41455_);
  or (_41560_, _41559_, _41556_);
  or (_41561_, _41560_, _41551_);
  and (_41562_, _41561_, _40571_);
  and (_41563_, _41546_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_41564_, _41546_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_41565_, _41564_, _41563_);
  nor (_41566_, _41565_, _40571_);
  or (_41567_, _41566_, _41562_);
  and (_05735_, _41567_, _39026_);
  and (_41568_, _41439_, ABINPUT[26]);
  and (_41569_, _40745_, _37300_);
  and (_41570_, _40587_, _40575_);
  or (_41571_, _41570_, _41569_);
  or (_41572_, _41571_, _41568_);
  or (_41573_, _40598_, _40599_);
  nand (_41574_, _41573_, _40677_);
  or (_41575_, _41573_, _40677_);
  and (_41576_, _41575_, _41574_);
  and (_41577_, _41576_, _41455_);
  or (_41578_, _41577_, _41572_);
  nand (_41579_, _40586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nand (_41580_, _41579_, _40571_);
  or (_41581_, _41580_, _41578_);
  and (_41582_, _40781_, _40774_);
  nor (_41583_, _41563_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_41584_, _41583_, _41582_);
  or (_41585_, _41584_, _40571_);
  and (_41586_, _41585_, _39026_);
  and (_05737_, _41586_, _41581_);
  and (_41587_, _40679_, _41266_);
  nor (_41588_, _40679_, _41266_);
  nor (_41589_, _41588_, _41587_);
  or (_41590_, _41589_, _40690_);
  nand (_41591_, _41589_, _40690_);
  and (_41592_, _41591_, _40730_);
  and (_41593_, _41592_, _41590_);
  and (_41594_, _40587_, _37586_);
  and (_41595_, _40725_, ABINPUT[11]);
  and (_41596_, _21601_, ABINPUT[19]);
  or (_41597_, _41596_, _41595_);
  nor (_41598_, _41597_, _41594_);
  and (_41599_, _40745_, _40942_);
  and (_41600_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_41601_, _41600_, _41599_);
  and (_41602_, _41601_, _41598_);
  nand (_41603_, _41602_, _40571_);
  or (_41604_, _41603_, _41593_);
  nor (_41605_, _41582_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_41606_, _41605_, _40784_);
  or (_41607_, _41606_, _40571_);
  and (_41608_, _41607_, _39026_);
  and (_05739_, _41608_, _41604_);
  and (_41609_, _40679_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_41610_, _41609_, _40690_);
  and (_41611_, _40698_, _40597_);
  nor (_41612_, _41611_, _41610_);
  nand (_41613_, _41612_, _40697_);
  or (_41614_, _41612_, _40697_);
  and (_41615_, _41614_, _40730_);
  and (_41616_, _41615_, _41613_);
  and (_41624_, _40587_, _37495_);
  and (_41631_, _40725_, ABINPUT[12]);
  and (_41635_, _21601_, ABINPUT[20]);
  or (_41641_, _41635_, _41631_);
  nor (_41649_, _41641_, _41624_);
  and (_41654_, _40745_, _40921_);
  and (_41658_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_41666_, _41658_, _41654_);
  and (_41673_, _41666_, _41649_);
  nand (_41677_, _41673_, _40571_);
  or (_41683_, _41677_, _41616_);
  nor (_41691_, _40784_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_41696_, _41691_, _40785_);
  or (_41700_, _41696_, _40571_);
  and (_41708_, _41700_, _39026_);
  and (_05741_, _41708_, _41683_);
  and (_41718_, _40699_, _40597_);
  and (_41724_, _41610_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_41732_, _41724_, _41718_);
  nand (_41737_, _41732_, _40695_);
  or (_41741_, _41732_, _40695_);
  and (_41749_, _41741_, _40730_);
  and (_41756_, _41749_, _41737_);
  and (_41760_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_41766_, _40725_, ABINPUT[13]);
  and (_41774_, _21601_, ABINPUT[21]);
  or (_41779_, _41774_, _41766_);
  nor (_41783_, _41779_, _41760_);
  and (_41791_, _40745_, _40932_);
  and (_41792_, _40587_, _37428_);
  nor (_41801_, _41792_, _41791_);
  and (_41809_, _41801_, _41783_);
  nand (_41816_, _41809_, _40571_);
  or (_41820_, _41816_, _41756_);
  nor (_41826_, _40785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_41834_, _41826_, _40786_);
  or (_41839_, _41834_, _40571_);
  and (_41843_, _41839_, _39026_);
  and (_05743_, _41843_, _41820_);
  and (_41844_, _40681_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_41845_, _41844_, _40679_);
  and (_41846_, _41845_, _40690_);
  and (_41847_, _40701_, _40597_);
  nor (_41848_, _41847_, _41846_);
  nand (_41849_, _41848_, _40694_);
  or (_41850_, _41848_, _40694_);
  and (_41851_, _41850_, _40730_);
  and (_41852_, _41851_, _41849_);
  and (_41853_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_41854_, _40725_, ABINPUT[14]);
  and (_41855_, _21601_, ABINPUT[22]);
  or (_41856_, _41855_, _41854_);
  or (_41857_, _41856_, _41853_);
  and (_41858_, _40587_, _37548_);
  and (_41859_, _40754_, _41844_);
  and (_41860_, _41859_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_41861_, _41859_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_41862_, _41861_, _41860_);
  and (_41863_, _41862_, _40745_);
  or (_41864_, _41863_, _41858_);
  nor (_41865_, _41864_, _41857_);
  nand (_41866_, _41865_, _40571_);
  or (_41867_, _41866_, _41852_);
  nor (_41868_, _40786_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_41869_, _41868_, _40788_);
  or (_41870_, _41869_, _40571_);
  and (_41871_, _41870_, _39026_);
  and (_05745_, _41871_, _41867_);
  and (_41872_, _40702_, _40597_);
  and (_41873_, _40685_, _40690_);
  nor (_41874_, _41873_, _41872_);
  nand (_41875_, _41874_, _40693_);
  or (_41876_, _41874_, _40693_);
  and (_41877_, _41876_, _40730_);
  and (_41878_, _41877_, _41875_);
  and (_41879_, _41860_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_41880_, _41860_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_41881_, _41880_, _41879_);
  and (_41882_, _41881_, _40745_);
  and (_41883_, _40725_, ABINPUT[15]);
  and (_41884_, _21601_, ABINPUT[23]);
  or (_41885_, _41884_, _41883_);
  nor (_41886_, _41885_, _41882_);
  and (_41887_, _40587_, _37456_);
  and (_41888_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_41889_, _41888_, _41887_);
  and (_41890_, _41889_, _41886_);
  nand (_41891_, _41890_, _40571_);
  or (_41892_, _41891_, _41878_);
  nor (_41893_, _40788_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_41894_, _41893_, _40789_);
  or (_41895_, _41894_, _40571_);
  and (_41896_, _41895_, _39026_);
  and (_05747_, _41896_, _41892_);
  and (_41897_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_41898_, _40587_, _37384_);
  and (_41899_, _40586_, ABINPUT[24]);
  or (_41900_, _41899_, _41898_);
  or (_41901_, _41900_, _41897_);
  and (_41902_, _40704_, _40597_);
  and (_41903_, _40686_, _40690_);
  nor (_41904_, _41903_, _41902_);
  nor (_41905_, _41904_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_41906_, _41904_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_41907_, _41906_, _41905_);
  and (_41908_, _41907_, _41455_);
  or (_41909_, _41908_, _41901_);
  and (_41910_, _41879_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_41911_, _41879_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_41912_, _41911_, _41910_);
  and (_41913_, _41912_, _40745_);
  and (_41914_, _40725_, ABINPUT[16]);
  nor (_41915_, _41914_, _41913_);
  nand (_41916_, _41915_, _40571_);
  or (_41917_, _41916_, _41909_);
  nor (_41918_, _40789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_41919_, _41918_, _40790_);
  or (_41920_, _41919_, _40571_);
  and (_41921_, _41920_, _39026_);
  and (_05749_, _41921_, _41917_);
  nand (_41922_, _40725_, ABINPUT[17]);
  nand (_41923_, _40586_, ABINPUT[25]);
  nand (_41924_, _40587_, _37612_);
  and (_41925_, _41924_, _41923_);
  and (_41926_, _41925_, _41922_);
  nand (_41927_, _40736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_41928_, _40757_, _41287_);
  nor (_41929_, _40757_, _41287_);
  or (_41930_, _41929_, _41928_);
  nand (_41931_, _41930_, _40745_);
  and (_41932_, _41931_, _41927_);
  and (_41933_, _40707_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_41934_, _40707_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_41935_, _41934_, _41933_);
  nand (_41936_, _41935_, _41455_);
  and (_41937_, _41936_, _41932_);
  and (_41938_, _41937_, _41926_);
  nand (_41939_, _41938_, _40571_);
  nor (_41940_, _40790_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_41941_, _41940_, _40792_);
  or (_41942_, _41941_, _40571_);
  and (_41943_, _41942_, _39026_);
  and (_05751_, _41943_, _41939_);
  or (_41944_, _41090_, _41088_);
  nor (_41945_, _40805_, _41091_);
  and (_41946_, _41945_, _41944_);
  nor (_41947_, _40804_, _41230_);
  or (_41948_, _41947_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_41949_, _41948_, _41946_);
  or (_41950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _18620_);
  and (_41951_, _41950_, _39026_);
  and (_05753_, _41951_, _41949_);
  and (_41952_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_41953_, _41093_, _41091_);
  nor (_41954_, _41953_, _41094_);
  or (_41955_, _41954_, _40805_);
  or (_41956_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_41957_, _41956_, _41125_);
  and (_41958_, _41957_, _41955_);
  or (_05755_, _41958_, _41952_);
  and (_41959_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_41960_, _41098_, _41096_);
  nor (_41961_, _41960_, _41099_);
  or (_41962_, _41961_, _40805_);
  or (_41963_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_41964_, _41963_, _41125_);
  and (_41965_, _41964_, _41962_);
  or (_05757_, _41965_, _41959_);
  and (_41966_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_41967_, _41099_, _40914_);
  nor (_41968_, _41967_, _41100_);
  or (_41969_, _41968_, _40805_);
  or (_41970_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_41971_, _41970_, _41125_);
  and (_41972_, _41971_, _41969_);
  or (_05759_, _41972_, _41966_);
  and (_41973_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_41974_, _41103_, _41100_);
  nor (_41975_, _41974_, _41104_);
  or (_41976_, _41975_, _40805_);
  or (_41977_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_41978_, _41977_, _41125_);
  and (_41979_, _41978_, _41976_);
  or (_05761_, _41979_, _41973_);
  and (_41980_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_41981_, _41104_, _40908_);
  nor (_41982_, _41981_, _41105_);
  or (_41983_, _41982_, _40805_);
  or (_41984_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_41985_, _41984_, _41125_);
  and (_41986_, _41985_, _41983_);
  or (_05763_, _41986_, _41980_);
  nor (_41987_, _41105_, _40902_);
  nor (_41988_, _41987_, _41106_);
  or (_41989_, _41988_, _40805_);
  or (_41990_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_41991_, _41990_, _41125_);
  and (_41992_, _41991_, _41989_);
  and (_41993_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_05765_, _41993_, _41992_);
  nor (_41994_, _41106_, _40899_);
  nor (_41995_, _41994_, _41107_);
  or (_41996_, _41995_, _40805_);
  or (_41997_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_41998_, _41997_, _41125_);
  and (_41999_, _41998_, _41996_);
  and (_42000_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_05767_, _42000_, _41999_);
  nor (_42001_, _41109_, _41107_);
  nor (_42002_, _42001_, _41110_);
  or (_42003_, _42002_, _40805_);
  or (_42004_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_42005_, _42004_, _41125_);
  and (_42006_, _42005_, _42003_);
  and (_42007_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_05769_, _42007_, _42006_);
  nor (_42008_, _41110_, _40892_);
  nor (_42009_, _42008_, _41111_);
  or (_42010_, _42009_, _40805_);
  or (_42011_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_42012_, _42011_, _41125_);
  and (_42013_, _42012_, _42010_);
  and (_42014_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_05771_, _42014_, _42013_);
  nor (_42015_, _41111_, _40882_);
  nor (_42016_, _42015_, _41112_);
  or (_42017_, _42016_, _40805_);
  or (_42018_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_42019_, _42018_, _41125_);
  and (_42020_, _42019_, _42017_);
  and (_42021_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_05773_, _42021_, _42020_);
  nor (_42022_, _41112_, _40880_);
  nor (_42023_, _42022_, _41113_);
  or (_42024_, _42023_, _40805_);
  or (_42025_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_42026_, _42025_, _41125_);
  and (_42027_, _42026_, _42024_);
  and (_42028_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_05775_, _42028_, _42027_);
  or (_42029_, _41115_, _41113_);
  nor (_42030_, _40805_, _41116_);
  and (_42031_, _42030_, _42029_);
  nor (_42032_, _40804_, _40693_);
  or (_42033_, _42032_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_42034_, _42033_, _42031_);
  or (_42035_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _18620_);
  and (_42036_, _42035_, _39026_);
  and (_05777_, _42036_, _42034_);
  nor (_42037_, _41116_, _40872_);
  nor (_42038_, _42037_, _41117_);
  or (_42039_, _42038_, _40805_);
  or (_42040_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_42041_, _42040_, _41125_);
  and (_42042_, _42041_, _42039_);
  and (_42043_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_05779_, _42043_, _42042_);
  and (_42044_, _40800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_42045_, _41117_, _40865_);
  nor (_42046_, _42045_, _41118_);
  or (_42047_, _42046_, _40805_);
  or (_42048_, _40804_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_42049_, _42048_, _41125_);
  and (_42050_, _42049_, _42047_);
  or (_05781_, _42050_, _42044_);
  and (_42051_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_42052_, _42051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_05783_, _42052_, _39026_);
  and (_42053_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_42054_, _42053_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_05785_, _42054_, _39026_);
  and (_42055_, _41136_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_42056_, _42055_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_05787_, _42056_, _39026_);
  and (_42057_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_42058_, _42057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_05789_, _42058_, _39026_);
  and (_42059_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_42060_, _42059_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_05791_, _42060_, _39026_);
  and (_42061_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_42062_, _42061_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_05793_, _42062_, _39026_);
  and (_42063_, _41137_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_42064_, _42063_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_05795_, _42064_, _39026_);
  nor (_42065_, _41087_, _37283_);
  nand (_42066_, _42065_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_42067_, _42065_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_42068_, _42067_, _41125_);
  and (_05797_, _42068_, _42066_);
  nor (_42069_, _41148_, _41146_);
  nor (_42070_, _42069_, _41149_);
  or (_42071_, _42070_, _37283_);
  or (_42072_, _18653_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_42073_, _42072_, _41125_);
  and (_05799_, _42073_, _42071_);
  and (_42074_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_42075_, _42074_, _41173_);
  or (_42076_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42077_, _42076_, _39026_);
  and (_05829_, _42077_, _42075_);
  or (_42078_, _41345_, _41173_);
  or (_42079_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42080_, _42079_, _39026_);
  and (_05831_, _42080_, _42078_);
  or (_42081_, _41349_, _41173_);
  or (_42082_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42083_, _42082_, _39026_);
  and (_05833_, _42083_, _42081_);
  and (_42084_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_42085_, _42084_, _41173_);
  or (_42086_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42087_, _42086_, _39026_);
  and (_05835_, _42087_, _42085_);
  or (_42088_, _41356_, _41173_);
  or (_42089_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42090_, _42089_, _39026_);
  and (_05837_, _42090_, _42088_);
  or (_42091_, _41360_, _41173_);
  or (_42092_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42093_, _42092_, _39026_);
  and (_05839_, _42093_, _42091_);
  or (_42094_, _41364_, _41173_);
  or (_42095_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_42096_, _42095_, _39026_);
  and (_05841_, _42096_, _42094_);
  and (_05843_, _41182_, _39026_);
  nor (_05845_, _41192_, rst);
  and (_05847_, _41188_, _39026_);
  and (_42097_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_42098_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_42099_, _42098_, _42097_);
  and (_05849_, _42099_, _39026_);
  and (_42100_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_42101_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_42102_, _42101_, _42100_);
  and (_05851_, _42102_, _39026_);
  and (_42103_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_42104_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_42105_, _42104_, _42103_);
  and (_05853_, _42105_, _39026_);
  and (_42106_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_42107_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_42108_, _42107_, _42106_);
  and (_05855_, _42108_, _39026_);
  and (_42109_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_42110_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_42111_, _42110_, _42109_);
  and (_05857_, _42111_, _39026_);
  and (_42112_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_42113_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_42114_, _42113_, _42112_);
  and (_05859_, _42114_, _39026_);
  and (_42115_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_42116_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_42117_, _42116_, _42115_);
  and (_05861_, _42117_, _39026_);
  and (_42118_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_42119_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_42120_, _42119_, _42118_);
  and (_05863_, _42120_, _39026_);
  and (_42121_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_42122_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_42123_, _42122_, _42121_);
  and (_05865_, _42123_, _39026_);
  and (_42124_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_42125_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_42126_, _42125_, _42124_);
  and (_05867_, _42126_, _39026_);
  and (_42127_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_42128_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_42129_, _42128_, _42127_);
  and (_05869_, _42129_, _39026_);
  and (_42130_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_42131_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_42132_, _42131_, _42130_);
  and (_05871_, _42132_, _39026_);
  and (_42133_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_42134_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_42135_, _42134_, _42133_);
  and (_05873_, _42135_, _39026_);
  and (_42136_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_42137_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_42138_, _42137_, _42136_);
  and (_05875_, _42138_, _39026_);
  and (_42139_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_42140_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_42141_, _42140_, _42139_);
  and (_05877_, _42141_, _39026_);
  and (_42142_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_42143_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_42144_, _42143_, _42142_);
  and (_05879_, _42144_, _39026_);
  and (_42145_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_42146_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_42147_, _42146_, _42145_);
  and (_05881_, _42147_, _39026_);
  and (_42148_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_42149_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_42150_, _42149_, _42148_);
  and (_05883_, _42150_, _39026_);
  and (_42151_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_42152_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_42153_, _42152_, _42151_);
  and (_05885_, _42153_, _39026_);
  and (_42154_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_42155_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_42156_, _42155_, _42154_);
  and (_05887_, _42156_, _39026_);
  and (_42157_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_42158_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_42159_, _42158_, _42157_);
  and (_05889_, _42159_, _39026_);
  and (_42160_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_42161_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_42162_, _42161_, _42160_);
  and (_05891_, _42162_, _39026_);
  and (_42163_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_42164_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_42165_, _42164_, _42163_);
  and (_05893_, _42165_, _39026_);
  and (_42166_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_42167_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_42168_, _42167_, _42166_);
  and (_05895_, _42168_, _39026_);
  and (_42169_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_42170_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_42171_, _42170_, _42169_);
  and (_05897_, _42171_, _39026_);
  and (_42172_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_42173_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_42174_, _42173_, _42172_);
  and (_05899_, _42174_, _39026_);
  and (_42175_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_42176_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_42177_, _42176_, _42175_);
  and (_05901_, _42177_, _39026_);
  and (_42178_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_42179_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_42180_, _42179_, _42178_);
  and (_05903_, _42180_, _39026_);
  and (_42181_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_42182_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_42183_, _42182_, _42181_);
  and (_05905_, _42183_, _39026_);
  and (_42184_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_42185_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_42186_, _42185_, _42184_);
  and (_05907_, _42186_, _39026_);
  and (_42187_, _41196_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_42188_, _41198_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_42189_, _42188_, _42187_);
  and (_05909_, _42189_, _39026_);
  and (_42190_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42191_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_42192_, _42191_, _42190_);
  and (_05911_, _42192_, _39026_);
  and (_42193_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42194_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_42195_, _42194_, _42193_);
  and (_05913_, _42195_, _39026_);
  and (_42196_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42197_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_42198_, _42197_, _42196_);
  and (_05915_, _42198_, _39026_);
  and (_42199_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42200_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_42201_, _42200_, _42199_);
  and (_05917_, _42201_, _39026_);
  and (_42202_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42203_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_42204_, _42203_, _42202_);
  and (_05919_, _42204_, _39026_);
  and (_42205_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42206_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_42207_, _42206_, _42205_);
  and (_05921_, _42207_, _39026_);
  and (_42208_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_42209_, _41206_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_42210_, _42209_, _42208_);
  and (_05923_, _42210_, _39026_);
  and (_42211_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42212_, _37569_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42213_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_42214_, _42213_, _41205_);
  and (_42215_, _42214_, _42212_);
  or (_42216_, _42215_, _42211_);
  and (_05925_, _42216_, _39026_);
  and (_42217_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42218_, _37510_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42219_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_42220_, _42219_, _41205_);
  and (_42221_, _42220_, _42218_);
  or (_42222_, _42221_, _42217_);
  and (_05927_, _42222_, _39026_);
  and (_42223_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42224_, _37411_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42225_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_42226_, _42225_, _41205_);
  and (_42227_, _42226_, _42224_);
  or (_42228_, _42227_, _42223_);
  and (_05929_, _42228_, _39026_);
  and (_42229_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42230_, _37531_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42231_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_42232_, _42231_, _41205_);
  and (_42233_, _42232_, _42230_);
  or (_42234_, _42233_, _42229_);
  and (_05931_, _42234_, _39026_);
  and (_42235_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42236_, _37471_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42237_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_42238_, _42237_, _41205_);
  and (_42239_, _42238_, _42236_);
  or (_42240_, _42239_, _42235_);
  and (_05933_, _42240_, _39026_);
  and (_42241_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42242_, _37366_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42243_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_42244_, _42243_, _41205_);
  and (_42245_, _42244_, _42242_);
  or (_42246_, _42245_, _42241_);
  and (_05935_, _42246_, _39026_);
  and (_42247_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42248_, _37625_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42249_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_42250_, _42249_, _41205_);
  and (_42251_, _42250_, _42248_);
  or (_42252_, _42251_, _42247_);
  and (_05937_, _42252_, _39026_);
  and (_42253_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_42254_, _37335_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_42255_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_42256_, _42255_, _41205_);
  and (_42257_, _42256_, _42254_);
  or (_42258_, _42257_, _42253_);
  and (_05939_, _42258_, _39026_);
  and (_42259_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_42260_, _42259_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42261_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _41205_);
  and (_42262_, _42261_, _39026_);
  and (_05941_, _42262_, _42260_);
  and (_42263_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_42264_, _42263_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42265_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _41205_);
  and (_42266_, _42265_, _39026_);
  and (_05943_, _42266_, _42264_);
  and (_42267_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_42268_, _42267_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42269_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _41205_);
  and (_42270_, _42269_, _39026_);
  and (_05945_, _42270_, _42268_);
  and (_42271_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_42272_, _42271_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42273_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _41205_);
  and (_42274_, _42273_, _39026_);
  and (_05947_, _42274_, _42272_);
  and (_42275_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_42276_, _42275_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42277_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _41205_);
  and (_42278_, _42277_, _39026_);
  and (_05949_, _42278_, _42276_);
  and (_42279_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_42280_, _42279_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42281_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _41205_);
  and (_42282_, _42281_, _39026_);
  and (_05951_, _42282_, _42280_);
  and (_42283_, _41212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_42284_, _42283_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_42285_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _41205_);
  and (_42286_, _42285_, _39026_);
  and (_05953_, _42286_, _42284_);
  not (_42287_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_42288_, _41220_, _42287_);
  and (_42289_, _41220_, ABINPUT[19]);
  or (_42290_, _42289_, _42288_);
  and (_05955_, _42290_, _39026_);
  not (_42291_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_42292_, _41220_, _42291_);
  and (_42293_, _41220_, ABINPUT[20]);
  or (_42294_, _42293_, _42292_);
  and (_05957_, _42294_, _39026_);
  not (_42295_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_42296_, _41220_, _42295_);
  and (_42297_, _41220_, ABINPUT[21]);
  or (_42298_, _42297_, _42296_);
  and (_05959_, _42298_, _39026_);
  not (_42299_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_42300_, _41220_, _42299_);
  and (_42301_, _41220_, ABINPUT[22]);
  or (_42302_, _42301_, _42300_);
  and (_05961_, _42302_, _39026_);
  or (_42303_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  nand (_42304_, _41220_, _24586_);
  and (_42305_, _42304_, _39026_);
  and (_05963_, _42305_, _42303_);
  or (_42306_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  nand (_42307_, _41220_, _24683_);
  and (_42308_, _42307_, _39026_);
  and (_05965_, _42308_, _42306_);
  or (_42309_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  nand (_42310_, _41220_, _24780_);
  and (_42311_, _42310_, _39026_);
  and (_05967_, _42311_, _42309_);
  or (_42312_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  nand (_42313_, _41220_, _24026_);
  and (_42314_, _42313_, _39026_);
  and (_05969_, _42314_, _42312_);
  or (_42315_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  nand (_42316_, _41220_, _24242_);
  and (_42317_, _42316_, _39026_);
  and (_05971_, _42317_, _42315_);
  or (_42318_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  nand (_42319_, _41220_, _24339_);
  and (_42320_, _42319_, _39026_);
  and (_05973_, _42320_, _42318_);
  or (_42321_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  nand (_42322_, _41220_, _24436_);
  and (_42323_, _42322_, _39026_);
  and (_05975_, _42323_, _42321_);
  or (_42324_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  nand (_42325_, _41220_, _24533_);
  and (_42326_, _42325_, _39026_);
  and (_05977_, _42326_, _42324_);
  or (_42327_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  nand (_42328_, _41220_, _24630_);
  and (_42329_, _42328_, _39026_);
  and (_05979_, _42329_, _42327_);
  or (_42330_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  nand (_42331_, _41220_, _24726_);
  and (_42332_, _42331_, _39026_);
  and (_05981_, _42332_, _42330_);
  or (_42333_, _41220_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  nand (_42334_, _41220_, _24823_);
  and (_42335_, _42334_, _39026_);
  and (_05983_, _42335_, _42333_);
  and (_08307_, _37689_, _39026_);
  and (_08310_, _37744_, _39026_);
  nor (_08316_, _37432_, rst);
  and (_08467_, _37766_, _39026_);
  and (_08469_, _37783_, _39026_);
  and (_08471_, _37799_, _39026_);
  and (_08473_, _37814_, _39026_);
  and (_08475_, _37829_, _39026_);
  and (_08477_, _37843_, _39026_);
  and (_08479_, _37858_, _39026_);
  nor (_08481_, _37590_, rst);
  nor (_08483_, _37514_, rst);
  nor (_12308_, _22830_, rst);
  nand (_42336_, _41166_, _21383_);
  nor (_42337_, _21230_, _21132_);
  or (_12311_, _42337_, _42336_);
  and (_42338_, _40949_, _41037_);
  and (_42339_, _40920_, _40945_);
  or (_42340_, _42339_, _42338_);
  and (_42341_, _41062_, _40971_);
  or (_42342_, _42341_, _41009_);
  or (_42343_, _42342_, _42340_);
  and (_42344_, _40977_, _40948_);
  or (_42345_, _41015_, _40987_);
  or (_42346_, _42345_, _42344_);
  or (_42347_, _42346_, _42343_);
  and (_42348_, _40972_, _40994_);
  and (_42349_, _42348_, _40971_);
  and (_42350_, _40933_, _19835_);
  and (_42351_, _42350_, _40920_);
  or (_42352_, _42351_, _42349_);
  and (_42353_, _40957_, _40942_);
  and (_42354_, _42353_, _40918_);
  or (_42355_, _42354_, _42352_);
  and (_42356_, _42353_, _40931_);
  or (_42357_, _42356_, _41080_);
  or (_42358_, _42357_, _40990_);
  or (_42359_, _41022_, _40974_);
  or (_42360_, _41064_, _40941_);
  or (_42361_, _42360_, _42359_);
  or (_42362_, _42361_, _42358_);
  or (_42363_, _42362_, _40964_);
  or (_42364_, _42363_, _42355_);
  or (_42365_, _42364_, _42347_);
  and (_42366_, _42365_, _18664_);
  not (_42367_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_42368_, _18642_, _15686_);
  and (_42369_, _42368_, _21536_);
  nor (_42370_, _42369_, _42367_);
  or (_42371_, _42370_, rst);
  or (_12313_, _42371_, _42366_);
  nand (_42372_, _20304_, _18598_);
  or (_42373_, _18598_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_42374_, _42373_, _39026_);
  and (_12316_, _42374_, _42372_);
  and (_42375_, \oc8051_top_1.oc8051_sfr1.wait_data , _39026_);
  and (_42376_, _42375_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_42377_, _21241_, _21143_);
  or (_42378_, _42377_, _22335_);
  nor (_42379_, _42378_, _22137_);
  nand (_42380_, _42379_, _21765_);
  and (_42381_, _22742_, _21797_);
  and (_42382_, _21241_, _21165_);
  or (_42383_, _42382_, _42381_);
  and (_42384_, _22126_, _21241_);
  or (_42385_, _42384_, _40511_);
  or (_42386_, _42385_, _22632_);
  or (_42387_, _42386_, _42383_);
  or (_42388_, _42387_, _42380_);
  and (_42389_, _42388_, _41166_);
  or (_12319_, _42389_, _42376_);
  and (_42390_, _21132_, _20762_);
  or (_42391_, _42390_, _21274_);
  and (_42392_, _22126_, _21776_);
  and (_42393_, _22368_, _20729_);
  or (_42394_, _42393_, _20740_);
  or (_42395_, _42394_, _42392_);
  or (_42396_, _42395_, _42391_);
  and (_42397_, _42396_, _18653_);
  nor (_42398_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42399_, _42398_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_42400_, _22775_);
  and (_42401_, _42400_, _42399_);
  and (_42402_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42403_, _42402_, _42401_);
  or (_42404_, _42403_, _42397_);
  and (_12321_, _42404_, _39026_);
  and (_42405_, _42375_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_42406_, _21732_, _21776_);
  and (_42407_, _22742_, _21961_);
  or (_42408_, _21972_, _22159_);
  or (_42409_, _42408_, _42407_);
  or (_42410_, _42409_, _42406_);
  or (_42411_, _40521_, _39625_);
  or (_42412_, _42411_, _42410_);
  and (_42413_, _22742_, _20762_);
  and (_42414_, _22742_, _21819_);
  or (_42415_, _42414_, _20707_);
  or (_42416_, _42415_, _42391_);
  or (_42417_, _42416_, _42413_);
  or (_42418_, _42417_, _42412_);
  and (_42419_, _42418_, _41166_);
  or (_12324_, _42419_, _42405_);
  and (_42420_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42421_, _22456_, _18653_);
  or (_42422_, _42421_, _42420_);
  or (_42423_, _42422_, _42401_);
  and (_12327_, _42423_, _39026_);
  and (_42424_, _21241_, _20751_);
  not (_42425_, _21797_);
  nor (_42426_, _42337_, _42425_);
  nor (_42427_, _42426_, _42424_);
  not (_42428_, _42427_);
  and (_42429_, _42428_, _42399_);
  or (_42430_, _42429_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42431_, _21732_, _21448_);
  and (_42432_, _40540_, _20620_);
  or (_42433_, _42432_, _42431_);
  or (_42434_, _42433_, _42382_);
  and (_42435_, _42433_, _21557_);
  or (_42436_, _42435_, _22731_);
  and (_42437_, _42436_, _42434_);
  or (_42438_, _42437_, _42430_);
  or (_42439_, _15686_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_42440_, _42439_, _39026_);
  and (_12329_, _42440_, _42438_);
  and (_42441_, _42375_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_42442_, _22159_, _21274_);
  and (_42443_, _21448_, _20685_);
  and (_42444_, _21230_, _21143_);
  or (_42445_, _42444_, _42406_);
  or (_42446_, _42445_, _42443_);
  or (_42447_, _42446_, _42442_);
  or (_42448_, _42393_, _22489_);
  or (_42449_, _20729_, _20347_);
  and (_42450_, _42449_, _39612_);
  or (_42451_, _22126_, _21732_);
  and (_42452_, _42451_, _19617_);
  or (_42453_, _42452_, _42450_);
  or (_42454_, _42453_, _42448_);
  or (_42455_, _42454_, _42447_);
  and (_42456_, _42455_, _41166_);
  or (_12332_, _42456_, _42441_);
  and (_42457_, _42375_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_42458_, _22742_, _22038_);
  and (_42459_, _22038_, _21230_);
  or (_42460_, _42459_, _22203_);
  or (_42461_, _42460_, _42458_);
  not (_42462_, _39627_);
  and (_42463_, _20805_, _21372_);
  or (_42464_, _42463_, _21470_);
  and (_42465_, _21143_, _19617_);
  or (_42466_, _42465_, _42464_);
  or (_42467_, _42466_, _42462_);
  or (_42468_, _42467_, _42461_);
  and (_42469_, _22368_, _20805_);
  and (_42470_, _39615_, _19857_);
  or (_42471_, _42470_, _42469_);
  and (_42472_, _21241_, _20337_);
  and (_42473_, _21776_, _22280_);
  or (_42474_, _42473_, _42472_);
  or (_42475_, _42474_, _42471_);
  nor (_42476_, _42392_, _22214_);
  nand (_42477_, _42476_, _22060_);
  or (_42478_, _42477_, _42475_);
  or (_42479_, _42478_, _42410_);
  or (_42480_, _42479_, _42468_);
  and (_42481_, _42480_, _41166_);
  or (_12335_, _42481_, _42457_);
  and (_42482_, _39612_, _20751_);
  and (_42483_, _21776_, _20838_);
  or (_42484_, _42483_, _42482_);
  or (_42485_, _42484_, _20849_);
  and (_42486_, _20838_, _19067_);
  or (_42487_, _42486_, _20773_);
  or (_42488_, _42487_, _42485_);
  and (_42489_, _21776_, _20762_);
  or (_42490_, _42489_, _42400_);
  or (_42491_, _42490_, _42488_);
  and (_42492_, _42491_, _41166_);
  and (_42493_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_42494_, _42493_, _22786_);
  and (_42495_, _42494_, _39026_);
  or (_12337_, _42495_, _42492_);
  and (_42496_, _21307_, _20620_);
  and (_42497_, _42496_, _19617_);
  or (_42498_, _42497_, _20358_);
  or (_42499_, _42498_, _21983_);
  not (_42500_, _22148_);
  and (_42501_, _42496_, _21786_);
  or (_42502_, _42501_, _42500_);
  or (_42503_, _42502_, _42408_);
  nor (_42504_, _42431_, _22170_);
  nand (_42505_, _42504_, _22467_);
  nor (_42506_, _22489_, _22335_);
  nand (_42507_, _42506_, _22093_);
  or (_42508_, _42507_, _42505_);
  nor (_42509_, _42508_, _42503_);
  nand (_42510_, _42509_, _22324_);
  and (_42511_, _39612_, _21307_);
  or (_42512_, _42511_, _21885_);
  and (_42513_, _20751_, _21372_);
  or (_42514_, _42432_, _42513_);
  and (_42515_, _22368_, _20751_);
  or (_42516_, _42515_, _22379_);
  or (_42517_, _42516_, _42514_);
  or (_42518_, _42517_, _42512_);
  or (_42519_, _42394_, _39625_);
  or (_42520_, _42519_, _42518_);
  or (_42521_, _42520_, _42510_);
  or (_42522_, _42521_, _42499_);
  and (_42523_, _42522_, _18653_);
  and (_42524_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42525_, _42435_, _42401_);
  and (_42526_, _21743_, _21557_);
  or (_42527_, _42526_, _42525_);
  or (_42528_, _42527_, _42524_);
  or (_42529_, _42528_, _42523_);
  and (_12340_, _42529_, _39026_);
  nor (_12382_, _21623_, rst);
  nor (_12384_, _22676_, rst);
  nand (_12387_, _42428_, _41166_);
  nand (_42530_, _42424_, _41166_);
  not (_42531_, _21132_);
  or (_42532_, _42336_, _42531_);
  and (_12389_, _42532_, _42530_);
  or (_42533_, _42338_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_42534_, _42533_, _42341_);
  or (_42535_, _42534_, _42352_);
  and (_42536_, _42535_, _42369_);
  nor (_42537_, _42368_, _21536_);
  or (_42538_, _42537_, rst);
  or (_12392_, _42538_, _42536_);
  nand (_42539_, _21089_, _18598_);
  or (_42540_, _18598_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_42541_, _42540_, _39026_);
  and (_12395_, _42541_, _42539_);
  not (_42542_, _18598_);
  or (_42543_, _19584_, _42542_);
  or (_42544_, _18598_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_42545_, _42544_, _39026_);
  and (_12397_, _42545_, _42543_);
  nand (_42546_, _19286_, _18598_);
  or (_42547_, _18598_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_42548_, _42547_, _39026_);
  and (_12400_, _42548_, _42546_);
  nand (_42549_, _19046_, _18598_);
  or (_42550_, _18598_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_42551_, _42550_, _39026_);
  and (_12403_, _42551_, _42549_);
  or (_42552_, _20598_, _42542_);
  or (_42553_, _18598_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_42554_, _42553_, _39026_);
  and (_12405_, _42554_, _42552_);
  nand (_42555_, _19835_, _18598_);
  or (_42556_, _18598_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_42557_, _42556_, _39026_);
  and (_12408_, _42557_, _42555_);
  nand (_42558_, _20075_, _18598_);
  or (_42559_, _18598_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_42560_, _42559_, _39026_);
  and (_12411_, _42560_, _42558_);
  or (_42561_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _15686_);
  and (_42562_, _42561_, _42430_);
  and (_42563_, _22742_, _20620_);
  and (_42564_, _42563_, _42449_);
  or (_42565_, _42564_, _42407_);
  and (_42566_, _22038_, _21776_);
  or (_42567_, _42566_, _42390_);
  or (_42568_, _42486_, _39613_);
  or (_42569_, _42568_, _42567_);
  or (_42570_, _42569_, _42565_);
  and (_42571_, _22280_, _19617_);
  or (_42572_, _42571_, _21274_);
  or (_42573_, _21808_, _21416_);
  or (_42574_, _42573_, _42572_);
  or (_42575_, _42470_, _20773_);
  or (_42576_, _42575_, _42489_);
  or (_42577_, _42576_, _42485_);
  or (_42578_, _42577_, _42574_);
  and (_42579_, _22368_, _21405_);
  and (_42580_, _42496_, _22742_);
  or (_42581_, _42580_, _42472_);
  or (_42582_, _42581_, _42579_);
  and (_42583_, _21874_, _19617_);
  or (_42584_, _39619_, _42583_);
  or (_42585_, _42473_, _42381_);
  or (_42586_, _42585_, _42584_);
  or (_42587_, _42586_, _42582_);
  or (_42588_, _42587_, _42578_);
  or (_42589_, _42588_, _42570_);
  and (_42590_, _42589_, _18653_);
  or (_42591_, _42590_, _42562_);
  and (_37213_, _42591_, _39026_);
  and (_42592_, _42375_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_42593_, _42567_, _42466_);
  and (_42594_, _22742_, _22280_);
  or (_42595_, _20816_, _20685_);
  and (_42596_, _42595_, _42563_);
  or (_42597_, _42596_, _42594_);
  or (_42598_, _42597_, _42383_);
  or (_42599_, _42598_, _42593_);
  not (_42600_, _22082_);
  nand (_42601_, _22500_, _42600_);
  nor (_42602_, _42471_, _22302_);
  nand (_42603_, _42602_, _40522_);
  or (_42604_, _42603_, _42601_);
  and (_42605_, _22742_, _20838_);
  or (_42606_, _42605_, _42413_);
  or (_42607_, _42606_, _42604_);
  or (_42608_, _42607_, _42599_);
  and (_42609_, _42608_, _41166_);
  or (_37214_, _42609_, _42592_);
  or (_42610_, _42515_, _21885_);
  or (_42611_, _42610_, _42514_);
  or (_42612_, _42611_, _42510_);
  and (_42613_, _42612_, _18653_);
  and (_42614_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_42615_, _42614_, _42527_);
  or (_42616_, _42615_, _42613_);
  and (_37215_, _42616_, _39026_);
  and (_42617_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_42618_, _22258_, _20631_);
  or (_42619_, _42618_, _20740_);
  or (_42620_, _42619_, _42499_);
  or (_42621_, _42620_, _42433_);
  and (_42622_, _42621_, _18653_);
  or (_42623_, _42622_, _42617_);
  or (_42624_, _42623_, _42525_);
  and (_37216_, _42624_, _39026_);
  and (_42625_, _22742_, _22126_);
  or (_42626_, _42489_, _42625_);
  and (_42627_, _42563_, _21383_);
  or (_42628_, _42627_, _42565_);
  or (_42629_, _42381_, _40517_);
  or (_42630_, _42629_, _22753_);
  or (_42631_, _42630_, _42628_);
  or (_42632_, _42631_, _42626_);
  or (_42633_, _42482_, _20860_);
  or (_42634_, _42568_, _42472_);
  or (_42635_, _39619_, _22764_);
  and (_42636_, _21776_, _21710_);
  or (_42637_, _42636_, _42424_);
  or (_42638_, _42637_, _42635_);
  or (_42639_, _42638_, _42634_);
  or (_42640_, _42639_, _42633_);
  and (_42641_, _42501_, _20326_);
  or (_42642_, _42497_, _20773_);
  or (_42643_, _42642_, _42511_);
  or (_42644_, _42458_, _21339_);
  or (_42645_, _42644_, _42643_);
  or (_42646_, _42645_, _42641_);
  and (_42647_, _21448_, _21874_);
  or (_42648_, _42594_, _42647_);
  and (_42649_, _22742_, _21329_);
  and (_42650_, _42483_, _20631_);
  or (_42651_, _42650_, _42649_);
  or (_42652_, _42651_, _42648_);
  or (_42653_, _42652_, _42433_);
  or (_42654_, _42653_, _42646_);
  or (_42655_, _42654_, _42640_);
  or (_42656_, _42655_, _42632_);
  and (_42657_, _42656_, _18653_);
  and (_42658_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_42659_, _42429_, _22786_);
  or (_42660_, _42659_, _42658_);
  or (_42661_, _42660_, _42657_);
  and (_37217_, _42661_, _39026_);
  or (_42662_, _42390_, _20773_);
  nor (_42663_, _42662_, _21885_);
  nand (_42664_, _42663_, _21350_);
  or (_42665_, _22038_, _22280_);
  and (_42666_, _42665_, _21241_);
  or (_42667_, _42666_, _21939_);
  or (_42668_, _42667_, _42664_);
  or (_42669_, _42501_, _22764_);
  and (_42670_, _42511_, _20326_);
  and (_42671_, _42497_, _20326_);
  or (_42672_, _42671_, _42670_);
  or (_42673_, _42672_, _42669_);
  or (_42674_, _42673_, _42634_);
  or (_42675_, _42674_, _42633_);
  or (_42676_, _42675_, _42668_);
  or (_42677_, _42676_, _42632_);
  and (_42678_, _42677_, _18653_);
  and (_42679_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_42680_, _42679_, _42659_);
  or (_42681_, _42680_, _42678_);
  and (_37218_, _42681_, _39026_);
  and (_42682_, _42375_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_42683_, _42406_, _21111_);
  or (_42684_, _42564_, _42683_);
  and (_42685_, _42392_, _21111_);
  or (_42686_, _42685_, _22335_);
  and (_42687_, _21732_, _21241_);
  or (_42688_, _42687_, _42377_);
  or (_00010_, _42688_, _42686_);
  or (_00011_, _00010_, _42684_);
  and (_00012_, _21710_, _20871_);
  or (_00013_, _42489_, _20773_);
  nor (_00014_, _00013_, _00012_);
  nand (_00015_, _00014_, _37347_);
  not (_00016_, _37346_);
  or (_00017_, _42442_, _00016_);
  or (_00018_, _00017_, _00015_);
  and (_00019_, _21710_, _21241_);
  or (_00020_, _00019_, _22445_);
  and (_00021_, _21241_, _21819_);
  or (_00022_, _42482_, _42393_);
  or (_00023_, _00022_, _00021_);
  or (_00024_, _00023_, _00020_);
  or (_00025_, _00024_, _42453_);
  or (_00026_, _00025_, _00018_);
  or (_00027_, _00026_, _00011_);
  and (_00028_, _00027_, _41166_);
  or (_37219_, _00028_, _42682_);
  and (_00029_, _42563_, _20729_);
  or (_00030_, _00029_, _00019_);
  or (_00031_, _42638_, _42461_);
  or (_00032_, _00031_, _00030_);
  or (_00033_, _21906_, _20860_);
  or (_00034_, _42568_, _42687_);
  or (_00035_, _00034_, _00033_);
  or (_00036_, _42463_, _42392_);
  or (_00037_, _42650_, _42465_);
  or (_00038_, _00037_, _00036_);
  or (_00039_, _22049_, _21339_);
  or (_00040_, _42469_, _21274_);
  or (_00041_, _00040_, _00039_);
  or (_00042_, _00041_, _00038_);
  or (_00043_, _00042_, _00035_);
  or (_00044_, _00043_, _00032_);
  and (_00045_, _00044_, _41166_);
  and (_00046_, _42375_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_00047_, _18609_, _39026_);
  and (_00049_, _00047_, _22764_);
  or (_00051_, _00049_, _00046_);
  or (_37220_, _00051_, _00045_);
  and (_00054_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00056_, _22764_, _15686_);
  or (_00058_, _00056_, _00054_);
  and (_00060_, _00058_, _39026_);
  or (_00061_, _39614_, _20794_);
  or (_00062_, _00061_, _42629_);
  or (_00063_, _00021_, _42627_);
  or (_00064_, _00063_, _22115_);
  or (_00065_, _42489_, _22027_);
  or (_00066_, _00065_, _42392_);
  and (_00068_, _21241_, _20838_);
  or (_00069_, _00068_, _00022_);
  nor (_00071_, _00069_, _00066_);
  nand (_00072_, _00071_, _39620_);
  or (_00073_, _00072_, _00064_);
  or (_00074_, _00073_, _00062_);
  or (_00075_, _00074_, _42412_);
  and (_00076_, _00075_, _41166_);
  or (_37221_, _00076_, _00060_);
  or (_00077_, _22753_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00078_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15686_);
  and (_00079_, _00078_, _39026_);
  and (_00080_, _00079_, _00077_);
  or (_00081_, _42684_, _42448_);
  or (_00082_, _00081_, _00064_);
  or (_00083_, _39614_, _21906_);
  or (_00084_, _00083_, _39625_);
  or (_00085_, _20740_, _20358_);
  or (_00086_, _00085_, _22214_);
  and (_00087_, _21241_, _20347_);
  or (_00088_, _00087_, _39619_);
  or (_00089_, _00088_, _00086_);
  or (_00090_, _00089_, _42409_);
  or (_00091_, _00090_, _00084_);
  or (_00092_, _00091_, _00082_);
  and (_00093_, _00092_, _41166_);
  or (_37222_, _00093_, _00080_);
  and (_00094_, _42375_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_00095_, _42384_, _00016_);
  or (_00096_, _42688_, _41448_);
  or (_00097_, _00096_, _42489_);
  and (_00099_, _00068_, _20620_);
  or (_00101_, _00029_, _00099_);
  or (_00103_, _00101_, _00021_);
  nor (_00105_, _40517_, _22346_);
  nand (_00107_, _00105_, _37347_);
  or (_00109_, _00107_, _00103_);
  or (_00111_, _00109_, _00097_);
  or (_00112_, _00111_, _00095_);
  or (_00113_, _00112_, _42488_);
  and (_00114_, _00113_, _41166_);
  or (_37224_, _00114_, _00094_);
  not (_00115_, _39364_);
  nor (_00116_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00118_, _42287_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00119_, _00118_, _00116_);
  nor (_00121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00122_, _42291_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00123_, _00122_, _00121_);
  nor (_00124_, _00123_, _00119_);
  nor (_00125_, _41493_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00126_, _42295_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00127_, _00126_, _00125_);
  and (_00128_, _00127_, _00124_);
  nor (_00129_, _41512_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00130_, _42299_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00131_, _00130_, _00129_);
  and (_00132_, _00131_, _00128_);
  and (_00133_, _00132_, _00115_);
  not (_00134_, _39323_);
  and (_00135_, _00123_, _00119_);
  not (_00136_, _00124_);
  nor (_00137_, _00127_, _00136_);
  and (_00138_, _00127_, _00136_);
  nor (_00139_, _00138_, _00137_);
  and (_00140_, _00131_, _00139_);
  and (_00141_, _00140_, _00135_);
  and (_00142_, _00141_, _00134_);
  not (_00143_, _39282_);
  not (_00144_, _00123_);
  nor (_00145_, _00144_, _00119_);
  and (_00146_, _00140_, _00145_);
  and (_00147_, _00146_, _00143_);
  or (_00148_, _00147_, _00142_);
  not (_00149_, _39200_);
  and (_00151_, _00131_, _00137_);
  and (_00153_, _00151_, _00149_);
  not (_00155_, _39241_);
  and (_00157_, _00144_, _00119_);
  and (_00159_, _00140_, _00157_);
  and (_00161_, _00159_, _00155_);
  or (_00163_, _00161_, _00153_);
  or (_00164_, _00163_, _00148_);
  not (_00165_, _39159_);
  not (_00166_, _00139_);
  nor (_00167_, _00131_, _00138_);
  and (_00168_, _00131_, _00138_);
  nor (_00169_, _00168_, _00167_);
  and (_00171_, _00169_, _00166_);
  and (_00172_, _00171_, _00135_);
  and (_00174_, _00172_, _00165_);
  not (_00175_, _39118_);
  and (_00176_, _00171_, _00145_);
  and (_00177_, _00176_, _00175_);
  or (_00178_, _00177_, _00174_);
  not (_00179_, _39077_);
  and (_00180_, _00157_, _00171_);
  and (_00181_, _00180_, _00179_);
  not (_00182_, _39036_);
  and (_00183_, _00167_, _00128_);
  and (_00184_, _00183_, _00182_);
  or (_00185_, _00184_, _00181_);
  or (_00186_, _00185_, _00178_);
  or (_00187_, _00186_, _00164_);
  not (_00188_, _38982_);
  and (_00189_, _00167_, _00135_);
  and (_00190_, _00189_, _00188_);
  not (_00191_, _38940_);
  and (_00192_, _00167_, _00145_);
  and (_00193_, _00192_, _00191_);
  or (_00194_, _00193_, _00190_);
  not (_00195_, _38857_);
  nor (_00196_, _00169_, _00139_);
  and (_00197_, _00196_, _00124_);
  and (_00198_, _00197_, _00195_);
  not (_00199_, _38898_);
  and (_00200_, _00157_, _00167_);
  and (_00201_, _00200_, _00199_);
  or (_00202_, _00201_, _00198_);
  or (_00204_, _00202_, _00194_);
  not (_00206_, _38580_);
  and (_00208_, _00157_, _00196_);
  and (_00210_, _00208_, _00206_);
  not (_00212_, _38659_);
  and (_00214_, _00196_, _00145_);
  and (_00216_, _00214_, _00212_);
  not (_00217_, _38793_);
  and (_00218_, _00196_, _00135_);
  and (_00219_, _00218_, _00217_);
  or (_00220_, _00219_, _00216_);
  or (_00221_, _00220_, _00210_);
  or (_00222_, _00221_, _00204_);
  or (_00224_, _00222_, _00187_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _00224_, _00133_);
  and (_00226_, _00208_, _00115_);
  and (_00227_, _00141_, _00143_);
  and (_00228_, _00146_, _00155_);
  and (_00229_, _00159_, _00149_);
  or (_00230_, _00229_, _00228_);
  or (_00231_, _00230_, _00227_);
  or (_00232_, _00231_, _00226_);
  and (_00233_, _00214_, _00206_);
  and (_00234_, _00197_, _00217_);
  or (_00235_, _00234_, _00233_);
  or (_00236_, _00235_, _00232_);
  and (_00237_, _00132_, _00134_);
  and (_00238_, _00151_, _00165_);
  and (_00239_, _00172_, _00175_);
  or (_00240_, _00239_, _00238_);
  and (_00241_, _00180_, _00182_);
  and (_00242_, _00176_, _00179_);
  or (_00243_, _00242_, _00241_);
  or (_00244_, _00243_, _00240_);
  and (_00245_, _00200_, _00195_);
  and (_00246_, _00183_, _00188_);
  and (_00247_, _00189_, _00191_);
  or (_00248_, _00247_, _00246_);
  or (_00249_, _00248_, _00245_);
  and (_00250_, _00218_, _00212_);
  and (_00251_, _00192_, _00199_);
  or (_00252_, _00251_, _00250_);
  or (_00253_, _00252_, _00249_);
  or (_00254_, _00253_, _00244_);
  or (_00256_, _00254_, _00237_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _00256_, _00236_);
  and (_00259_, _00214_, _00115_);
  and (_00261_, _00159_, _00165_);
  and (_00263_, _00151_, _00175_);
  or (_00265_, _00263_, _00261_);
  and (_00267_, _00172_, _00179_);
  and (_00268_, _00176_, _00182_);
  or (_00269_, _00268_, _00267_);
  or (_00270_, _00269_, _00265_);
  and (_00271_, _00141_, _00155_);
  and (_00272_, _00146_, _00149_);
  or (_00273_, _00272_, _00271_);
  and (_00275_, _00132_, _00143_);
  and (_00276_, _00208_, _00134_);
  or (_00278_, _00276_, _00275_);
  or (_00279_, _00278_, _00273_);
  or (_00280_, _00279_, _00270_);
  and (_00281_, _00218_, _00206_);
  and (_00282_, _00197_, _00212_);
  and (_00283_, _00200_, _00217_);
  or (_00284_, _00283_, _00282_);
  or (_00285_, _00284_, _00281_);
  and (_00286_, _00192_, _00195_);
  and (_00287_, _00189_, _00199_);
  or (_00288_, _00287_, _00286_);
  and (_00289_, _00180_, _00188_);
  and (_00290_, _00183_, _00191_);
  or (_00291_, _00290_, _00289_);
  or (_00292_, _00291_, _00288_);
  or (_00293_, _00292_, _00285_);
  or (_00294_, _00293_, _00280_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _00294_, _00259_);
  and (_00295_, _00218_, _00115_);
  and (_00296_, _00180_, _00191_);
  and (_00297_, _00183_, _00199_);
  and (_00298_, _00189_, _00195_);
  or (_00299_, _00298_, _00297_);
  or (_00300_, _00299_, _00296_);
  and (_00301_, _00176_, _00188_);
  and (_00302_, _00197_, _00206_);
  and (_00303_, _00192_, _00217_);
  and (_00304_, _00200_, _00212_);
  or (_00305_, _00304_, _00303_);
  or (_00307_, _00305_, _00302_);
  or (_00309_, _00307_, _00301_);
  or (_00311_, _00309_, _00300_);
  and (_00313_, _00172_, _00182_);
  and (_00315_, _00151_, _00179_);
  and (_00317_, _00146_, _00165_);
  and (_00319_, _00159_, _00175_);
  or (_00320_, _00319_, _00317_);
  or (_00321_, _00320_, _00315_);
  or (_00322_, _00321_, _00313_);
  and (_00323_, _00214_, _00134_);
  and (_00324_, _00208_, _00143_);
  or (_00325_, _00324_, _00323_);
  and (_00327_, _00132_, _00155_);
  and (_00328_, _00141_, _00149_);
  or (_00330_, _00328_, _00327_);
  or (_00331_, _00330_, _00325_);
  or (_00332_, _00331_, _00322_);
  or (_00333_, _00332_, _00311_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _00333_, _00295_);
  not (_00334_, _39369_);
  and (_00335_, _00218_, _00334_);
  not (_00336_, _38945_);
  and (_00337_, _00180_, _00336_);
  not (_00338_, _38903_);
  and (_00339_, _00183_, _00338_);
  not (_00340_, _38862_);
  and (_00341_, _00189_, _00340_);
  or (_00342_, _00341_, _00339_);
  or (_00343_, _00342_, _00337_);
  not (_00344_, _38987_);
  and (_00345_, _00176_, _00344_);
  not (_00346_, _38612_);
  and (_00347_, _00197_, _00346_);
  not (_00348_, _38807_);
  and (_00349_, _00192_, _00348_);
  not (_00350_, _38677_);
  and (_00351_, _00200_, _00350_);
  or (_00352_, _00351_, _00349_);
  or (_00353_, _00352_, _00347_);
  or (_00354_, _00353_, _00345_);
  or (_00355_, _00354_, _00343_);
  not (_00356_, _39041_);
  and (_00357_, _00172_, _00356_);
  not (_00359_, _39164_);
  and (_00361_, _00146_, _00359_);
  not (_00363_, _39123_);
  and (_00365_, _00159_, _00363_);
  or (_00367_, _00365_, _00361_);
  not (_00369_, _39082_);
  and (_00371_, _00151_, _00369_);
  or (_00372_, _00371_, _00367_);
  or (_00373_, _00372_, _00357_);
  not (_00374_, _39287_);
  and (_00375_, _00208_, _00374_);
  not (_00376_, _39328_);
  and (_00377_, _00214_, _00376_);
  or (_00379_, _00377_, _00375_);
  not (_00380_, _39205_);
  and (_00382_, _00141_, _00380_);
  not (_00383_, _39246_);
  and (_00384_, _00132_, _00383_);
  or (_00385_, _00384_, _00382_);
  or (_00386_, _00385_, _00379_);
  or (_00387_, _00386_, _00373_);
  or (_00388_, _00387_, _00355_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _00388_, _00335_);
  not (_00389_, _38950_);
  and (_00390_, _00180_, _00389_);
  not (_00391_, _38867_);
  and (_00392_, _00189_, _00391_);
  not (_00393_, _38908_);
  and (_00394_, _00183_, _00393_);
  or (_00395_, _00394_, _00392_);
  or (_00396_, _00395_, _00390_);
  not (_00397_, _39210_);
  and (_00398_, _00141_, _00397_);
  not (_00399_, _39333_);
  and (_00400_, _00214_, _00399_);
  not (_00401_, _39374_);
  and (_00402_, _00218_, _00401_);
  or (_00403_, _00402_, _00400_);
  or (_00404_, _00403_, _00398_);
  or (_00405_, _00404_, _00396_);
  not (_00406_, _39251_);
  and (_00407_, _00132_, _00406_);
  not (_00408_, _39087_);
  and (_00409_, _00151_, _00408_);
  not (_00411_, _39128_);
  and (_00413_, _00159_, _00411_);
  not (_00415_, _39169_);
  and (_00417_, _00146_, _00415_);
  or (_00419_, _00417_, _00413_);
  or (_00421_, _00419_, _00409_);
  not (_00423_, _39046_);
  and (_00424_, _00172_, _00423_);
  not (_00425_, _39292_);
  and (_00426_, _00208_, _00425_);
  or (_00427_, _00426_, _00424_);
  or (_00428_, _00427_, _00421_);
  not (_00429_, _38992_);
  and (_00431_, _00176_, _00429_);
  not (_00432_, _38617_);
  and (_00434_, _00197_, _00432_);
  not (_00435_, _38826_);
  and (_00436_, _00192_, _00435_);
  not (_00437_, _38690_);
  and (_00438_, _00200_, _00437_);
  or (_00439_, _00438_, _00436_);
  or (_00440_, _00439_, _00434_);
  or (_00441_, _00440_, _00431_);
  or (_00442_, _00441_, _00428_);
  or (_00443_, _00442_, _00407_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _00443_, _00405_);
  not (_00444_, _38955_);
  and (_00445_, _00180_, _00444_);
  not (_00446_, _38913_);
  and (_00447_, _00183_, _00446_);
  not (_00448_, _38872_);
  and (_00449_, _00189_, _00448_);
  or (_00450_, _00449_, _00447_);
  or (_00451_, _00450_, _00445_);
  not (_00452_, _39297_);
  and (_00453_, _00208_, _00452_);
  not (_00454_, _39338_);
  and (_00455_, _00214_, _00454_);
  not (_00456_, _39379_);
  and (_00457_, _00218_, _00456_);
  or (_00458_, _00457_, _00455_);
  or (_00459_, _00458_, _00453_);
  or (_00460_, _00459_, _00451_);
  not (_00461_, _39256_);
  and (_00463_, _00132_, _00461_);
  not (_00465_, _39051_);
  and (_00467_, _00172_, _00465_);
  not (_00469_, _39133_);
  and (_00471_, _00159_, _00469_);
  not (_00473_, _39174_);
  and (_00475_, _00146_, _00473_);
  or (_00476_, _00475_, _00471_);
  or (_00477_, _00476_, _00467_);
  not (_00478_, _39092_);
  and (_00479_, _00151_, _00478_);
  not (_00480_, _39215_);
  and (_00481_, _00141_, _00480_);
  or (_00483_, _00481_, _00479_);
  or (_00484_, _00483_, _00477_);
  not (_00486_, _39000_);
  and (_00487_, _00176_, _00486_);
  not (_00488_, _38622_);
  and (_00489_, _00197_, _00488_);
  not (_00490_, _38831_);
  and (_00491_, _00192_, _00490_);
  not (_00492_, _38707_);
  and (_00493_, _00200_, _00492_);
  or (_00494_, _00493_, _00491_);
  or (_00495_, _00494_, _00489_);
  or (_00496_, _00495_, _00487_);
  or (_00497_, _00496_, _00484_);
  or (_00498_, _00497_, _00463_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _00498_, _00460_);
  not (_00499_, _39384_);
  and (_00500_, _00218_, _00499_);
  not (_00501_, _38960_);
  and (_00502_, _00180_, _00501_);
  not (_00503_, _38918_);
  and (_00504_, _00183_, _00503_);
  not (_00505_, _38877_);
  and (_00506_, _00189_, _00505_);
  or (_00507_, _00506_, _00504_);
  or (_00508_, _00507_, _00502_);
  not (_00509_, _39005_);
  and (_00510_, _00176_, _00509_);
  not (_00511_, _38627_);
  and (_00512_, _00197_, _00511_);
  not (_00513_, _38836_);
  and (_00515_, _00192_, _00513_);
  not (_00517_, _38724_);
  and (_00519_, _00200_, _00517_);
  or (_00521_, _00519_, _00515_);
  or (_00523_, _00521_, _00512_);
  or (_00525_, _00523_, _00510_);
  or (_00527_, _00525_, _00508_);
  not (_00528_, _39056_);
  and (_00529_, _00172_, _00528_);
  not (_00530_, _39097_);
  and (_00531_, _00151_, _00530_);
  not (_00532_, _39179_);
  and (_00533_, _00146_, _00532_);
  not (_00535_, _39138_);
  and (_00536_, _00159_, _00535_);
  or (_00538_, _00536_, _00533_);
  or (_00539_, _00538_, _00531_);
  or (_00540_, _00539_, _00529_);
  not (_00541_, _39343_);
  and (_00542_, _00214_, _00541_);
  not (_00543_, _39302_);
  and (_00544_, _00208_, _00543_);
  or (_00545_, _00544_, _00542_);
  not (_00546_, _39261_);
  and (_00547_, _00132_, _00546_);
  not (_00548_, _39220_);
  and (_00549_, _00141_, _00548_);
  or (_00550_, _00549_, _00547_);
  or (_00551_, _00550_, _00545_);
  or (_00552_, _00551_, _00540_);
  or (_00553_, _00552_, _00527_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _00553_, _00500_);
  not (_00554_, _38965_);
  and (_00555_, _00180_, _00554_);
  not (_00556_, _38882_);
  and (_00557_, _00189_, _00556_);
  not (_00558_, _38923_);
  and (_00559_, _00183_, _00558_);
  or (_00560_, _00559_, _00557_);
  or (_00561_, _00560_, _00555_);
  not (_00562_, _39307_);
  and (_00563_, _00208_, _00562_);
  not (_00564_, _39348_);
  and (_00565_, _00214_, _00564_);
  not (_00567_, _39389_);
  and (_00569_, _00218_, _00567_);
  or (_00571_, _00569_, _00565_);
  or (_00573_, _00571_, _00563_);
  or (_00575_, _00573_, _00561_);
  not (_00577_, _39266_);
  and (_00579_, _00132_, _00577_);
  not (_00580_, _39061_);
  and (_00581_, _00172_, _00580_);
  not (_00582_, _39184_);
  and (_00583_, _00146_, _00582_);
  not (_00584_, _39143_);
  and (_00585_, _00159_, _00584_);
  or (_00587_, _00585_, _00583_);
  or (_00588_, _00587_, _00581_);
  not (_00590_, _39225_);
  and (_00591_, _00141_, _00590_);
  not (_00592_, _39102_);
  and (_00593_, _00151_, _00592_);
  or (_00594_, _00593_, _00591_);
  or (_00595_, _00594_, _00588_);
  not (_00596_, _39010_);
  and (_00597_, _00176_, _00596_);
  not (_00598_, _38632_);
  and (_00599_, _00197_, _00598_);
  not (_00600_, _38841_);
  and (_00601_, _00192_, _00600_);
  not (_00602_, _38737_);
  and (_00603_, _00200_, _00602_);
  or (_00604_, _00603_, _00601_);
  or (_00605_, _00604_, _00599_);
  or (_00606_, _00605_, _00597_);
  or (_00607_, _00606_, _00595_);
  or (_00608_, _00607_, _00579_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _00608_, _00575_);
  not (_00609_, _38970_);
  and (_00610_, _00180_, _00609_);
  not (_00611_, _38928_);
  and (_00612_, _00183_, _00611_);
  not (_00613_, _38887_);
  and (_00614_, _00189_, _00613_);
  or (_00615_, _00614_, _00612_);
  or (_00616_, _00615_, _00610_);
  not (_00617_, _39230_);
  and (_00619_, _00141_, _00617_);
  not (_00621_, _39394_);
  and (_00623_, _00218_, _00621_);
  not (_00625_, _39353_);
  and (_00627_, _00214_, _00625_);
  or (_00629_, _00627_, _00623_);
  or (_00631_, _00629_, _00619_);
  or (_00632_, _00631_, _00616_);
  not (_00633_, _39271_);
  and (_00634_, _00132_, _00633_);
  not (_00635_, _39066_);
  and (_00636_, _00172_, _00635_);
  not (_00637_, _39189_);
  and (_00639_, _00146_, _00637_);
  not (_00640_, _39148_);
  and (_00642_, _00159_, _00640_);
  or (_00643_, _00642_, _00639_);
  or (_00644_, _00643_, _00636_);
  not (_00645_, _39107_);
  and (_00646_, _00151_, _00645_);
  not (_00647_, _39312_);
  and (_00648_, _00208_, _00647_);
  or (_00649_, _00648_, _00646_);
  or (_00650_, _00649_, _00644_);
  not (_00651_, _39015_);
  and (_00652_, _00176_, _00651_);
  not (_00653_, _38637_);
  and (_00654_, _00197_, _00653_);
  not (_00655_, _38846_);
  and (_00656_, _00192_, _00655_);
  not (_00657_, _38758_);
  and (_00658_, _00200_, _00657_);
  or (_00659_, _00658_, _00656_);
  or (_00660_, _00659_, _00654_);
  or (_00661_, _00660_, _00652_);
  or (_00662_, _00661_, _00650_);
  or (_00663_, _00662_, _00634_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _00663_, _00632_);
  not (_00664_, _39399_);
  and (_00665_, _00218_, _00664_);
  not (_00666_, _38976_);
  and (_00667_, _00180_, _00666_);
  not (_00668_, _38933_);
  and (_00669_, _00183_, _00668_);
  not (_00671_, _38892_);
  and (_00673_, _00189_, _00671_);
  or (_00675_, _00673_, _00669_);
  or (_00677_, _00675_, _00667_);
  not (_00679_, _39025_);
  and (_00681_, _00176_, _00679_);
  not (_00683_, _38642_);
  and (_00684_, _00197_, _00683_);
  not (_00685_, _38851_);
  and (_00686_, _00192_, _00685_);
  not (_00687_, _38771_);
  and (_00688_, _00200_, _00687_);
  or (_00689_, _00688_, _00686_);
  or (_00691_, _00689_, _00684_);
  or (_00692_, _00691_, _00681_);
  or (_00694_, _00692_, _00677_);
  not (_00695_, _39112_);
  and (_00696_, _00151_, _00695_);
  not (_00697_, _39194_);
  and (_00698_, _00146_, _00697_);
  not (_00699_, _39153_);
  and (_00700_, _00159_, _00699_);
  or (_00701_, _00700_, _00698_);
  not (_00702_, _39071_);
  and (_00703_, _00172_, _00702_);
  or (_00704_, _00703_, _00701_);
  or (_00705_, _00704_, _00696_);
  not (_00706_, _39317_);
  and (_00707_, _00208_, _00706_);
  not (_00708_, _39358_);
  and (_00709_, _00214_, _00708_);
  or (_00710_, _00709_, _00707_);
  not (_00711_, _39235_);
  and (_00712_, _00141_, _00711_);
  not (_00713_, _39276_);
  and (_00714_, _00132_, _00713_);
  or (_00715_, _00714_, _00712_);
  or (_00716_, _00715_, _00710_);
  or (_00717_, _00716_, _00705_);
  or (_00718_, _00717_, _00694_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _00718_, _00665_);
  and (_00719_, _00200_, _00348_);
  and (_00720_, _00218_, _00346_);
  or (_00721_, _00720_, _00719_);
  and (_00723_, _00172_, _00369_);
  and (_00725_, _00159_, _00359_);
  and (_00727_, _00151_, _00363_);
  or (_00729_, _00727_, _00725_);
  or (_00731_, _00729_, _00723_);
  or (_00733_, _00731_, _00721_);
  and (_00735_, _00132_, _00374_);
  and (_00736_, _00141_, _00383_);
  and (_00737_, _00146_, _00380_);
  or (_00738_, _00737_, _00736_);
  and (_00739_, _00208_, _00376_);
  or (_00740_, _00739_, _00738_);
  and (_00741_, _00176_, _00356_);
  and (_00743_, _00214_, _00334_);
  or (_00744_, _00743_, _00741_);
  or (_00746_, _00744_, _00740_);
  and (_00747_, _00183_, _00336_);
  and (_00748_, _00189_, _00338_);
  and (_00749_, _00192_, _00340_);
  or (_00750_, _00749_, _00748_);
  or (_00751_, _00750_, _00747_);
  and (_00752_, _00180_, _00344_);
  and (_00753_, _00197_, _00350_);
  or (_00754_, _00753_, _00752_);
  or (_00755_, _00754_, _00751_);
  or (_00756_, _00755_, _00746_);
  or (_00757_, _00756_, _00735_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _00757_, _00733_);
  and (_00758_, _00214_, _00401_);
  and (_00759_, _00146_, _00397_);
  and (_00760_, _00141_, _00406_);
  or (_00761_, _00760_, _00759_);
  and (_00762_, _00132_, _00425_);
  and (_00763_, _00208_, _00399_);
  or (_00764_, _00763_, _00762_);
  or (_00765_, _00764_, _00761_);
  and (_00766_, _00151_, _00411_);
  and (_00767_, _00159_, _00415_);
  or (_00768_, _00767_, _00766_);
  and (_00769_, _00172_, _00408_);
  and (_00770_, _00176_, _00423_);
  or (_00771_, _00770_, _00769_);
  or (_00772_, _00771_, _00768_);
  or (_00773_, _00772_, _00765_);
  and (_00775_, _00218_, _00432_);
  and (_00777_, _00197_, _00437_);
  and (_00779_, _00200_, _00435_);
  or (_00781_, _00779_, _00777_);
  or (_00783_, _00781_, _00775_);
  and (_00785_, _00192_, _00391_);
  and (_00787_, _00189_, _00393_);
  or (_00788_, _00787_, _00785_);
  and (_00789_, _00180_, _00429_);
  and (_00790_, _00183_, _00389_);
  or (_00791_, _00790_, _00789_);
  or (_00792_, _00791_, _00788_);
  or (_00793_, _00792_, _00783_);
  or (_00795_, _00793_, _00773_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _00795_, _00758_);
  and (_00797_, _00172_, _00478_);
  and (_00798_, _00176_, _00465_);
  and (_00799_, _00151_, _00469_);
  and (_00800_, _00159_, _00473_);
  or (_00801_, _00800_, _00799_);
  or (_00802_, _00801_, _00798_);
  or (_00803_, _00802_, _00797_);
  and (_00804_, _00218_, _00488_);
  and (_00805_, _00200_, _00490_);
  or (_00806_, _00805_, _00804_);
  or (_00807_, _00806_, _00803_);
  and (_00808_, _00132_, _00452_);
  and (_00809_, _00141_, _00461_);
  and (_00810_, _00146_, _00480_);
  or (_00811_, _00810_, _00809_);
  and (_00812_, _00208_, _00454_);
  and (_00813_, _00214_, _00456_);
  or (_00814_, _00813_, _00812_);
  or (_00815_, _00814_, _00811_);
  and (_00816_, _00183_, _00444_);
  and (_00817_, _00189_, _00446_);
  and (_00818_, _00192_, _00448_);
  or (_00819_, _00818_, _00817_);
  or (_00820_, _00819_, _00816_);
  and (_00821_, _00180_, _00486_);
  and (_00822_, _00197_, _00492_);
  or (_00823_, _00822_, _00821_);
  or (_00824_, _00823_, _00820_);
  or (_00825_, _00824_, _00815_);
  or (_00827_, _00825_, _00808_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _00827_, _00807_);
  and (_00830_, _00214_, _00499_);
  and (_00832_, _00146_, _00548_);
  and (_00834_, _00141_, _00546_);
  or (_00836_, _00834_, _00832_);
  and (_00838_, _00132_, _00543_);
  and (_00839_, _00208_, _00541_);
  or (_00840_, _00839_, _00838_);
  or (_00841_, _00840_, _00836_);
  and (_00842_, _00151_, _00535_);
  and (_00843_, _00159_, _00532_);
  or (_00844_, _00843_, _00842_);
  and (_00846_, _00176_, _00528_);
  and (_00847_, _00172_, _00530_);
  or (_00849_, _00847_, _00846_);
  or (_00850_, _00849_, _00844_);
  or (_00851_, _00850_, _00841_);
  and (_00852_, _00218_, _00511_);
  and (_00853_, _00197_, _00517_);
  and (_00854_, _00200_, _00513_);
  or (_00855_, _00854_, _00853_);
  or (_00856_, _00855_, _00852_);
  and (_00857_, _00192_, _00505_);
  and (_00858_, _00189_, _00503_);
  or (_00859_, _00858_, _00857_);
  and (_00860_, _00180_, _00509_);
  and (_00861_, _00183_, _00501_);
  or (_00862_, _00861_, _00860_);
  or (_00863_, _00862_, _00859_);
  or (_00864_, _00863_, _00856_);
  or (_00865_, _00864_, _00851_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _00865_, _00830_);
  and (_00866_, _00214_, _00567_);
  and (_00867_, _00146_, _00590_);
  and (_00868_, _00141_, _00577_);
  or (_00869_, _00868_, _00867_);
  and (_00870_, _00208_, _00564_);
  and (_00871_, _00132_, _00562_);
  or (_00872_, _00871_, _00870_);
  or (_00873_, _00872_, _00869_);
  and (_00874_, _00151_, _00584_);
  and (_00875_, _00159_, _00582_);
  or (_00876_, _00875_, _00874_);
  and (_00878_, _00176_, _00580_);
  and (_00880_, _00172_, _00592_);
  or (_00882_, _00880_, _00878_);
  or (_00884_, _00882_, _00876_);
  or (_00886_, _00884_, _00873_);
  and (_00888_, _00218_, _00598_);
  and (_00890_, _00197_, _00602_);
  and (_00891_, _00200_, _00600_);
  or (_00892_, _00891_, _00890_);
  or (_00893_, _00892_, _00888_);
  and (_00894_, _00189_, _00558_);
  and (_00895_, _00192_, _00556_);
  or (_00896_, _00895_, _00894_);
  and (_00897_, _00183_, _00554_);
  and (_00898_, _00180_, _00596_);
  or (_00899_, _00898_, _00897_);
  or (_00900_, _00899_, _00896_);
  or (_00901_, _00900_, _00893_);
  or (_00902_, _00901_, _00886_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _00902_, _00866_);
  and (_00903_, _00214_, _00621_);
  and (_00904_, _00159_, _00637_);
  and (_00905_, _00151_, _00640_);
  or (_00906_, _00905_, _00904_);
  and (_00907_, _00176_, _00635_);
  and (_00908_, _00172_, _00645_);
  or (_00909_, _00908_, _00907_);
  or (_00910_, _00909_, _00906_);
  and (_00911_, _00146_, _00617_);
  and (_00912_, _00141_, _00633_);
  or (_00913_, _00912_, _00911_);
  and (_00914_, _00132_, _00647_);
  and (_00915_, _00208_, _00625_);
  or (_00916_, _00915_, _00914_);
  or (_00917_, _00916_, _00913_);
  or (_00918_, _00917_, _00910_);
  and (_00919_, _00218_, _00653_);
  and (_00921_, _00197_, _00657_);
  and (_00922_, _00200_, _00655_);
  or (_00923_, _00922_, _00921_);
  or (_00925_, _00923_, _00919_);
  and (_00926_, _00192_, _00613_);
  and (_00927_, _00189_, _00611_);
  or (_00929_, _00927_, _00926_);
  and (_00930_, _00180_, _00651_);
  and (_00931_, _00183_, _00609_);
  or (_00932_, _00931_, _00930_);
  or (_00933_, _00932_, _00929_);
  or (_00934_, _00933_, _00925_);
  or (_00935_, _00934_, _00918_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _00935_, _00903_);
  and (_00936_, _00200_, _00685_);
  and (_00937_, _00218_, _00683_);
  or (_00938_, _00937_, _00936_);
  and (_00939_, _00176_, _00702_);
  and (_00940_, _00159_, _00697_);
  and (_00941_, _00151_, _00699_);
  or (_00942_, _00941_, _00940_);
  or (_00943_, _00942_, _00939_);
  or (_00944_, _00943_, _00938_);
  and (_00945_, _00132_, _00706_);
  and (_00946_, _00141_, _00713_);
  and (_00947_, _00146_, _00711_);
  or (_00948_, _00947_, _00946_);
  and (_00949_, _00208_, _00708_);
  or (_00950_, _00949_, _00948_);
  and (_00951_, _00172_, _00695_);
  and (_00952_, _00214_, _00664_);
  or (_00953_, _00952_, _00951_);
  or (_00954_, _00953_, _00950_);
  and (_00955_, _00183_, _00666_);
  and (_00956_, _00192_, _00671_);
  and (_00957_, _00189_, _00668_);
  or (_00958_, _00957_, _00956_);
  or (_00959_, _00958_, _00955_);
  and (_00960_, _00180_, _00679_);
  and (_00961_, _00197_, _00687_);
  or (_00962_, _00961_, _00960_);
  or (_00963_, _00962_, _00959_);
  or (_00964_, _00963_, _00954_);
  or (_00965_, _00964_, _00945_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _00965_, _00944_);
  and (_00966_, _00180_, _00356_);
  and (_00967_, _00214_, _00346_);
  and (_00968_, _00218_, _00350_);
  or (_00969_, _00968_, _00967_);
  or (_00970_, _00969_, _00966_);
  and (_00971_, _00146_, _00383_);
  and (_00972_, _00197_, _00348_);
  and (_00973_, _00151_, _00359_);
  and (_00974_, _00132_, _00376_);
  or (_00975_, _00974_, _00973_);
  or (_00976_, _00975_, _00972_);
  or (_00977_, _00976_, _00971_);
  and (_00978_, _00159_, _00380_);
  and (_00979_, _00141_, _00374_);
  or (_00980_, _00979_, _00978_);
  or (_00981_, _00980_, _00977_);
  and (_00982_, _00172_, _00363_);
  and (_00983_, _00200_, _00340_);
  and (_00984_, _00192_, _00338_);
  or (_00985_, _00984_, _00983_);
  and (_00986_, _00183_, _00344_);
  and (_00987_, _00189_, _00336_);
  or (_00988_, _00987_, _00986_);
  or (_00989_, _00988_, _00985_);
  or (_00990_, _00989_, _00982_);
  and (_00991_, _00208_, _00334_);
  and (_00992_, _00176_, _00369_);
  or (_00993_, _00992_, _00991_);
  or (_00994_, _00993_, _00990_);
  or (_00995_, _00994_, _00981_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _00995_, _00970_);
  and (_00996_, _00208_, _00401_);
  and (_00997_, _00197_, _00435_);
  and (_00998_, _00214_, _00432_);
  or (_00999_, _00998_, _00997_);
  and (_01000_, _00218_, _00437_);
  and (_01001_, _00183_, _00429_);
  and (_01002_, _00192_, _00393_);
  or (_01003_, _01002_, _01001_);
  and (_01004_, _00189_, _00389_);
  and (_01005_, _00200_, _00391_);
  or (_01006_, _01005_, _01004_);
  or (_01007_, _01006_, _01003_);
  or (_01008_, _01007_, _01000_);
  or (_01009_, _01008_, _00999_);
  and (_01010_, _00151_, _00415_);
  and (_01011_, _00172_, _00411_);
  or (_01012_, _01011_, _01010_);
  and (_01013_, _00180_, _00423_);
  and (_01014_, _00176_, _00408_);
  or (_01015_, _01014_, _01013_);
  or (_01016_, _01015_, _01012_);
  and (_01017_, _00146_, _00406_);
  and (_01018_, _00159_, _00397_);
  or (_01019_, _01018_, _01017_);
  and (_01020_, _00132_, _00399_);
  and (_01021_, _00141_, _00425_);
  or (_01022_, _01021_, _01020_);
  or (_01023_, _01022_, _01019_);
  or (_01024_, _01023_, _01016_);
  or (_01025_, _01024_, _01009_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01025_, _00996_);
  and (_01026_, _00214_, _00488_);
  and (_01027_, _00197_, _00490_);
  or (_01028_, _01027_, _01026_);
  and (_01029_, _00218_, _00492_);
  and (_01030_, _00189_, _00444_);
  and (_01031_, _00192_, _00446_);
  or (_01032_, _01031_, _01030_);
  and (_01033_, _00183_, _00486_);
  and (_01034_, _00200_, _00448_);
  or (_01035_, _01034_, _01033_);
  or (_01036_, _01035_, _01032_);
  or (_01037_, _01036_, _01029_);
  or (_01038_, _01037_, _01028_);
  and (_01039_, _00132_, _00454_);
  and (_01040_, _00180_, _00465_);
  and (_01041_, _00151_, _00473_);
  and (_01042_, _00172_, _00469_);
  or (_01043_, _01042_, _01041_);
  or (_01044_, _01043_, _01040_);
  and (_01045_, _00208_, _00456_);
  and (_01046_, _00176_, _00478_);
  or (_01047_, _01046_, _01045_);
  and (_01048_, _00141_, _00452_);
  and (_01050_, _00159_, _00480_);
  and (_01051_, _00146_, _00461_);
  or (_01053_, _01051_, _01050_);
  or (_01054_, _01053_, _01048_);
  or (_01056_, _01054_, _01047_);
  or (_01057_, _01056_, _01044_);
  or (_01059_, _01057_, _01039_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01059_, _01038_);
  and (_01061_, _00214_, _00511_);
  and (_01062_, _00197_, _00513_);
  or (_01064_, _01062_, _01061_);
  and (_01065_, _00218_, _00517_);
  and (_01067_, _00183_, _00509_);
  and (_01068_, _00192_, _00503_);
  or (_01070_, _01068_, _01067_);
  and (_01071_, _00189_, _00501_);
  and (_01073_, _00200_, _00505_);
  or (_01074_, _01073_, _01071_);
  or (_01076_, _01074_, _01070_);
  or (_01077_, _01076_, _01065_);
  or (_01079_, _01077_, _01064_);
  and (_01080_, _00132_, _00541_);
  and (_01082_, _00176_, _00530_);
  and (_01083_, _00172_, _00535_);
  and (_01085_, _00151_, _00532_);
  or (_01086_, _01085_, _01083_);
  or (_01088_, _01086_, _01082_);
  and (_01089_, _00208_, _00499_);
  and (_01091_, _00180_, _00528_);
  or (_01092_, _01091_, _01089_);
  and (_01094_, _00159_, _00548_);
  and (_01095_, _00146_, _00546_);
  or (_01097_, _01095_, _01094_);
  and (_01098_, _00141_, _00543_);
  or (_01100_, _01098_, _01097_);
  or (_01101_, _01100_, _01092_);
  or (_01103_, _01101_, _01088_);
  or (_01104_, _01103_, _01080_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _01104_, _01079_);
  and (_01106_, _00214_, _00598_);
  and (_01108_, _00197_, _00600_);
  or (_01109_, _01108_, _01106_);
  and (_01110_, _00218_, _00602_);
  and (_01111_, _00183_, _00596_);
  and (_01112_, _00192_, _00558_);
  or (_01113_, _01112_, _01111_);
  and (_01114_, _00189_, _00554_);
  and (_01115_, _00200_, _00556_);
  or (_01116_, _01115_, _01114_);
  or (_01117_, _01116_, _01113_);
  or (_01118_, _01117_, _01110_);
  or (_01119_, _01118_, _01109_);
  and (_01120_, _00132_, _00564_);
  and (_01121_, _00180_, _00580_);
  and (_01122_, _00172_, _00584_);
  and (_01123_, _00151_, _00582_);
  or (_01124_, _01123_, _01122_);
  or (_01125_, _01124_, _01121_);
  and (_01126_, _00208_, _00567_);
  and (_01127_, _00176_, _00592_);
  or (_01128_, _01127_, _01126_);
  and (_01129_, _00159_, _00590_);
  and (_01130_, _00146_, _00577_);
  or (_01131_, _01130_, _01129_);
  and (_01132_, _00141_, _00562_);
  or (_01133_, _01132_, _01131_);
  or (_01134_, _01133_, _01128_);
  or (_01135_, _01134_, _01125_);
  or (_01136_, _01135_, _01120_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _01136_, _01119_);
  and (_01137_, _00208_, _00621_);
  and (_01138_, _00197_, _00655_);
  and (_01139_, _00214_, _00653_);
  or (_01140_, _01139_, _01138_);
  and (_01141_, _00218_, _00657_);
  and (_01142_, _00183_, _00651_);
  and (_01143_, _00192_, _00611_);
  or (_01144_, _01143_, _01142_);
  and (_01145_, _00189_, _00609_);
  and (_01146_, _00200_, _00613_);
  or (_01147_, _01146_, _01145_);
  or (_01148_, _01147_, _01144_);
  or (_01149_, _01148_, _01141_);
  or (_01150_, _01149_, _01140_);
  and (_01151_, _00146_, _00633_);
  and (_01152_, _00159_, _00617_);
  or (_01153_, _01152_, _01151_);
  and (_01154_, _00132_, _00625_);
  and (_01155_, _00141_, _00647_);
  or (_01156_, _01155_, _01154_);
  or (_01157_, _01156_, _01153_);
  and (_01158_, _00151_, _00637_);
  and (_01159_, _00172_, _00640_);
  or (_01160_, _01159_, _01158_);
  and (_01161_, _00176_, _00645_);
  and (_01162_, _00180_, _00635_);
  or (_01163_, _01162_, _01161_);
  or (_01164_, _01163_, _01160_);
  or (_01165_, _01164_, _01157_);
  or (_01166_, _01165_, _01150_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _01166_, _01137_);
  and (_01167_, _00218_, _00687_);
  and (_01168_, _00180_, _00702_);
  and (_01169_, _00214_, _00683_);
  or (_01170_, _01169_, _01168_);
  or (_01171_, _01170_, _01167_);
  and (_01172_, _00146_, _00713_);
  and (_01173_, _00197_, _00685_);
  and (_01174_, _00151_, _00697_);
  and (_01175_, _00132_, _00708_);
  or (_01176_, _01175_, _01174_);
  or (_01177_, _01176_, _01173_);
  or (_01178_, _01177_, _01172_);
  and (_01179_, _00159_, _00711_);
  and (_01180_, _00141_, _00706_);
  or (_01181_, _01180_, _01179_);
  or (_01182_, _01181_, _01178_);
  and (_01183_, _00172_, _00699_);
  and (_01184_, _00192_, _00668_);
  and (_01185_, _00200_, _00671_);
  or (_01186_, _01185_, _01184_);
  and (_01187_, _00183_, _00679_);
  and (_01188_, _00189_, _00666_);
  or (_01189_, _01188_, _01187_);
  or (_01190_, _01189_, _01186_);
  or (_01191_, _01190_, _01183_);
  and (_01192_, _00208_, _00664_);
  and (_01193_, _00176_, _00695_);
  or (_01194_, _01193_, _01192_);
  or (_01195_, _01194_, _01191_);
  or (_01196_, _01195_, _01182_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _01196_, _01171_);
  and (_01197_, _00214_, _00350_);
  and (_01198_, _00176_, _00363_);
  and (_01199_, _00218_, _00348_);
  or (_01200_, _01199_, _01198_);
  or (_01201_, _01200_, _01197_);
  and (_01202_, _00141_, _00376_);
  and (_01203_, _00146_, _00374_);
  or (_01204_, _01203_, _01202_);
  and (_01205_, _00159_, _00383_);
  and (_01206_, _00197_, _00340_);
  and (_01207_, _00132_, _00334_);
  and (_01208_, _00151_, _00380_);
  or (_01209_, _01208_, _01207_);
  or (_01210_, _01209_, _01206_);
  or (_01211_, _01210_, _01205_);
  or (_01212_, _01211_, _01204_);
  and (_01213_, _00180_, _00369_);
  and (_01214_, _00189_, _00344_);
  and (_01215_, _00192_, _00336_);
  or (_01216_, _01215_, _01214_);
  and (_01217_, _00183_, _00356_);
  and (_01218_, _00200_, _00338_);
  or (_01219_, _01218_, _01217_);
  or (_01220_, _01219_, _01216_);
  or (_01221_, _01220_, _01213_);
  and (_01222_, _00172_, _00359_);
  and (_01223_, _00208_, _00346_);
  or (_01224_, _01223_, _01222_);
  or (_01225_, _01224_, _01221_);
  or (_01226_, _01225_, _01212_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01226_, _01201_);
  and (_01227_, _00132_, _00401_);
  and (_01228_, _00146_, _00425_);
  and (_01229_, _00141_, _00399_);
  or (_01230_, _01229_, _01228_);
  and (_01231_, _00151_, _00397_);
  and (_01232_, _00159_, _00406_);
  or (_01233_, _01232_, _01231_);
  or (_01234_, _01233_, _01230_);
  and (_01235_, _00172_, _00415_);
  and (_01236_, _00176_, _00411_);
  or (_01237_, _01236_, _01235_);
  and (_01238_, _00180_, _00408_);
  and (_01239_, _00183_, _00423_);
  or (_01240_, _01239_, _01238_);
  or (_01241_, _01240_, _01237_);
  or (_01242_, _01241_, _01234_);
  and (_01243_, _00192_, _00389_);
  and (_01244_, _00189_, _00429_);
  or (_01245_, _01244_, _01243_);
  and (_01246_, _00197_, _00391_);
  and (_01247_, _00200_, _00393_);
  or (_01248_, _01247_, _01246_);
  or (_01249_, _01248_, _01245_);
  and (_01250_, _00218_, _00435_);
  and (_01251_, _00214_, _00437_);
  or (_01252_, _01251_, _01250_);
  and (_01253_, _00208_, _00432_);
  or (_01254_, _01253_, _01252_);
  or (_01255_, _01254_, _01249_);
  or (_01256_, _01255_, _01242_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01256_, _01227_);
  and (_01257_, _00208_, _00488_);
  and (_01258_, _00218_, _00490_);
  or (_01259_, _01258_, _01257_);
  and (_01260_, _00180_, _00478_);
  and (_01261_, _00176_, _00469_);
  and (_01262_, _00172_, _00473_);
  or (_01263_, _01262_, _01261_);
  or (_01264_, _01263_, _01260_);
  or (_01265_, _01264_, _01259_);
  and (_01266_, _00132_, _00456_);
  and (_01267_, _00159_, _00461_);
  and (_01268_, _00141_, _00454_);
  and (_01269_, _00146_, _00452_);
  or (_01270_, _01269_, _01268_);
  or (_01271_, _01270_, _01267_);
  and (_01272_, _00151_, _00480_);
  and (_01273_, _00183_, _00465_);
  or (_01274_, _01273_, _01272_);
  or (_01275_, _01274_, _01271_);
  and (_01276_, _00200_, _00446_);
  and (_01277_, _00192_, _00444_);
  and (_01278_, _00189_, _00486_);
  or (_01279_, _01278_, _01277_);
  or (_01280_, _01279_, _01276_);
  and (_01281_, _00214_, _00492_);
  and (_01282_, _00197_, _00448_);
  or (_01283_, _01282_, _01281_);
  or (_01284_, _01283_, _01280_);
  or (_01285_, _01284_, _01275_);
  or (_01286_, _01285_, _01266_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01286_, _01265_);
  and (_01287_, _00208_, _00511_);
  and (_01288_, _00218_, _00513_);
  or (_01289_, _01288_, _01287_);
  and (_01290_, _00180_, _00530_);
  and (_01291_, _00176_, _00535_);
  and (_01292_, _00172_, _00532_);
  or (_01293_, _01292_, _01291_);
  or (_01294_, _01293_, _01290_);
  or (_01295_, _01294_, _01289_);
  and (_01296_, _00132_, _00499_);
  and (_01297_, _00159_, _00546_);
  and (_01298_, _00141_, _00541_);
  and (_01299_, _00146_, _00543_);
  or (_01300_, _01299_, _01298_);
  or (_01301_, _01300_, _01297_);
  and (_01302_, _00151_, _00548_);
  and (_01303_, _00183_, _00528_);
  or (_01304_, _01303_, _01302_);
  or (_01305_, _01304_, _01301_);
  and (_01306_, _00200_, _00503_);
  and (_01307_, _00192_, _00501_);
  and (_01308_, _00189_, _00509_);
  or (_01309_, _01308_, _01307_);
  or (_01310_, _01309_, _01306_);
  and (_01311_, _00214_, _00517_);
  and (_01312_, _00197_, _00505_);
  or (_01313_, _01312_, _01311_);
  or (_01314_, _01313_, _01310_);
  or (_01315_, _01314_, _01305_);
  or (_01316_, _01315_, _01296_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01316_, _01295_);
  and (_01317_, _00214_, _00602_);
  and (_01318_, _00176_, _00584_);
  and (_01319_, _00208_, _00598_);
  or (_01320_, _01319_, _01318_);
  or (_01321_, _01320_, _01317_);
  and (_01322_, _00141_, _00564_);
  and (_01323_, _00197_, _00556_);
  and (_01324_, _00132_, _00567_);
  and (_01325_, _00151_, _00590_);
  or (_01326_, _01325_, _01324_);
  or (_01327_, _01326_, _01323_);
  or (_01328_, _01327_, _01322_);
  and (_01329_, _00146_, _00562_);
  and (_01330_, _00159_, _00577_);
  or (_01331_, _01330_, _01329_);
  or (_01332_, _01331_, _01328_);
  and (_01333_, _00180_, _00592_);
  and (_01334_, _00183_, _00580_);
  and (_01335_, _00192_, _00554_);
  or (_01336_, _01335_, _01334_);
  and (_01337_, _00189_, _00596_);
  and (_01338_, _00200_, _00558_);
  or (_01339_, _01338_, _01337_);
  or (_01340_, _01339_, _01336_);
  or (_01341_, _01340_, _01333_);
  and (_01342_, _00172_, _00582_);
  and (_01343_, _00218_, _00600_);
  or (_01344_, _01343_, _01342_);
  or (_01345_, _01344_, _01341_);
  or (_01346_, _01345_, _01332_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01346_, _01321_);
  and (_01347_, _00214_, _00657_);
  and (_01348_, _00176_, _00640_);
  and (_01349_, _00218_, _00655_);
  or (_01350_, _01349_, _01348_);
  or (_01351_, _01350_, _01347_);
  and (_01352_, _00141_, _00625_);
  and (_01353_, _00146_, _00647_);
  or (_01354_, _01353_, _01352_);
  and (_01355_, _00159_, _00633_);
  and (_01356_, _00197_, _00613_);
  and (_01357_, _00132_, _00621_);
  and (_01358_, _00151_, _00617_);
  or (_01359_, _01358_, _01357_);
  or (_01360_, _01359_, _01356_);
  or (_01361_, _01360_, _01355_);
  or (_01362_, _01361_, _01354_);
  and (_01363_, _00180_, _00645_);
  and (_01364_, _00189_, _00651_);
  and (_01365_, _00192_, _00609_);
  or (_01366_, _01365_, _01364_);
  and (_01367_, _00183_, _00635_);
  and (_01368_, _00200_, _00611_);
  or (_01369_, _01368_, _01367_);
  or (_01370_, _01369_, _01366_);
  or (_01371_, _01370_, _01363_);
  and (_01372_, _00172_, _00637_);
  and (_01373_, _00208_, _00653_);
  or (_01374_, _01373_, _01372_);
  or (_01375_, _01374_, _01371_);
  or (_01376_, _01375_, _01362_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01376_, _01351_);
  and (_01377_, _00132_, _00664_);
  and (_01378_, _00141_, _00708_);
  and (_01379_, _00146_, _00706_);
  or (_01380_, _01379_, _01378_);
  and (_01381_, _00151_, _00711_);
  and (_01382_, _00159_, _00713_);
  or (_01383_, _01382_, _01381_);
  or (_01384_, _01383_, _01380_);
  and (_01385_, _00172_, _00697_);
  and (_01386_, _00176_, _00699_);
  or (_01387_, _01386_, _01385_);
  and (_01388_, _00180_, _00695_);
  and (_01389_, _00183_, _00702_);
  or (_01390_, _01389_, _01388_);
  or (_01391_, _01390_, _01387_);
  or (_01392_, _01391_, _01384_);
  and (_01393_, _00189_, _00679_);
  and (_01394_, _00192_, _00666_);
  or (_01395_, _01394_, _01393_);
  and (_01396_, _00197_, _00671_);
  and (_01397_, _00200_, _00668_);
  or (_01398_, _01397_, _01396_);
  or (_01399_, _01398_, _01395_);
  and (_01400_, _00208_, _00683_);
  and (_01401_, _00214_, _00687_);
  and (_01402_, _00218_, _00685_);
  or (_01403_, _01402_, _01401_);
  or (_01404_, _01403_, _01400_);
  or (_01405_, _01404_, _01399_);
  or (_01406_, _01405_, _01392_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01406_, _01377_);
  nand (_01407_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_01408_, \oc8051_golden_model_1.PC [3]);
  or (_01409_, \oc8051_golden_model_1.PC [2], _01408_);
  or (_01410_, _01409_, _01407_);
  or (_01411_, _01410_, _39235_);
  not (_01412_, \oc8051_golden_model_1.PC [1]);
  or (_01413_, _01412_, \oc8051_golden_model_1.PC [0]);
  or (_01414_, _01413_, _01409_);
  or (_01415_, _01414_, _39194_);
  and (_01416_, _01415_, _01411_);
  not (_01417_, \oc8051_golden_model_1.PC [2]);
  or (_01418_, _01417_, \oc8051_golden_model_1.PC [3]);
  or (_01419_, _01418_, _01407_);
  or (_01420_, _01419_, _39071_);
  or (_01421_, _01418_, _01413_);
  or (_01422_, _01421_, _39025_);
  and (_01423_, _01422_, _01420_);
  and (_01424_, _01423_, _01416_);
  nand (_01425_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01426_, _01425_, _01407_);
  or (_01427_, _01426_, _39399_);
  or (_01428_, _01425_, _01413_);
  or (_01429_, _01428_, _39358_);
  and (_01430_, _01429_, _01427_);
  or (_01431_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01432_, _01431_, _01407_);
  or (_01433_, _01432_, _38892_);
  or (_01434_, _01431_, _01413_);
  or (_01435_, _01434_, _38851_);
  and (_01436_, _01435_, _01433_);
  and (_01437_, _01436_, _01430_);
  and (_01438_, _01437_, _01424_);
  not (_01439_, \oc8051_golden_model_1.PC [0]);
  or (_01440_, \oc8051_golden_model_1.PC [1], _01439_);
  or (_01441_, _01440_, _01425_);
  or (_01442_, _01441_, _39317_);
  or (_01443_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_01444_, _01443_, _01425_);
  or (_01445_, _01444_, _39276_);
  and (_01446_, _01445_, _01442_);
  or (_01447_, _01431_, _01443_);
  or (_01448_, _01447_, _38642_);
  or (_01449_, _01431_, _01440_);
  or (_01450_, _01449_, _38771_);
  and (_01451_, _01450_, _01448_);
  and (_01452_, _01451_, _01446_);
  or (_01453_, _01440_, _01409_);
  or (_01454_, _01453_, _39153_);
  or (_01455_, _01443_, _01409_);
  or (_01456_, _01455_, _39112_);
  and (_01457_, _01456_, _01454_);
  or (_01458_, _01440_, _01418_);
  or (_01459_, _01458_, _38976_);
  or (_01460_, _01443_, _01418_);
  or (_01461_, _01460_, _38933_);
  and (_01462_, _01461_, _01459_);
  and (_01463_, _01462_, _01457_);
  and (_01464_, _01463_, _01452_);
  and (_01465_, _01464_, _01438_);
  or (_01466_, _01410_, _39200_);
  or (_01467_, _01414_, _39159_);
  and (_01468_, _01467_, _01466_);
  or (_01469_, _01419_, _39036_);
  or (_01470_, _01421_, _38982_);
  and (_01471_, _01470_, _01469_);
  and (_01472_, _01471_, _01468_);
  or (_01473_, _01426_, _39364_);
  or (_01474_, _01428_, _39323_);
  and (_01475_, _01474_, _01473_);
  or (_01476_, _01432_, _38857_);
  or (_01477_, _01434_, _38793_);
  and (_01478_, _01477_, _01476_);
  and (_01479_, _01478_, _01475_);
  and (_01480_, _01479_, _01472_);
  or (_01481_, _01441_, _39282_);
  or (_01482_, _01444_, _39241_);
  and (_01483_, _01482_, _01481_);
  or (_01484_, _01447_, _38580_);
  or (_01485_, _01449_, _38659_);
  and (_01486_, _01485_, _01484_);
  and (_01487_, _01486_, _01483_);
  or (_01488_, _01453_, _39118_);
  or (_01489_, _01455_, _39077_);
  and (_01490_, _01489_, _01488_);
  or (_01491_, _01458_, _38940_);
  or (_01492_, _01460_, _38898_);
  and (_01493_, _01492_, _01491_);
  and (_01494_, _01493_, _01490_);
  and (_01495_, _01494_, _01487_);
  and (_01496_, _01495_, _01480_);
  and (_01497_, _01496_, _01465_);
  or (_01498_, _01410_, _39225_);
  or (_01499_, _01414_, _39184_);
  and (_01500_, _01499_, _01498_);
  or (_01501_, _01419_, _39061_);
  or (_01502_, _01421_, _39010_);
  and (_01503_, _01502_, _01501_);
  and (_01504_, _01503_, _01500_);
  or (_01505_, _01426_, _39389_);
  or (_01506_, _01428_, _39348_);
  and (_01507_, _01506_, _01505_);
  or (_01508_, _01432_, _38882_);
  or (_01509_, _01434_, _38841_);
  and (_01510_, _01509_, _01508_);
  and (_01511_, _01510_, _01507_);
  and (_01512_, _01511_, _01504_);
  or (_01513_, _01441_, _39307_);
  or (_01514_, _01444_, _39266_);
  and (_01515_, _01514_, _01513_);
  or (_01516_, _01447_, _38632_);
  or (_01517_, _01449_, _38737_);
  and (_01518_, _01517_, _01516_);
  and (_01519_, _01518_, _01515_);
  or (_01520_, _01453_, _39143_);
  or (_01521_, _01455_, _39102_);
  and (_01523_, _01521_, _01520_);
  or (_01525_, _01458_, _38965_);
  or (_01527_, _01460_, _38923_);
  and (_01528_, _01527_, _01525_);
  and (_01530_, _01528_, _01523_);
  and (_01531_, _01530_, _01519_);
  and (_01532_, _01531_, _01512_);
  or (_01533_, _01410_, _39230_);
  or (_01534_, _01414_, _39189_);
  and (_01535_, _01534_, _01533_);
  or (_01536_, _01419_, _39066_);
  or (_01537_, _01421_, _39015_);
  and (_01538_, _01537_, _01536_);
  and (_01539_, _01538_, _01535_);
  or (_01540_, _01426_, _39394_);
  or (_01541_, _01428_, _39353_);
  and (_01542_, _01541_, _01540_);
  or (_01543_, _01432_, _38887_);
  or (_01544_, _01434_, _38846_);
  and (_01545_, _01544_, _01543_);
  and (_01546_, _01545_, _01542_);
  and (_01547_, _01546_, _01539_);
  or (_01548_, _01441_, _39312_);
  or (_01549_, _01444_, _39271_);
  and (_01550_, _01549_, _01548_);
  or (_01551_, _01447_, _38637_);
  or (_01552_, _01449_, _38758_);
  and (_01553_, _01552_, _01551_);
  and (_01554_, _01553_, _01550_);
  or (_01555_, _01453_, _39148_);
  or (_01556_, _01455_, _39107_);
  and (_01557_, _01556_, _01555_);
  or (_01558_, _01458_, _38970_);
  or (_01559_, _01460_, _38928_);
  and (_01560_, _01559_, _01558_);
  and (_01561_, _01560_, _01557_);
  and (_01562_, _01561_, _01554_);
  nand (_01563_, _01562_, _01547_);
  or (_01564_, _01563_, _01532_);
  not (_01565_, _01564_);
  and (_01566_, _01565_, _01497_);
  or (_01567_, _01410_, _39205_);
  or (_01568_, _01414_, _39164_);
  and (_01569_, _01568_, _01567_);
  or (_01570_, _01419_, _39041_);
  or (_01571_, _01421_, _38987_);
  and (_01573_, _01571_, _01570_);
  and (_01574_, _01573_, _01569_);
  or (_01575_, _01426_, _39369_);
  or (_01576_, _01428_, _39328_);
  and (_01577_, _01576_, _01575_);
  or (_01578_, _01432_, _38862_);
  or (_01579_, _01434_, _38807_);
  and (_01580_, _01579_, _01578_);
  and (_01581_, _01580_, _01577_);
  and (_01582_, _01581_, _01574_);
  or (_01583_, _01441_, _39287_);
  or (_01584_, _01444_, _39246_);
  and (_01585_, _01584_, _01583_);
  or (_01586_, _01447_, _38612_);
  or (_01587_, _01449_, _38677_);
  and (_01588_, _01587_, _01586_);
  and (_01589_, _01588_, _01585_);
  or (_01590_, _01453_, _39123_);
  or (_01591_, _01455_, _39082_);
  and (_01592_, _01591_, _01590_);
  or (_01593_, _01458_, _38945_);
  or (_01594_, _01460_, _38903_);
  and (_01595_, _01594_, _01593_);
  and (_01596_, _01595_, _01592_);
  and (_01597_, _01596_, _01589_);
  and (_01598_, _01597_, _01582_);
  or (_01599_, _01410_, _39210_);
  or (_01600_, _01414_, _39169_);
  and (_01601_, _01600_, _01599_);
  or (_01602_, _01419_, _39046_);
  or (_01603_, _01421_, _38992_);
  and (_01604_, _01603_, _01602_);
  and (_01605_, _01604_, _01601_);
  or (_01606_, _01426_, _39374_);
  or (_01607_, _01428_, _39333_);
  and (_01608_, _01607_, _01606_);
  or (_01609_, _01432_, _38867_);
  or (_01610_, _01434_, _38826_);
  and (_01611_, _01610_, _01609_);
  and (_01612_, _01611_, _01608_);
  and (_01613_, _01612_, _01605_);
  or (_01614_, _01441_, _39292_);
  or (_01615_, _01444_, _39251_);
  and (_01616_, _01615_, _01614_);
  or (_01617_, _01447_, _38617_);
  or (_01618_, _01449_, _38690_);
  and (_01619_, _01618_, _01617_);
  and (_01620_, _01619_, _01616_);
  or (_01621_, _01453_, _39128_);
  or (_01622_, _01455_, _39087_);
  and (_01623_, _01622_, _01621_);
  or (_01624_, _01458_, _38950_);
  or (_01625_, _01460_, _38908_);
  and (_01626_, _01625_, _01624_);
  and (_01627_, _01626_, _01623_);
  and (_01628_, _01627_, _01620_);
  nand (_01629_, _01628_, _01613_);
  not (_01630_, _01629_);
  and (_01631_, _01630_, _01598_);
  or (_01632_, _01410_, _39215_);
  or (_01633_, _01414_, _39174_);
  and (_01634_, _01633_, _01632_);
  or (_01635_, _01419_, _39051_);
  or (_01636_, _01421_, _39000_);
  and (_01637_, _01636_, _01635_);
  and (_01638_, _01637_, _01634_);
  or (_01639_, _01426_, _39379_);
  or (_01640_, _01428_, _39338_);
  and (_01641_, _01640_, _01639_);
  or (_01642_, _01432_, _38872_);
  or (_01643_, _01434_, _38831_);
  and (_01644_, _01643_, _01642_);
  and (_01645_, _01644_, _01641_);
  and (_01646_, _01645_, _01638_);
  or (_01647_, _01441_, _39297_);
  or (_01648_, _01444_, _39256_);
  and (_01649_, _01648_, _01647_);
  or (_01650_, _01447_, _38622_);
  or (_01651_, _01449_, _38707_);
  and (_01652_, _01651_, _01650_);
  and (_01653_, _01652_, _01649_);
  or (_01654_, _01453_, _39133_);
  or (_01655_, _01455_, _39092_);
  and (_01656_, _01655_, _01654_);
  or (_01657_, _01458_, _38955_);
  or (_01658_, _01460_, _38913_);
  and (_01659_, _01658_, _01657_);
  and (_01660_, _01659_, _01656_);
  and (_01661_, _01660_, _01653_);
  nand (_01662_, _01661_, _01646_);
  or (_01663_, _01410_, _39220_);
  or (_01664_, _01414_, _39179_);
  and (_01665_, _01664_, _01663_);
  or (_01666_, _01419_, _39056_);
  or (_01667_, _01421_, _39005_);
  and (_01668_, _01667_, _01666_);
  and (_01669_, _01668_, _01665_);
  or (_01670_, _01426_, _39384_);
  or (_01671_, _01428_, _39343_);
  and (_01672_, _01671_, _01670_);
  or (_01673_, _01432_, _38877_);
  or (_01674_, _01434_, _38836_);
  and (_01675_, _01674_, _01673_);
  and (_01676_, _01675_, _01672_);
  and (_01677_, _01676_, _01669_);
  or (_01678_, _01441_, _39302_);
  or (_01679_, _01444_, _39261_);
  and (_01680_, _01679_, _01678_);
  or (_01681_, _01447_, _38627_);
  or (_01682_, _01449_, _38724_);
  and (_01683_, _01682_, _01681_);
  and (_01684_, _01683_, _01680_);
  or (_01685_, _01453_, _39138_);
  or (_01686_, _01455_, _39097_);
  and (_01687_, _01686_, _01685_);
  or (_01688_, _01458_, _38960_);
  or (_01689_, _01460_, _38918_);
  and (_01690_, _01689_, _01688_);
  and (_01691_, _01690_, _01687_);
  and (_01692_, _01691_, _01684_);
  nand (_01693_, _01692_, _01677_);
  or (_01694_, _01693_, _01662_);
  not (_01695_, _01694_);
  and (_01696_, _01695_, _01631_);
  and (_01697_, _01696_, _01566_);
  not (_01698_, _01697_);
  and (_01699_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_01700_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_01701_, _01700_, _01699_);
  not (_01702_, _01701_);
  or (_01703_, _01629_, _01598_);
  or (_01704_, _01703_, _01694_);
  not (_01705_, _01704_);
  nand (_01706_, _01531_, _01512_);
  or (_01707_, _01563_, _01706_);
  nand (_01708_, _01464_, _01438_);
  or (_01709_, _01496_, _01708_);
  nor (_01710_, _01709_, _01707_);
  and (_01711_, _01710_, _01705_);
  not (_01712_, _01711_);
  and (_01713_, _01496_, _01708_);
  and (_01714_, _01562_, _01547_);
  or (_01715_, _01714_, _01532_);
  not (_01716_, _01715_);
  and (_01717_, _01716_, _01713_);
  and (_01718_, _01717_, _01705_);
  or (_01719_, _01714_, _01706_);
  not (_01720_, _01719_);
  and (_01721_, _01720_, _01713_);
  and (_01722_, _01721_, _01705_);
  nor (_01723_, _01722_, _01718_);
  and (_01724_, _01723_, _01712_);
  and (_01725_, _01716_, _01497_);
  and (_01726_, _01725_, _01705_);
  and (_01727_, _01713_, _01565_);
  and (_01728_, _01727_, _01705_);
  nor (_01729_, _01728_, _01726_);
  not (_01730_, _01707_);
  and (_01731_, _01730_, _01497_);
  and (_01732_, _01731_, _01705_);
  and (_01733_, _01705_, _01566_);
  nor (_01734_, _01733_, _01732_);
  and (_01735_, _01713_, _01730_);
  and (_01736_, _01735_, _01705_);
  and (_01737_, _01720_, _01497_);
  and (_01738_, _01737_, _01705_);
  nor (_01739_, _01738_, _01736_);
  and (_01740_, _01739_, _01734_);
  and (_01741_, _01740_, _01729_);
  and (_01742_, _01741_, _01724_);
  or (_01743_, _01496_, _01465_);
  or (_01744_, _01743_, _01564_);
  or (_01745_, _01744_, _01704_);
  or (_01746_, _01743_, _01715_);
  or (_01747_, _01746_, _01704_);
  and (_01748_, _01747_, _01745_);
  or (_01749_, _01709_, _01715_);
  or (_01750_, _01749_, _01704_);
  or (_01751_, _01743_, _01719_);
  or (_01752_, _01751_, _01704_);
  and (_01753_, _01752_, _01750_);
  or (_01754_, _01709_, _01719_);
  or (_01755_, _01754_, _01704_);
  or (_01756_, _01743_, _01707_);
  or (_01757_, _01756_, _01704_);
  and (_01758_, _01757_, _01755_);
  and (_01759_, _01758_, _01753_);
  and (_01760_, _01759_, _01748_);
  not (_01761_, _01703_);
  not (_01762_, _01693_);
  and (_01763_, _01762_, _01662_);
  and (_01764_, _01763_, _01761_);
  and (_01765_, _01764_, _01710_);
  nor (_01766_, _01709_, _01564_);
  and (_01767_, _01766_, _01705_);
  nor (_01768_, _01767_, _01765_);
  and (_01769_, _01768_, _01760_);
  and (_01770_, _01769_, _01742_);
  or (_01771_, _01770_, _01702_);
  not (_01772_, _01710_);
  or (_01773_, _01630_, _01598_);
  or (_01774_, _01773_, _01694_);
  nor (_01775_, _01774_, _01772_);
  not (_01776_, _01775_);
  not (_01777_, _01766_);
  or (_01778_, _01774_, _01777_);
  nand (_01779_, _01759_, _01748_);
  nor (_01780_, _01407_, _01417_);
  and (_01781_, _01407_, _01417_);
  nor (_01782_, _01781_, _01780_);
  not (_01783_, _01782_);
  or (_01784_, _01783_, _01779_);
  nand (_01785_, _01784_, _01778_);
  and (_01786_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_01787_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_01788_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_01789_, _01788_, _01786_);
  and (_01790_, _01789_, _01787_);
  nor (_01791_, _01790_, _01786_);
  and (_01792_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_01793_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_01794_, _01793_, _01792_);
  not (_01795_, _01794_);
  nor (_01796_, _01795_, _01791_);
  and (_01797_, _01795_, _01791_);
  nor (_01798_, _01797_, _01796_);
  or (_01799_, _01798_, _01778_);
  and (_01800_, _01799_, _01768_);
  nand (_01801_, _01800_, _01785_);
  nand (_01802_, _01801_, _01776_);
  not (_01803_, _01742_);
  not (_01804_, \oc8051_golden_model_1.ACC [1]);
  and (_01805_, _01440_, _01413_);
  nor (_01806_, _01805_, _01804_);
  and (_01807_, \oc8051_golden_model_1.ACC [0], _01439_);
  and (_01808_, _01805_, _01804_);
  nor (_01809_, _01808_, _01806_);
  and (_01810_, _01809_, _01807_);
  nor (_01811_, _01810_, _01806_);
  and (_01812_, _01782_, \oc8051_golden_model_1.ACC [2]);
  nor (_01813_, _01782_, \oc8051_golden_model_1.ACC [2]);
  nor (_01814_, _01813_, _01812_);
  not (_01815_, _01814_);
  nor (_01816_, _01815_, _01811_);
  and (_01817_, _01815_, _01811_);
  nor (_01818_, _01817_, _01816_);
  nor (_01819_, _01818_, _01776_);
  nor (_01820_, _01819_, _01803_);
  nand (_01821_, _01820_, _01802_);
  and (_01822_, _01821_, _01771_);
  nor (_01823_, _01699_, \oc8051_golden_model_1.PC [3]);
  and (_01824_, _01699_, \oc8051_golden_model_1.PC [3]);
  nor (_01825_, _01824_, _01823_);
  or (_01826_, _01825_, _01770_);
  nor (_01827_, _01816_, _01812_);
  not (_01828_, _01419_);
  nor (_01829_, _01780_, _01408_);
  nor (_01830_, _01829_, _01828_);
  nor (_01831_, _01830_, \oc8051_golden_model_1.ACC [3]);
  and (_01832_, _01830_, \oc8051_golden_model_1.ACC [3]);
  nor (_01833_, _01832_, _01831_);
  and (_01834_, _01833_, _01827_);
  nor (_01835_, _01833_, _01827_);
  nor (_01836_, _01835_, _01834_);
  nor (_01837_, _01836_, _01776_);
  nor (_01838_, _01796_, _01792_);
  and (_01839_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_01840_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_01841_, _01840_, _01839_);
  not (_01842_, _01841_);
  nor (_01843_, _01842_, _01838_);
  and (_01844_, _01842_, _01838_);
  nor (_01845_, _01844_, _01843_);
  or (_01846_, _01845_, _01778_);
  and (_01847_, _01778_, _01830_);
  nand (_01848_, _01847_, _01760_);
  nand (_01849_, _01848_, _01846_);
  and (_01850_, _01776_, _01768_);
  and (_01851_, _01850_, _01849_);
  or (_01852_, _01851_, _01837_);
  nand (_01853_, _01852_, _01742_);
  nand (_01854_, _01853_, _01826_);
  or (_01855_, _01854_, _01822_);
  or (_01856_, _01742_, _01412_);
  or (_01857_, _01760_, \oc8051_golden_model_1.PC [1]);
  or (_01858_, _01805_, _01779_);
  nand (_01859_, _01858_, _01857_);
  nand (_01860_, _01859_, _01778_);
  nor (_01861_, _01789_, _01787_);
  nor (_01862_, _01861_, _01790_);
  not (_01863_, _01862_);
  or (_01864_, _01863_, _01778_);
  and (_01865_, _01864_, _01768_);
  nand (_01866_, _01865_, _01860_);
  or (_01867_, _01768_, _01412_);
  and (_01868_, _01867_, _01776_);
  nand (_01869_, _01868_, _01866_);
  nor (_01870_, _01809_, _01807_);
  nor (_01871_, _01870_, _01810_);
  and (_01872_, _01871_, _01775_);
  nor (_01873_, _01872_, _01803_);
  nand (_01874_, _01873_, _01869_);
  nand (_01875_, _01874_, _01856_);
  not (_01876_, _01778_);
  nor (_01877_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_01878_, _01877_, _01787_);
  nand (_01879_, _01878_, _01876_);
  and (_01880_, _01778_, _01439_);
  nand (_01881_, _01880_, _01760_);
  nand (_01882_, _01881_, _01879_);
  nand (_01883_, _01882_, _01768_);
  or (_01884_, _01769_, _01439_);
  nand (_01885_, _01884_, _01883_);
  nand (_01886_, _01885_, _01776_);
  not (_01887_, \oc8051_golden_model_1.ACC [0]);
  and (_01888_, _01887_, \oc8051_golden_model_1.PC [0]);
  or (_01889_, _01807_, _01776_);
  or (_01890_, _01889_, _01888_);
  and (_01891_, _01890_, _01742_);
  nand (_01892_, _01891_, _01886_);
  or (_01893_, _01742_, \oc8051_golden_model_1.PC [0]);
  nand (_01894_, _01893_, _01892_);
  or (_01895_, _01894_, _01875_);
  or (_01896_, _01895_, _01855_);
  or (_01897_, _01896_, _39364_);
  and (_01898_, _01874_, _01856_);
  or (_01899_, _01894_, _01898_);
  nand (_01900_, _01821_, _01771_);
  or (_01901_, _01854_, _01900_);
  or (_01902_, _01901_, _01899_);
  or (_01903_, _01902_, _39118_);
  and (_01904_, _01903_, _01897_);
  and (_01905_, _01893_, _01892_);
  or (_01906_, _01905_, _01875_);
  or (_01907_, _01901_, _01906_);
  or (_01908_, _01907_, _39159_);
  and (_01909_, _01853_, _01826_);
  or (_01910_, _01909_, _01900_);
  or (_01911_, _01910_, _01899_);
  or (_01912_, _01911_, _38659_);
  and (_01913_, _01912_, _01908_);
  and (_01914_, _01913_, _01904_);
  or (_01915_, _01906_, _01855_);
  or (_01916_, _01915_, _39323_);
  or (_01917_, _01899_, _01855_);
  or (_01918_, _01917_, _39282_);
  and (_01919_, _01918_, _01916_);
  or (_01920_, _01909_, _01822_);
  or (_01921_, _01920_, _01895_);
  or (_01922_, _01921_, _39036_);
  or (_01923_, _01905_, _01898_);
  or (_01924_, _01920_, _01923_);
  or (_01925_, _01924_, _38898_);
  and (_01926_, _01925_, _01922_);
  and (_01927_, _01926_, _01919_);
  and (_01928_, _01927_, _01914_);
  or (_01929_, _01920_, _01899_);
  or (_01930_, _01929_, _38940_);
  or (_01931_, _01910_, _01906_);
  or (_01932_, _01931_, _38793_);
  and (_01933_, _01932_, _01930_);
  or (_01934_, _01910_, _01895_);
  or (_01935_, _01934_, _38857_);
  or (_01936_, _01910_, _01923_);
  or (_01937_, _01936_, _38580_);
  and (_01938_, _01937_, _01935_);
  and (_01939_, _01938_, _01933_);
  or (_01940_, _01923_, _01855_);
  or (_01941_, _01940_, _39241_);
  or (_01942_, _01920_, _01906_);
  or (_01943_, _01942_, _38982_);
  and (_01944_, _01943_, _01941_);
  or (_01945_, _01901_, _01895_);
  or (_01946_, _01945_, _39200_);
  or (_01947_, _01901_, _01923_);
  or (_01948_, _01947_, _39077_);
  and (_01949_, _01948_, _01946_);
  and (_01950_, _01949_, _01944_);
  and (_01951_, _01950_, _01939_);
  nand (_01952_, _01951_, _01928_);
  or (_01953_, _01917_, _39302_);
  or (_01954_, _01921_, _39056_);
  and (_01955_, _01954_, _01953_);
  or (_01956_, _01929_, _38960_);
  or (_01957_, _01911_, _38724_);
  and (_01958_, _01957_, _01956_);
  and (_01959_, _01958_, _01955_);
  or (_01960_, _01945_, _39220_);
  or (_01961_, _01934_, _38877_);
  and (_01962_, _01961_, _01960_);
  or (_01963_, _01907_, _39179_);
  or (_01964_, _01947_, _39097_);
  and (_01965_, _01964_, _01963_);
  and (_01966_, _01965_, _01962_);
  and (_01967_, _01966_, _01959_);
  or (_01968_, _01942_, _39005_);
  or (_01969_, _01924_, _38918_);
  and (_01970_, _01969_, _01968_);
  or (_01971_, _01915_, _39343_);
  or (_01972_, _01936_, _38627_);
  and (_01973_, _01972_, _01971_);
  and (_01974_, _01973_, _01970_);
  or (_01975_, _01896_, _39384_);
  or (_01976_, _01931_, _38836_);
  and (_01977_, _01976_, _01975_);
  or (_01978_, _01940_, _39261_);
  or (_01979_, _01902_, _39138_);
  and (_01980_, _01979_, _01978_);
  and (_01981_, _01980_, _01977_);
  and (_01982_, _01981_, _01974_);
  and (_01983_, _01982_, _01967_);
  or (_01984_, _01983_, _01952_);
  nor (_01985_, _01984_, _01698_);
  not (_01986_, \oc8051_golden_model_1.SP [0]);
  and (_01987_, _01629_, _01598_);
  and (_01988_, _01987_, _01695_);
  and (_01989_, _01988_, _01566_);
  nor (_01990_, _01989_, _01733_);
  nor (_01991_, _01990_, _01986_);
  nor (_01992_, _01952_, _01698_);
  and (_01993_, _01726_, _01986_);
  and (_01994_, _01764_, _01717_);
  not (_01995_, _01994_);
  nor (_01996_, _01995_, _01952_);
  or (_01997_, _01934_, _38862_);
  or (_01998_, _01911_, _38677_);
  and (_01999_, _01998_, _01997_);
  or (_02000_, _01902_, _39123_);
  or (_02001_, _01931_, _38807_);
  and (_02002_, _02001_, _02000_);
  and (_02003_, _02002_, _01999_);
  or (_02004_, _01921_, _39041_);
  or (_02005_, _01942_, _38987_);
  and (_02006_, _02005_, _02004_);
  or (_02007_, _01896_, _39369_);
  or (_02008_, _01917_, _39287_);
  and (_02009_, _02008_, _02007_);
  and (_02010_, _02009_, _02006_);
  and (_02011_, _02010_, _02003_);
  or (_02012_, _01929_, _38945_);
  or (_02013_, _01936_, _38612_);
  and (_02014_, _02013_, _02012_);
  or (_02015_, _01945_, _39205_);
  or (_02016_, _01907_, _39164_);
  and (_02017_, _02016_, _02015_);
  and (_02018_, _02017_, _02014_);
  or (_02019_, _01915_, _39328_);
  or (_02020_, _01940_, _39246_);
  and (_02021_, _02020_, _02019_);
  or (_02022_, _01947_, _39082_);
  or (_02023_, _01924_, _38903_);
  and (_02024_, _02023_, _02022_);
  and (_02025_, _02024_, _02021_);
  and (_02026_, _02025_, _02018_);
  and (_02027_, _02026_, _02011_);
  not (_02028_, _02027_);
  and (_02029_, _02028_, _01996_);
  and (_02030_, _01763_, _01629_);
  and (_02031_, _02030_, _01710_);
  not (_02032_, _02031_);
  nor (_02033_, _02032_, _01952_);
  nor (_02034_, _01952_, _01772_);
  and (_02035_, _02034_, _01693_);
  nor (_02036_, _02035_, _02033_);
  not (_02037_, _01765_);
  nor (_02038_, _01952_, _02037_);
  not (_02039_, _02038_);
  and (_02040_, _02039_, _02036_);
  nor (_02041_, _02040_, _02028_);
  and (_02042_, _01988_, _01766_);
  not (_02043_, _02042_);
  nor (_02044_, _02043_, _01984_);
  not (_02045_, _01749_);
  and (_02046_, _01988_, _02045_);
  not (_02047_, _02046_);
  nor (_02048_, _02047_, _01984_);
  nor (_02049_, _02047_, _01952_);
  not (_02050_, _02049_);
  not (_02051_, _01756_);
  and (_02052_, _02051_, _01696_);
  and (_02053_, _01988_, _02051_);
  not (_02054_, _02053_);
  nor (_02055_, _02054_, _01984_);
  not (_02056_, _01744_);
  and (_02057_, _01988_, _02056_);
  not (_02058_, _02057_);
  or (_02059_, _02058_, _01984_);
  not (_02060_, _01747_);
  not (_02061_, _01746_);
  and (_02062_, _01764_, _02061_);
  not (_02063_, _02062_);
  nor (_02064_, _02063_, _01952_);
  and (_02065_, _02064_, _02028_);
  nor (_02066_, _02065_, _02060_);
  and (_02067_, _01693_, _01598_);
  and (_02068_, _02067_, _02061_);
  nor (_02069_, _02068_, _02064_);
  not (_02070_, _02069_);
  and (_02071_, _02070_, _02066_);
  nor (_02072_, _01747_, _01986_);
  and (_02073_, _02067_, _02056_);
  nor (_02074_, _02073_, _02072_);
  not (_02075_, _02074_);
  nor (_02076_, _02075_, _02071_);
  not (_02077_, _02076_);
  and (_02078_, _02030_, _02061_);
  and (_02079_, _02030_, _02056_);
  nor (_02080_, _02079_, _02078_);
  and (_02081_, _01764_, _01731_);
  not (_02082_, _02081_);
  and (_02083_, _01988_, _01737_);
  not (_02084_, _02083_);
  and (_02085_, _01764_, _01737_);
  and (_02086_, _02085_, _01983_);
  not (_02087_, _02085_);
  nor (_02088_, _01945_, _39235_);
  nor (_02089_, _01921_, _39071_);
  nor (_02090_, _02089_, _02088_);
  nor (_02091_, _01942_, _39025_);
  nor (_02092_, _01911_, _38771_);
  nor (_02093_, _02092_, _02091_);
  and (_02094_, _02093_, _02090_);
  nor (_02095_, _01896_, _39399_);
  nor (_02096_, _01934_, _38892_);
  nor (_02097_, _02096_, _02095_);
  nor (_02098_, _01915_, _39358_);
  nor (_02099_, _01902_, _39153_);
  nor (_02100_, _02099_, _02098_);
  and (_02101_, _02100_, _02097_);
  and (_02102_, _02101_, _02094_);
  nor (_02103_, _01929_, _38976_);
  nor (_02104_, _01924_, _38933_);
  nor (_02105_, _02104_, _02103_);
  nor (_02106_, _01907_, _39194_);
  nor (_02107_, _01936_, _38642_);
  nor (_02108_, _02107_, _02106_);
  and (_02109_, _02108_, _02105_);
  nor (_02110_, _01917_, _39317_);
  nor (_02111_, _01931_, _38851_);
  nor (_02112_, _02111_, _02110_);
  nor (_02113_, _01940_, _39276_);
  nor (_02114_, _01947_, _39112_);
  nor (_02115_, _02114_, _02113_);
  and (_02116_, _02115_, _02112_);
  and (_02117_, _02116_, _02109_);
  and (_02118_, _02117_, _02102_);
  nor (_02119_, _02118_, _01952_);
  not (_02120_, _01983_);
  and (_02121_, _02120_, _01952_);
  nor (_02122_, _02121_, _02119_);
  and (_02123_, _01988_, _01717_);
  and (_02124_, _01988_, _01710_);
  nor (_02125_, _02124_, _02123_);
  not (_02126_, _02125_);
  and (_02127_, _02126_, _02122_);
  not (_02128_, _01754_);
  nor (_02129_, _01762_, _01662_);
  and (_02130_, _02129_, _01629_);
  and (_02131_, _02130_, _02128_);
  and (_02132_, _02129_, _01631_);
  and (_02133_, _02129_, _01761_);
  nor (_02134_, _02133_, _02132_);
  nor (_02135_, _02134_, _01754_);
  nor (_02136_, _02135_, _02131_);
  and (_02137_, _01693_, _01662_);
  and (_02138_, _02137_, _01631_);
  and (_02139_, _02138_, _02128_);
  not (_02140_, _02137_);
  or (_02141_, _02140_, _01631_);
  nor (_02142_, _02141_, _01754_);
  nor (_02143_, _02142_, _02139_);
  and (_02144_, _02143_, _02136_);
  not (_02145_, _02144_);
  and (_02146_, _02145_, _01983_);
  and (_02147_, _02045_, _01696_);
  nor (_02148_, _02147_, _02046_);
  nor (_02149_, _02148_, _02122_);
  nor (_02150_, _02057_, _02053_);
  not (_02151_, _02150_);
  and (_02152_, _02151_, _02122_);
  and (_02153_, _01764_, _02051_);
  and (_02154_, _02153_, _01983_);
  and (_02155_, _02056_, _01696_);
  and (_02156_, _02155_, \oc8051_golden_model_1.SP [3]);
  nor (_02157_, _02156_, _02153_);
  and (_02158_, _01764_, _02056_);
  not (_02159_, _01751_);
  and (_02160_, _01764_, _02159_);
  nor (_02161_, _02160_, _02158_);
  or (_02162_, _02161_, _01983_);
  nand (_02163_, _02161_, \oc8051_golden_model_1.PSW [3]);
  and (_02164_, _02163_, _02058_);
  and (_02165_, _02164_, _02162_);
  or (_02166_, _02165_, _02155_);
  and (_02167_, _02166_, _02157_);
  or (_02168_, _02167_, _02154_);
  and (_02169_, _02168_, _02054_);
  nor (_02170_, _02169_, _02152_);
  and (_02171_, _01764_, _02045_);
  nor (_02172_, _02171_, _02052_);
  not (_02173_, _02172_);
  nor (_02174_, _02173_, _02170_);
  and (_02175_, _02173_, _01983_);
  nor (_02176_, _02175_, _02174_);
  and (_02177_, _02176_, _02148_);
  or (_02178_, _02177_, _02145_);
  nor (_02179_, _02178_, _02149_);
  nor (_02180_, _02179_, _02146_);
  and (_02181_, _02128_, _01696_);
  and (_02182_, _01988_, _02128_);
  nor (_02183_, _02182_, _02181_);
  not (_02184_, _02183_);
  nor (_02185_, _02184_, _02180_);
  and (_02186_, _01766_, _01764_);
  and (_02187_, _02184_, _02122_);
  nor (_02188_, _02187_, _02186_);
  not (_02189_, _02188_);
  or (_02190_, _02189_, _02185_);
  not (_02191_, _02186_);
  nor (_02192_, _02191_, _01983_);
  nor (_02193_, _02192_, _02042_);
  nand (_02194_, _02193_, _02190_);
  and (_02195_, _02122_, _02042_);
  nor (_02196_, _02195_, _01765_);
  nand (_02197_, _02196_, _02194_);
  and (_02198_, _01988_, _01731_);
  nor (_02199_, _02198_, _01697_);
  and (_02200_, _01725_, _01696_);
  not (_02201_, _01774_);
  and (_02202_, _02201_, _01735_);
  nor (_02203_, _02202_, _02200_);
  and (_02204_, _02203_, _02199_);
  and (_02206_, _02201_, _01727_);
  not (_02208_, _02206_);
  and (_02210_, _02201_, _01721_);
  nor (_02212_, _02210_, _01994_);
  and (_02214_, _02212_, _02208_);
  and (_02216_, _02214_, _02204_);
  and (_02218_, _01766_, _01696_);
  and (_02219_, _02137_, _01987_);
  and (_02220_, _02219_, _02045_);
  nor (_02221_, _02220_, _02218_);
  and (_02222_, _01987_, _01763_);
  and (_02223_, _02222_, _02045_);
  nor (_02224_, _02223_, _02171_);
  and (_02225_, _02224_, _02221_);
  and (_02226_, _02225_, _02216_);
  and (_02227_, _02130_, _02045_);
  and (_02228_, _02138_, _02045_);
  nor (_02229_, _02228_, _02227_);
  and (_02230_, _02132_, _02045_);
  and (_02231_, _02133_, _02045_);
  or (_02232_, _02231_, _02230_);
  not (_02233_, _02232_);
  and (_02234_, _02233_, _02229_);
  not (_02235_, _01773_);
  and (_02236_, _02235_, _01763_);
  and (_02237_, _02236_, _02045_);
  not (_02238_, _02237_);
  nor (_02239_, _02140_, _01773_);
  and (_02240_, _02239_, _02045_);
  nor (_02241_, _02240_, _02158_);
  and (_02242_, _02241_, _02238_);
  and (_02243_, _01737_, _01696_);
  nor (_02244_, _02243_, _01989_);
  and (_02245_, _01763_, _01631_);
  and (_02246_, _02245_, _02045_);
  and (_02247_, _02137_, _01761_);
  and (_02248_, _02247_, _02045_);
  nor (_02249_, _02248_, _02246_);
  and (_02250_, _02249_, _02244_);
  and (_02251_, _02250_, _02242_);
  and (_02252_, _02251_, _02234_);
  and (_02253_, _02252_, _02226_);
  nor (_02254_, _02253_, _01439_);
  and (_02255_, _02253_, _01439_);
  nor (_02256_, _02255_, _02254_);
  nor (_02257_, _02255_, _01412_);
  and (_02258_, _02255_, _01412_);
  nor (_02259_, _02258_, _02257_);
  nor (_02260_, _02259_, _02256_);
  nor (_02261_, _02253_, _01702_);
  and (_02262_, _02253_, _01782_);
  nor (_02263_, _02262_, _02261_);
  not (_02264_, _01825_);
  nor (_02265_, _02253_, _02264_);
  not (_02266_, _01830_);
  and (_02267_, _02253_, _02266_);
  nor (_02268_, _02267_, _02265_);
  and (_02269_, _02268_, _02263_);
  and (_02270_, _02269_, _02260_);
  and (_02271_, _02270_, _00517_);
  and (_02272_, _02259_, _02256_);
  and (_02273_, _02272_, _02269_);
  and (_02274_, _02273_, _00513_);
  nor (_02275_, _02274_, _02271_);
  nor (_02276_, _02268_, _02263_);
  and (_02277_, _02276_, _02260_);
  and (_02278_, _02277_, _00543_);
  not (_02279_, _02256_);
  nor (_02280_, _02259_, _02279_);
  and (_02281_, _02280_, _02276_);
  and (_02282_, _02281_, _00546_);
  nor (_02283_, _02282_, _02278_);
  and (_02284_, _02283_, _02275_);
  and (_02285_, _02259_, _02279_);
  and (_02286_, _02285_, _02269_);
  and (_02287_, _02286_, _00505_);
  not (_02288_, _02268_);
  nor (_02289_, _02288_, _02263_);
  and (_02290_, _02289_, _02280_);
  and (_02291_, _02290_, _00503_);
  nor (_02292_, _02291_, _02287_);
  and (_02293_, _02288_, _02263_);
  and (_02294_, _02293_, _02285_);
  and (_02295_, _02294_, _00548_);
  and (_02296_, _02293_, _02280_);
  and (_02297_, _02296_, _00530_);
  nor (_02298_, _02297_, _02295_);
  and (_02299_, _02298_, _02292_);
  and (_02300_, _02299_, _02284_);
  and (_02301_, _02289_, _02272_);
  and (_02302_, _02301_, _00509_);
  and (_02303_, _02289_, _02260_);
  and (_02304_, _02303_, _00501_);
  nor (_02305_, _02304_, _02302_);
  and (_02306_, _02285_, _02276_);
  and (_02307_, _02306_, _00499_);
  and (_02308_, _02276_, _02272_);
  and (_02309_, _02308_, _00541_);
  nor (_02310_, _02309_, _02307_);
  and (_02311_, _02310_, _02305_);
  and (_02312_, _02293_, _02272_);
  and (_02313_, _02312_, _00532_);
  and (_02314_, _02280_, _02269_);
  and (_02315_, _02314_, _00511_);
  nor (_02316_, _02315_, _02313_);
  and (_02317_, _02293_, _02260_);
  and (_02318_, _02317_, _00535_);
  and (_02319_, _02289_, _02285_);
  and (_02320_, _02319_, _00528_);
  nor (_02321_, _02320_, _02318_);
  and (_02322_, _02321_, _02316_);
  and (_02323_, _02322_, _02311_);
  and (_02324_, _02323_, _02300_);
  nor (_02325_, _02324_, _02037_);
  nor (_02326_, _02325_, _02126_);
  and (_02327_, _02326_, _02197_);
  or (_02328_, _02327_, _02127_);
  and (_02329_, _01764_, _01721_);
  not (_02330_, _02329_);
  and (_02331_, _01988_, _01721_);
  nor (_02332_, _02331_, _02210_);
  and (_02333_, _02332_, _02330_);
  and (_02334_, _01988_, _01735_);
  nor (_02335_, _02334_, _02202_);
  and (_02336_, _01764_, _01735_);
  not (_02337_, _02336_);
  and (_02338_, _02337_, _02335_);
  and (_02339_, _02338_, _02333_);
  and (_02340_, _01764_, _01727_);
  not (_02341_, _02340_);
  and (_02342_, _01988_, _01727_);
  nor (_02343_, _02342_, _02206_);
  and (_02344_, _02343_, _02341_);
  and (_02345_, _01764_, _01725_);
  not (_02346_, _02345_);
  and (_02347_, _02346_, _02344_);
  and (_02348_, _02347_, _02339_);
  nand (_02349_, _02348_, _02328_);
  and (_02350_, _01988_, _01725_);
  nor (_02351_, _02348_, _02120_);
  nor (_02352_, _02351_, _02350_);
  and (_02353_, _02352_, _02349_);
  and (_02354_, _02350_, \oc8051_golden_model_1.SP [3]);
  or (_02355_, _02354_, _02200_);
  nor (_02356_, _02355_, _02353_);
  and (_02357_, _02122_, _02200_);
  or (_02358_, _02357_, _02356_);
  and (_02359_, _02358_, _02087_);
  or (_02360_, _02359_, _02086_);
  nand (_02361_, _02360_, _02084_);
  not (_02362_, \oc8051_golden_model_1.SP [3]);
  and (_02363_, _02083_, _02362_);
  nor (_02364_, _02363_, _02243_);
  nand (_02365_, _02364_, _02361_);
  and (_02366_, _01764_, _01566_);
  not (_02367_, _02243_);
  nor (_02368_, _02367_, _02122_);
  nor (_02369_, _02368_, _02366_);
  nand (_02370_, _02369_, _02365_);
  and (_02371_, _02366_, _01983_);
  nor (_02372_, _02371_, _01697_);
  and (_02373_, _02372_, _02370_);
  nor (_02374_, _02122_, _01698_);
  or (_02375_, _02374_, _02373_);
  nand (_02376_, _02375_, _02082_);
  nor (_02377_, _02082_, _01983_);
  not (_02378_, _02377_);
  and (_02379_, _02378_, _02376_);
  nor (_02380_, _01945_, _39230_);
  nor (_02381_, _01907_, _39189_);
  nor (_02382_, _02381_, _02380_);
  nor (_02383_, _01940_, _39271_);
  nor (_02384_, _01902_, _39148_);
  nor (_02385_, _02384_, _02383_);
  and (_02386_, _02385_, _02382_);
  nor (_02387_, _01921_, _39066_);
  nor (_02388_, _01942_, _39015_);
  nor (_02389_, _02388_, _02387_);
  nor (_02390_, _01929_, _38970_);
  nor (_02391_, _01931_, _38846_);
  nor (_02392_, _02391_, _02390_);
  and (_02393_, _02392_, _02389_);
  and (_02394_, _02393_, _02386_);
  nor (_02395_, _01917_, _39312_);
  nor (_02396_, _01936_, _38637_);
  nor (_02397_, _02396_, _02395_);
  nor (_02398_, _01947_, _39107_);
  nor (_02399_, _01934_, _38887_);
  nor (_02400_, _02399_, _02398_);
  and (_02401_, _02400_, _02397_);
  nor (_02402_, _01896_, _39394_);
  nor (_02403_, _01911_, _38758_);
  nor (_02404_, _02403_, _02402_);
  nor (_02405_, _01915_, _39353_);
  nor (_02406_, _01924_, _38928_);
  nor (_02407_, _02406_, _02405_);
  and (_02408_, _02407_, _02404_);
  and (_02409_, _02408_, _02401_);
  and (_02410_, _02409_, _02394_);
  nor (_02411_, _02410_, _01952_);
  and (_02412_, _02183_, _02148_);
  and (_02413_, _02150_, _02125_);
  and (_02414_, _02413_, _02412_);
  nor (_02415_, _02042_, _01697_);
  nor (_02416_, _02243_, _02200_);
  and (_02417_, _02416_, _02415_);
  and (_02418_, _02417_, _02414_);
  not (_02419_, _02418_);
  and (_02420_, _02419_, _02411_);
  not (_02421_, _02420_);
  nor (_02422_, _01917_, _39297_);
  nor (_02423_, _01911_, _38707_);
  nor (_02424_, _02423_, _02422_);
  nor (_02425_, _01940_, _39256_);
  nor (_02426_, _01921_, _39051_);
  nor (_02427_, _02426_, _02425_);
  and (_02428_, _02427_, _02424_);
  nor (_02429_, _01915_, _39338_);
  nor (_02430_, _01907_, _39174_);
  nor (_02431_, _02430_, _02429_);
  nor (_02432_, _01934_, _38872_);
  nor (_02433_, _01936_, _38622_);
  nor (_02434_, _02433_, _02432_);
  and (_02435_, _02434_, _02431_);
  and (_02436_, _02435_, _02428_);
  nor (_02437_, _01902_, _39133_);
  nor (_02438_, _01929_, _38955_);
  nor (_02439_, _02438_, _02437_);
  nor (_02440_, _01896_, _39379_);
  nor (_02441_, _01945_, _39215_);
  nor (_02442_, _02441_, _02440_);
  and (_02443_, _02442_, _02439_);
  nor (_02444_, _01947_, _39092_);
  nor (_02445_, _01924_, _38913_);
  nor (_02446_, _02445_, _02444_);
  nor (_02447_, _01942_, _39000_);
  nor (_02448_, _01931_, _38831_);
  nor (_02449_, _02448_, _02447_);
  and (_02450_, _02449_, _02446_);
  and (_02451_, _02450_, _02443_);
  and (_02452_, _02451_, _02436_);
  not (_02453_, _02452_);
  nor (_02454_, _02186_, _02153_);
  and (_02455_, _02454_, _02172_);
  and (_02456_, _02455_, _02161_);
  nand (_02457_, _02456_, _02144_);
  nor (_02458_, _02366_, _02081_);
  and (_02459_, _02458_, _02087_);
  nand (_02460_, _02459_, _02348_);
  or (_02461_, _02460_, _02457_);
  and (_02462_, _02461_, _02453_);
  not (_02463_, _02462_);
  and (_02464_, _02308_, _00454_);
  and (_02465_, _02277_, _00452_);
  nor (_02466_, _02465_, _02464_);
  and (_02467_, _02314_, _00488_);
  and (_02468_, _02273_, _00490_);
  nor (_02469_, _02468_, _02467_);
  and (_02470_, _02469_, _02466_);
  and (_02471_, _02294_, _00480_);
  and (_02472_, _02317_, _00469_);
  nor (_02473_, _02472_, _02471_);
  and (_02474_, _02290_, _00446_);
  and (_02475_, _02270_, _00492_);
  nor (_02476_, _02475_, _02474_);
  and (_02477_, _02476_, _02473_);
  and (_02478_, _02477_, _02470_);
  and (_02479_, _02301_, _00486_);
  and (_02480_, _02303_, _00444_);
  nor (_02481_, _02480_, _02479_);
  and (_02482_, _02306_, _00456_);
  and (_02483_, _02281_, _00461_);
  nor (_02484_, _02483_, _02482_);
  and (_02485_, _02484_, _02481_);
  and (_02486_, _02319_, _00465_);
  and (_02487_, _02296_, _00478_);
  nor (_02488_, _02487_, _02486_);
  and (_02489_, _02312_, _00473_);
  and (_02490_, _02286_, _00448_);
  nor (_02491_, _02490_, _02489_);
  and (_02492_, _02491_, _02488_);
  and (_02493_, _02492_, _02485_);
  and (_02494_, _02493_, _02478_);
  nor (_02495_, _02494_, _02037_);
  and (_02496_, _01693_, _01630_);
  and (_02497_, _02496_, _01662_);
  not (_02498_, _02497_);
  not (_02499_, _01737_);
  nor (_02500_, _01721_, _01725_);
  and (_02501_, _02500_, _02499_);
  nor (_02502_, _02501_, _02498_);
  not (_02503_, _02502_);
  nor (_02504_, _02045_, _01735_);
  nor (_02505_, _02159_, _01566_);
  and (_02506_, _02505_, _02504_);
  nor (_02507_, _02506_, _02140_);
  not (_02508_, _02507_);
  and (_02509_, _02497_, _01766_);
  not (_02510_, _02509_);
  nor (_02511_, _02140_, _01744_);
  and (_02512_, _02137_, _01629_);
  and (_02513_, _02512_, _01737_);
  nor (_02514_, _02513_, _02511_);
  and (_02515_, _02514_, _02510_);
  and (_02516_, _02515_, _02508_);
  and (_02517_, _02516_, _02503_);
  not (_02518_, \oc8051_golden_model_1.SP [2]);
  not (_02519_, _02155_);
  nor (_02520_, _02350_, _02083_);
  and (_02521_, _02520_, _02519_);
  nor (_02522_, _02521_, _02518_);
  not (_02523_, _02522_);
  not (_02524_, _02512_);
  nor (_02525_, _02500_, _02524_);
  not (_02526_, _02525_);
  and (_02527_, _02137_, _01731_);
  and (_02528_, _02497_, _02051_);
  nor (_02529_, _02528_, _02527_);
  and (_02530_, _02529_, _02526_);
  and (_02531_, _01777_, _01756_);
  nor (_02532_, _02531_, _02524_);
  nor (_02533_, _01710_, _01727_);
  nor (_02534_, _02533_, _02140_);
  nor (_02535_, _02534_, _02532_);
  and (_02536_, _02535_, _02530_);
  and (_02537_, _02536_, _02523_);
  and (_02538_, _02537_, _02517_);
  not (_02539_, _02538_);
  nor (_02540_, _02539_, _02495_);
  and (_02541_, _02540_, _02463_);
  and (_02542_, _02541_, _02421_);
  not (_02543_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_02544_, _02082_, _02027_);
  not (_02545_, _02544_);
  nor (_02546_, _02183_, _01984_);
  not (_02547_, _02171_);
  nor (_02548_, _02547_, _02027_);
  not (_02549_, _02153_);
  or (_02550_, _02549_, _02027_);
  nor (_02551_, _02161_, _02027_);
  and (_02552_, _02030_, _02159_);
  nand (_02553_, _01693_, _01629_);
  nor (_02554_, _02553_, _01751_);
  or (_02555_, _02554_, _02078_);
  or (_02556_, _02555_, _02552_);
  and (_02557_, _02556_, _01598_);
  and (_02558_, _02138_, _02159_);
  and (_02559_, _01988_, _02061_);
  and (_02560_, _02132_, _02159_);
  or (_02561_, _02560_, _02160_);
  or (_02562_, _02561_, _02559_);
  or (_02563_, _02562_, _02558_);
  nor (_02564_, _02563_, _02557_);
  and (_02565_, _02512_, _02056_);
  or (_02566_, _02565_, _02079_);
  and (_02567_, _02566_, _01598_);
  and (_02568_, _02138_, _02056_);
  and (_02569_, _01988_, _02159_);
  and (_02570_, _02129_, _01598_);
  and (_02571_, _02570_, _02056_);
  or (_02572_, _02571_, _02158_);
  or (_02573_, _02572_, _02569_);
  or (_02574_, _02573_, _02568_);
  nor (_02575_, _02574_, _02567_);
  and (_02576_, _02575_, _02564_);
  or (_02577_, _02576_, _02551_);
  nand (_02578_, _02577_, _02058_);
  nand (_02579_, _02059_, _02578_);
  and (_02580_, _02130_, _02051_);
  and (_02581_, _02512_, _02051_);
  and (_02582_, _02030_, _02051_);
  or (_02583_, _02582_, _02581_);
  or (_02584_, _02583_, _02580_);
  and (_02585_, _02584_, _01598_);
  not (_02586_, _02585_);
  and (_02587_, _02155_, _01986_);
  nor (_02588_, _02587_, _02153_);
  and (_02589_, _02138_, _02051_);
  and (_02590_, _02132_, _02051_);
  nor (_02591_, _02590_, _02589_);
  and (_02592_, _02591_, _02588_);
  and (_02593_, _02592_, _02586_);
  nand (_02594_, _02593_, _02579_);
  nand (_02595_, _02594_, _02550_);
  and (_02596_, _02595_, _02054_);
  or (_02597_, _02055_, _02596_);
  and (_02598_, _02052_, _02027_);
  and (_02599_, _02129_, _01987_);
  and (_02600_, _02599_, _02045_);
  nor (_02601_, _02600_, _02228_);
  nor (_02602_, _02230_, _02220_);
  and (_02603_, _02602_, _02601_);
  and (_02604_, _02603_, _02224_);
  not (_02605_, _02604_);
  nor (_02606_, _02605_, _02598_);
  and (_02607_, _02606_, _02597_);
  or (_02608_, _02607_, _02548_);
  nand (_02609_, _02608_, _02148_);
  nor (_02610_, _02148_, _01984_);
  nor (_02611_, _02610_, _02145_);
  nand (_02612_, _02611_, _02609_);
  and (_02613_, _02145_, _02027_);
  and (_02614_, _02222_, _02128_);
  not (_02615_, _02614_);
  and (_02616_, _02615_, _02183_);
  not (_02617_, _02616_);
  nor (_02618_, _02617_, _02613_);
  and (_02619_, _02618_, _02612_);
  or (_02620_, _02619_, _02546_);
  and (_02621_, _02219_, _01766_);
  nor (_02622_, _02621_, _02186_);
  and (_02623_, _02222_, _01766_);
  not (_02624_, _02623_);
  and (_02625_, _02132_, _01766_);
  not (_02626_, _02625_);
  and (_02627_, _02138_, _01766_);
  and (_02628_, _02599_, _01766_);
  nor (_02629_, _02628_, _02627_);
  and (_02630_, _02629_, _02626_);
  and (_02631_, _02630_, _02624_);
  and (_02632_, _02631_, _02622_);
  and (_02633_, _02632_, _02620_);
  nor (_02634_, _02191_, _02027_);
  or (_02635_, _02634_, _02633_);
  and (_02636_, _02635_, _02043_);
  or (_02637_, _02636_, _02044_);
  and (_02638_, _02512_, _01710_);
  and (_02639_, _02130_, _01710_);
  or (_02640_, _02639_, _02031_);
  or (_02641_, _02640_, _02638_);
  and (_02642_, _02641_, _01598_);
  and (_02643_, _02138_, _01710_);
  and (_02644_, _02132_, _01710_);
  or (_02645_, _02644_, _01765_);
  or (_02646_, _02645_, _02643_);
  nor (_02647_, _02646_, _02642_);
  and (_02648_, _02647_, _02637_);
  and (_02649_, _02306_, _00334_);
  and (_02650_, _02294_, _00380_);
  nor (_02651_, _02650_, _02649_);
  and (_02652_, _02290_, _00338_);
  and (_02653_, _02270_, _00350_);
  nor (_02654_, _02653_, _02652_);
  and (_02655_, _02654_, _02651_);
  and (_02656_, _02312_, _00359_);
  and (_02657_, _02317_, _00363_);
  nor (_02658_, _02657_, _02656_);
  and (_02659_, _02308_, _00376_);
  and (_02660_, _02281_, _00383_);
  nor (_02661_, _02660_, _02659_);
  and (_02662_, _02661_, _02658_);
  and (_02663_, _02662_, _02655_);
  and (_02664_, _02319_, _00356_);
  and (_02665_, _02301_, _00344_);
  nor (_02666_, _02665_, _02664_);
  and (_02667_, _02303_, _00336_);
  and (_02668_, _02286_, _00340_);
  nor (_02669_, _02668_, _02667_);
  and (_02670_, _02669_, _02666_);
  and (_02671_, _02277_, _00374_);
  and (_02672_, _02296_, _00369_);
  nor (_02673_, _02672_, _02671_);
  and (_02674_, _02314_, _00346_);
  and (_02675_, _02273_, _00348_);
  nor (_02676_, _02675_, _02674_);
  and (_02677_, _02676_, _02673_);
  and (_02678_, _02677_, _02670_);
  and (_02679_, _02678_, _02663_);
  nor (_02680_, _02679_, _02037_);
  or (_02681_, _02680_, _02648_);
  and (_02682_, _02124_, _01984_);
  and (_02683_, _02030_, _01717_);
  and (_02684_, _02683_, _01598_);
  or (_02685_, _02684_, _02123_);
  nor (_02686_, _02685_, _02682_);
  and (_02687_, _02686_, _02681_);
  not (_02688_, _02123_);
  nor (_02689_, _02688_, _01984_);
  or (_02690_, _02689_, _02687_);
  and (_02691_, _02570_, _01721_);
  not (_02692_, _02691_);
  and (_02693_, _02138_, _01721_);
  not (_02694_, _02693_);
  and (_02695_, _02219_, _01721_);
  and (_02696_, _02222_, _01721_);
  nor (_02697_, _02696_, _02695_);
  and (_02698_, _02697_, _02694_);
  and (_02699_, _02698_, _02692_);
  and (_02700_, _02699_, _02690_);
  nor (_02701_, _02333_, _02028_);
  and (_02702_, _02132_, _01727_);
  not (_02703_, _02702_);
  and (_02704_, _02222_, _01727_);
  not (_02705_, _02704_);
  and (_02706_, _02599_, _01727_);
  and (_02707_, _02137_, _01598_);
  and (_02708_, _02707_, _01727_);
  nor (_02709_, _02708_, _02706_);
  and (_02710_, _02709_, _02705_);
  and (_02711_, _02710_, _02703_);
  not (_02712_, _02711_);
  nor (_02713_, _02712_, _02701_);
  nor (_02714_, _02344_, _02028_);
  or (_02715_, _02599_, _02707_);
  and (_02716_, _02715_, _01735_);
  not (_02717_, _02716_);
  and (_02718_, _02222_, _01735_);
  and (_02719_, _02132_, _01735_);
  nor (_02720_, _02719_, _02718_);
  and (_02721_, _02720_, _02717_);
  not (_02722_, _02721_);
  nor (_02723_, _02722_, _02714_);
  and (_02724_, _02723_, _02713_);
  and (_02725_, _02724_, _02700_);
  nor (_02726_, _02338_, _02028_);
  and (_02727_, _02707_, _01725_);
  not (_02728_, _01598_);
  not (_02729_, _01725_);
  nor (_02730_, _02030_, _02132_);
  or (_02731_, _02730_, _02729_);
  nor (_02732_, _02731_, _02728_);
  and (_02733_, _02599_, _01725_);
  or (_02734_, _02733_, _02732_);
  or (_02735_, _02734_, _02345_);
  nor (_02736_, _02735_, _02727_);
  not (_02737_, _02736_);
  nor (_02738_, _02737_, _02726_);
  and (_02739_, _02738_, _02725_);
  nor (_02740_, _02346_, _02027_);
  nor (_02741_, _02740_, _02739_);
  and (_02742_, _02350_, _01986_);
  nor (_02743_, _02742_, _02741_);
  and (_02744_, _02200_, _01984_);
  and (_02745_, _02599_, _01737_);
  not (_02746_, _02745_);
  and (_02747_, _02132_, _01737_);
  and (_02748_, _02222_, _01737_);
  nor (_02749_, _02748_, _02747_);
  and (_02750_, _02749_, _02746_);
  and (_02751_, _02219_, _01737_);
  not (_02752_, _02751_);
  and (_02753_, _02138_, _01737_);
  nor (_02754_, _02753_, _02085_);
  and (_02755_, _02754_, _02752_);
  and (_02756_, _02755_, _02750_);
  not (_02757_, _02756_);
  nor (_02758_, _02757_, _02744_);
  and (_02759_, _02758_, _02743_);
  nor (_02760_, _02087_, _02027_);
  nor (_02761_, _02760_, _02759_);
  and (_02762_, _02083_, _01986_);
  nor (_02763_, _02762_, _02761_);
  and (_02764_, _02243_, _01984_);
  and (_02765_, _02570_, _01566_);
  nor (_02766_, _02765_, _02366_);
  and (_02767_, _02138_, _01566_);
  and (_02768_, _02219_, _01566_);
  and (_02769_, _02222_, _01566_);
  or (_02770_, _02769_, _02768_);
  nor (_02771_, _02770_, _02767_);
  and (_02772_, _02771_, _02766_);
  not (_02774_, _02772_);
  nor (_02775_, _02774_, _02764_);
  and (_02776_, _02775_, _02763_);
  not (_02778_, _02366_);
  nor (_02779_, _02778_, _02027_);
  or (_02780_, _02779_, _02776_);
  and (_02781_, _02780_, _01698_);
  or (_02782_, _02781_, _01985_);
  and (_02783_, _02527_, _01598_);
  not (_02784_, _02783_);
  and (_02785_, _02030_, _01731_);
  and (_02786_, _02785_, _01598_);
  not (_02787_, _02786_);
  and (_02788_, _02570_, _01731_);
  nor (_02789_, _02788_, _02081_);
  and (_02790_, _02789_, _02787_);
  and (_02791_, _02790_, _02784_);
  nand (_02792_, _02791_, _02782_);
  nand (_02793_, _02792_, _02545_);
  or (_02794_, _02793_, _02543_);
  nor (_02795_, _01896_, _39389_);
  nor (_02796_, _01945_, _39225_);
  nor (_02797_, _02796_, _02795_);
  nor (_02798_, _01929_, _38965_);
  nor (_02799_, _01924_, _38923_);
  nor (_02800_, _02799_, _02798_);
  and (_02801_, _02800_, _02797_);
  nor (_02802_, _01915_, _39348_);
  nor (_02803_, _01917_, _39307_);
  nor (_02804_, _02803_, _02802_);
  nor (_02805_, _01907_, _39184_);
  nor (_02806_, _01902_, _39143_);
  nor (_02807_, _02806_, _02805_);
  and (_02808_, _02807_, _02804_);
  and (_02809_, _02808_, _02801_);
  nor (_02810_, _01934_, _38882_);
  nor (_02811_, _01931_, _38841_);
  nor (_02812_, _02811_, _02810_);
  nor (_02813_, _01921_, _39061_);
  nor (_02814_, _01936_, _38632_);
  nor (_02815_, _02814_, _02813_);
  and (_02816_, _02815_, _02812_);
  nor (_02817_, _01940_, _39266_);
  nor (_02818_, _01947_, _39102_);
  nor (_02819_, _02818_, _02817_);
  nor (_02820_, _01942_, _39010_);
  nor (_02821_, _01911_, _38737_);
  nor (_02822_, _02821_, _02820_);
  and (_02823_, _02822_, _02819_);
  and (_02824_, _02823_, _02816_);
  and (_02825_, _02824_, _02809_);
  nor (_02826_, _02825_, _01952_);
  and (_02827_, _02826_, _02419_);
  not (_02828_, _02827_);
  nor (_02829_, _01896_, _39374_);
  nor (_02830_, _01947_, _39087_);
  nor (_02831_, _02830_, _02829_);
  nor (_02832_, _01945_, _39210_);
  nor (_02833_, _01934_, _38867_);
  nor (_02834_, _02833_, _02832_);
  and (_02835_, _02834_, _02831_);
  nor (_02836_, _01921_, _39046_);
  nor (_02837_, _01924_, _38908_);
  nor (_02838_, _02837_, _02836_);
  nor (_02839_, _01917_, _39292_);
  nor (_02840_, _01940_, _39251_);
  nor (_02841_, _02840_, _02839_);
  and (_02842_, _02841_, _02838_);
  and (_02843_, _02842_, _02835_);
  nor (_02844_, _01929_, _38950_);
  nor (_02845_, _01931_, _38826_);
  nor (_02846_, _02845_, _02844_);
  nor (_02847_, _01936_, _38617_);
  nor (_02848_, _01911_, _38690_);
  nor (_02849_, _02848_, _02847_);
  and (_02850_, _02849_, _02846_);
  nor (_02851_, _01902_, _39128_);
  nor (_02852_, _01907_, _39169_);
  nor (_02853_, _02852_, _02851_);
  nor (_02854_, _01915_, _39333_);
  nor (_02855_, _01942_, _38992_);
  nor (_02856_, _02855_, _02854_);
  and (_02857_, _02856_, _02853_);
  and (_02858_, _02857_, _02850_);
  and (_02859_, _02858_, _02843_);
  not (_02860_, _02859_);
  and (_02861_, _02860_, _02461_);
  not (_02862_, _02861_);
  and (_02863_, _02314_, _00432_);
  and (_02864_, _02273_, _00435_);
  nor (_02865_, _02864_, _02863_);
  and (_02866_, _02277_, _00425_);
  and (_02867_, _02301_, _00429_);
  nor (_02868_, _02867_, _02866_);
  and (_02869_, _02868_, _02865_);
  and (_02870_, _02294_, _00397_);
  and (_02871_, _02317_, _00411_);
  nor (_02872_, _02871_, _02870_);
  and (_02873_, _02303_, _00389_);
  and (_02874_, _02286_, _00391_);
  nor (_02875_, _02874_, _02873_);
  and (_02876_, _02875_, _02872_);
  and (_02877_, _02876_, _02869_);
  and (_02878_, _02306_, _00401_);
  and (_02879_, _02308_, _00399_);
  nor (_02880_, _02879_, _02878_);
  and (_02881_, _02281_, _00406_);
  and (_02882_, _02296_, _00408_);
  nor (_02883_, _02882_, _02881_);
  and (_02884_, _02883_, _02880_);
  and (_02885_, _02312_, _00415_);
  and (_02886_, _02270_, _00437_);
  nor (_02887_, _02886_, _02885_);
  and (_02888_, _02319_, _00423_);
  and (_02889_, _02290_, _00393_);
  nor (_02890_, _02889_, _02888_);
  and (_02891_, _02890_, _02887_);
  and (_02892_, _02891_, _02884_);
  and (_02893_, _02892_, _02877_);
  nor (_02894_, _02893_, _02037_);
  and (_02895_, _02512_, _01727_);
  and (_02896_, _01714_, _01497_);
  and (_02897_, _02896_, _02512_);
  nor (_02898_, _02897_, _02895_);
  and (_02899_, _02130_, _01766_);
  nor (_02900_, _02638_, _02899_);
  and (_02901_, _02900_, _02898_);
  and (_02902_, _02130_, _01721_);
  nor (_02903_, _02902_, _02580_);
  and (_02904_, _02130_, _01727_);
  and (_02905_, _02130_, _01735_);
  nor (_02906_, _02905_, _02904_);
  and (_02907_, _02906_, _02903_);
  and (_02908_, _02907_, _02901_);
  and (_02909_, _02531_, _02504_);
  nor (_02910_, _02909_, _02524_);
  not (_02911_, _02910_);
  and (_02912_, _02130_, _01725_);
  not (_02913_, _02912_);
  and (_02914_, _02130_, _01737_);
  nor (_02915_, _02914_, _02554_);
  and (_02916_, _02915_, _02913_);
  and (_02917_, _02916_, _02911_);
  and (_02918_, _02917_, _02908_);
  and (_02919_, _02083_, \oc8051_golden_model_1.SP [1]);
  nor (_02920_, _02919_, _02565_);
  and (_02921_, _02350_, \oc8051_golden_model_1.SP [1]);
  and (_02922_, _02155_, \oc8051_golden_model_1.SP [1]);
  nor (_02923_, _02922_, _02921_);
  and (_02924_, _02923_, _02920_);
  and (_02925_, _02130_, _01731_);
  and (_02926_, _02130_, _02056_);
  nor (_02927_, _02926_, _02925_);
  nor (_02928_, _02513_, _02227_);
  and (_02929_, _02928_, _02927_);
  and (_02930_, _02130_, _01566_);
  nor (_02931_, _02930_, _02639_);
  and (_02932_, _02931_, _02526_);
  and (_02933_, _02932_, _02929_);
  and (_02934_, _02933_, _02924_);
  and (_02935_, _02934_, _02918_);
  not (_02936_, _02935_);
  nor (_02937_, _02936_, _02894_);
  and (_02938_, _02937_, _02862_);
  and (_02939_, _02938_, _02828_);
  not (_02940_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_02941_, _02792_, _02545_);
  or (_02942_, _02941_, _02940_);
  and (_02943_, _02942_, _02939_);
  nand (_02944_, _02943_, _02794_);
  not (_02945_, \oc8051_golden_model_1.IRAM[3] [0]);
  or (_02946_, _02941_, _02945_);
  not (_02947_, _02939_);
  not (_02948_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_02949_, _02793_, _02948_);
  and (_02950_, _02949_, _02947_);
  nand (_02951_, _02950_, _02946_);
  nand (_02952_, _02951_, _02944_);
  nand (_02953_, _02952_, _02542_);
  not (_02954_, _02542_);
  not (_02955_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_02956_, _02941_, _02955_);
  not (_02957_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_02958_, _02793_, _02957_);
  and (_02959_, _02958_, _02947_);
  nand (_02960_, _02959_, _02956_);
  not (_02961_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_02962_, _02793_, _02961_);
  not (_02963_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_02964_, _02941_, _02963_);
  and (_02965_, _02964_, _02939_);
  nand (_02966_, _02965_, _02962_);
  nand (_02967_, _02966_, _02960_);
  nand (_02968_, _02967_, _02954_);
  nand (_02969_, _02968_, _02953_);
  nand (_02970_, _02969_, _02379_);
  not (_02971_, _02379_);
  not (_02972_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_02973_, _02941_, _02972_);
  not (_02974_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_02975_, _02793_, _02974_);
  and (_02976_, _02975_, _02947_);
  nand (_02977_, _02976_, _02973_);
  not (_02978_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_02979_, _02793_, _02978_);
  not (_02980_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_02981_, _02941_, _02980_);
  and (_02982_, _02981_, _02939_);
  nand (_02983_, _02982_, _02979_);
  nand (_02984_, _02983_, _02977_);
  nand (_02985_, _02984_, _02542_);
  not (_02986_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_02987_, _02941_, _02986_);
  not (_02988_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_02989_, _02793_, _02988_);
  and (_02990_, _02989_, _02947_);
  nand (_02991_, _02990_, _02987_);
  not (_02992_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_02993_, _02793_, _02992_);
  not (_02994_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_02995_, _02941_, _02994_);
  and (_02996_, _02995_, _02939_);
  nand (_02997_, _02996_, _02993_);
  nand (_02998_, _02997_, _02991_);
  nand (_02999_, _02998_, _02954_);
  nand (_03000_, _02999_, _02985_);
  nand (_03001_, _03000_, _02971_);
  and (_03002_, _03001_, _02970_);
  nor (_03003_, _03002_, _02080_);
  nor (_03004_, _03003_, _02077_);
  nor (_03005_, _02058_, _01952_);
  not (_03006_, _02158_);
  nor (_03007_, _03006_, _01952_);
  and (_03008_, _03007_, _02027_);
  nor (_03009_, _03008_, _03005_);
  and (_03010_, _03009_, _03004_);
  not (_03011_, _03010_);
  and (_03012_, _03011_, _02059_);
  nor (_03013_, _01745_, _01986_);
  nor (_03014_, _03013_, _03012_);
  nor (_03015_, _02519_, _01952_);
  and (_03016_, _03015_, _02027_);
  and (_03017_, _02067_, _02051_);
  nor (_03018_, _03017_, _03016_);
  and (_03019_, _03018_, _03014_);
  nand (_03020_, _03001_, _02970_);
  and (_03021_, _03020_, _02582_);
  not (_03022_, _03021_);
  and (_03023_, _03022_, _03019_);
  nor (_03024_, _02054_, _01952_);
  nor (_03025_, _02549_, _01952_);
  and (_03026_, _03025_, _02027_);
  nor (_03027_, _03026_, _03024_);
  and (_03028_, _03027_, _03023_);
  nor (_03029_, _03028_, _02055_);
  nor (_03030_, _03029_, _02052_);
  and (_03031_, _02052_, _01986_);
  or (_03032_, _03031_, _03030_);
  and (_03033_, _03032_, _02050_);
  nor (_03034_, _03033_, _02048_);
  nor (_03035_, _01750_, _01986_);
  and (_03036_, _02067_, _02128_);
  nor (_03037_, _03036_, _03035_);
  not (_03038_, _03037_);
  nor (_03039_, _03038_, _03034_);
  nor (_03040_, _02043_, _01952_);
  and (_03041_, _02030_, _02128_);
  and (_03042_, _03020_, _03041_);
  nor (_03043_, _03042_, _03040_);
  and (_03044_, _03043_, _03039_);
  nor (_03045_, _03044_, _02044_);
  nor (_03046_, _03045_, _01767_);
  and (_03047_, _01767_, _01986_);
  nor (_03048_, _03047_, _03046_);
  and (_03049_, _02067_, _01717_);
  or (_03050_, _03049_, _03048_);
  nor (_03051_, _03050_, _02041_);
  and (_03052_, _03020_, _02683_);
  nor (_03053_, _03052_, _01996_);
  and (_03054_, _03053_, _03051_);
  nor (_03055_, _03054_, _02029_);
  nor (_03056_, _03055_, _01718_);
  and (_03057_, _01718_, _01986_);
  nor (_03058_, _03057_, _03056_);
  not (_03059_, _02210_);
  nor (_03060_, _03059_, _01952_);
  not (_03061_, _02331_);
  nor (_03062_, _03061_, _01952_);
  nor (_03063_, _03062_, _03060_);
  nor (_03064_, _02208_, _01952_);
  not (_03065_, _02342_);
  nor (_03066_, _03065_, _01952_);
  nor (_03067_, _03066_, _03064_);
  and (_03068_, _03067_, _03063_);
  nor (_03069_, _03068_, _02028_);
  nor (_03070_, _03069_, _01728_);
  not (_03071_, _03070_);
  nor (_03072_, _03071_, _03058_);
  and (_03073_, _01728_, _01986_);
  nor (_03074_, _03073_, _03072_);
  nor (_03075_, _02335_, _01952_);
  and (_03076_, _03075_, _02027_);
  nor (_03077_, _03076_, _01726_);
  not (_03078_, _03077_);
  nor (_03079_, _03078_, _03074_);
  nor (_03080_, _03079_, _01993_);
  and (_03081_, _02067_, _01566_);
  nor (_03082_, _03081_, _03080_);
  nor (_03083_, _02778_, _01952_);
  and (_03084_, _02030_, _01566_);
  and (_03085_, _03020_, _03084_);
  nor (_03086_, _03085_, _03083_);
  and (_03087_, _03086_, _03082_);
  and (_03088_, _03083_, _02028_);
  nor (_03089_, _03088_, _03087_);
  or (_03090_, _03089_, _01992_);
  nor (_03091_, _03090_, _01991_);
  nor (_03092_, _03091_, _01985_);
  and (_03093_, _02067_, _01731_);
  nor (_03094_, _03093_, _03092_);
  and (_03095_, _03020_, _02785_);
  not (_03096_, _03095_);
  and (_03097_, _03096_, _03094_);
  nor (_03098_, _02082_, _01952_);
  and (_03099_, _03098_, _02027_);
  not (_03100_, _03099_);
  and (_03101_, _03100_, _03097_);
  and (_03102_, _03098_, _02860_);
  and (_03103_, _02826_, _01697_);
  not (_03104_, \oc8051_golden_model_1.SP [1]);
  and (_03105_, _03104_, \oc8051_golden_model_1.SP [0]);
  and (_03106_, \oc8051_golden_model_1.SP [1], _01986_);
  nor (_03107_, _03106_, _03105_);
  not (_03108_, _03107_);
  nor (_03109_, _03108_, _01990_);
  and (_03110_, _03108_, _01726_);
  and (_03111_, _02860_, _01996_);
  and (_03112_, _02826_, _02042_);
  and (_03113_, _03108_, _02052_);
  not (_03114_, _02052_);
  nand (_03115_, _02941_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand (_03116_, _02793_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_03117_, _03116_, _02939_);
  nand (_03118_, _03117_, _03115_);
  nand (_03119_, _02793_, \oc8051_golden_model_1.IRAM[3] [1]);
  nand (_03120_, _02941_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_03121_, _03120_, _02947_);
  nand (_03122_, _03121_, _03119_);
  nand (_03123_, _03122_, _03118_);
  nand (_03124_, _03123_, _02542_);
  nand (_03125_, _02793_, \oc8051_golden_model_1.IRAM[7] [1]);
  nand (_03126_, _02941_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_03127_, _03126_, _02947_);
  nand (_03128_, _03127_, _03125_);
  nand (_03129_, _02941_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand (_03130_, _02793_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_03131_, _03130_, _02939_);
  nand (_03132_, _03131_, _03129_);
  nand (_03133_, _03132_, _03128_);
  nand (_03134_, _03133_, _02954_);
  nand (_03135_, _03134_, _03124_);
  nand (_03136_, _03135_, _02379_);
  nand (_03137_, _02793_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_03138_, _02941_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03139_, _03138_, _02947_);
  nand (_03140_, _03139_, _03137_);
  nand (_03141_, _02941_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_03142_, _02793_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03143_, _03142_, _02939_);
  nand (_03144_, _03143_, _03141_);
  nand (_03145_, _03144_, _03140_);
  nand (_03146_, _03145_, _02542_);
  nand (_03147_, _02793_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_03148_, _02941_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_03149_, _03148_, _02947_);
  nand (_03150_, _03149_, _03147_);
  nand (_03151_, _02941_, \oc8051_golden_model_1.IRAM[12] [1]);
  not (_03152_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_03153_, _02941_, _03152_);
  and (_03154_, _03153_, _02939_);
  nand (_03156_, _03154_, _03151_);
  nand (_03157_, _03156_, _03150_);
  nand (_03158_, _03157_, _02954_);
  nand (_03159_, _03158_, _03146_);
  nand (_03160_, _03159_, _02971_);
  nand (_03161_, _03160_, _03136_);
  not (_03163_, _03161_);
  or (_03164_, _03163_, _02080_);
  not (_03165_, _03007_);
  and (_03167_, _02496_, _02061_);
  nor (_03168_, _03167_, _02064_);
  and (_03170_, _02860_, _02064_);
  or (_03171_, _03170_, _02060_);
  or (_03173_, _03171_, _03168_);
  and (_03174_, _02132_, _02056_);
  and (_03176_, _02133_, _02056_);
  nor (_03177_, _03176_, _03174_);
  nor (_03178_, _03108_, _01747_);
  and (_03180_, _02497_, _02056_);
  nor (_03181_, _03180_, _03178_);
  and (_03183_, _03181_, _03177_);
  and (_03184_, _03183_, _03173_);
  and (_03186_, _03184_, _03165_);
  and (_03187_, _03186_, _03164_);
  and (_03189_, _03007_, _02860_);
  nor (_03190_, _03189_, _03187_);
  and (_03191_, _02825_, _03005_);
  nor (_03192_, _03191_, _03190_);
  or (_03194_, _03108_, _01745_);
  nand (_03195_, _03194_, _03192_);
  and (_03197_, _03015_, _02859_);
  and (_03198_, _02496_, _02051_);
  nor (_03200_, _03198_, _03197_);
  not (_03201_, _03200_);
  nor (_03203_, _03201_, _03195_);
  and (_03205_, _03161_, _02582_);
  nor (_03207_, _03205_, _03025_);
  and (_03208_, _03207_, _03203_);
  and (_03210_, _03025_, _02860_);
  nor (_03211_, _03210_, _03208_);
  and (_03213_, _02825_, _03024_);
  nor (_03215_, _03213_, _03211_);
  and (_03216_, _03215_, _03114_);
  nor (_03218_, _03216_, _03113_);
  and (_03219_, _02049_, _02825_);
  or (_03221_, _03219_, _03218_);
  not (_03222_, _02135_);
  nor (_03224_, _03108_, _01750_);
  not (_03225_, _03224_);
  and (_03227_, _02247_, _02128_);
  nor (_03229_, _03227_, _02139_);
  and (_03231_, _03229_, _03225_);
  and (_03233_, _03231_, _03222_);
  not (_03235_, _03233_);
  nor (_03237_, _03235_, _03221_);
  and (_03239_, _03161_, _03041_);
  nor (_03241_, _03239_, _03040_);
  and (_03243_, _03241_, _03237_);
  nor (_03245_, _03243_, _03112_);
  nor (_03247_, _03245_, _01767_);
  and (_03248_, _03108_, _01767_);
  nor (_03249_, _03248_, _03247_);
  nor (_03250_, _02040_, _02860_);
  and (_03251_, _02496_, _01717_);
  nor (_03252_, _03251_, _03250_);
  not (_03253_, _03252_);
  nor (_03254_, _03253_, _03249_);
  and (_03255_, _03161_, _02683_);
  nor (_03256_, _03255_, _01996_);
  and (_03257_, _03256_, _03254_);
  nor (_03258_, _03257_, _03111_);
  nor (_03259_, _03258_, _01718_);
  and (_03260_, _03108_, _01718_);
  nor (_03261_, _03260_, _03259_);
  nor (_03262_, _03068_, _02860_);
  nor (_03263_, _03262_, _01728_);
  not (_03264_, _03263_);
  nor (_03265_, _03264_, _03261_);
  and (_03266_, _03108_, _01728_);
  nor (_03267_, _03266_, _03265_);
  and (_03268_, _03075_, _02859_);
  nor (_03269_, _03268_, _01726_);
  not (_03270_, _03269_);
  nor (_03271_, _03270_, _03267_);
  nor (_03272_, _03271_, _03110_);
  and (_03273_, _02132_, _01566_);
  and (_03274_, _02133_, _01566_);
  nor (_03275_, _03274_, _03273_);
  and (_03276_, _02497_, _01566_);
  not (_03277_, _03276_);
  and (_03278_, _03277_, _03275_);
  not (_03279_, _03278_);
  nor (_03280_, _03279_, _03272_);
  and (_03281_, _03161_, _03084_);
  nor (_03282_, _03281_, _03083_);
  and (_03283_, _03282_, _03280_);
  and (_03284_, _03083_, _02860_);
  nor (_03285_, _03284_, _03283_);
  or (_03286_, _03285_, _01992_);
  nor (_03287_, _03286_, _03109_);
  nor (_03288_, _03287_, _03103_);
  and (_03289_, _02497_, _01731_);
  and (_03290_, _02132_, _01731_);
  and (_03291_, _02133_, _01731_);
  nor (_03292_, _03291_, _03290_);
  not (_03293_, _03292_);
  nor (_03294_, _03293_, _03289_);
  not (_03295_, _03294_);
  nor (_03296_, _03295_, _03288_);
  and (_03297_, _03161_, _02785_);
  nor (_03298_, _03297_, _03098_);
  and (_03299_, _03298_, _03296_);
  nor (_03300_, _03299_, _03102_);
  not (_03301_, _01764_);
  and (_03302_, _02134_, _03301_);
  not (_03303_, _03302_);
  and (_03304_, _03303_, _02034_);
  not (_03305_, _03304_);
  and (_03306_, _02034_, _02137_);
  not (_03307_, _03306_);
  not (_03308_, _01718_);
  and (_03309_, _01748_, _03308_);
  not (_03310_, _01750_);
  nor (_03311_, _01767_, _03310_);
  and (_03312_, _03311_, _01729_);
  and (_03313_, _03312_, _03309_);
  or (_03314_, _02133_, _02130_);
  and (_03315_, _03314_, _02051_);
  and (_03316_, _03314_, _02128_);
  nor (_03317_, _03316_, _03315_);
  and (_03318_, _02129_, _02061_);
  nor (_03319_, _03318_, _02527_);
  and (_03320_, _03319_, _03317_);
  and (_03321_, _01990_, _02787_);
  and (_03322_, _03321_, _03320_);
  and (_03323_, _03322_, _03313_);
  and (_03324_, _02236_, _01731_);
  not (_03325_, _03324_);
  and (_03326_, _03292_, _03325_);
  nor (_03327_, _02132_, _02138_);
  and (_03328_, _03327_, _02141_);
  nor (_03329_, _03328_, _01754_);
  not (_03330_, _03329_);
  and (_03331_, _03330_, _03326_);
  and (_03332_, _03331_, _03323_);
  not (_03333_, _01717_);
  nor (_03334_, _03327_, _03333_);
  not (_03335_, _03334_);
  not (_03336_, _02590_);
  nor (_03337_, _02511_, _02052_);
  and (_03338_, _03337_, _03336_);
  and (_03339_, _03338_, _03335_);
  and (_03340_, _03275_, _03177_);
  and (_03341_, _03340_, _03339_);
  nor (_03342_, _03276_, _02930_);
  and (_03343_, _03342_, _02080_);
  nor (_03344_, _02141_, _03333_);
  nor (_03345_, _03344_, _03084_);
  nor (_03346_, _02140_, _01746_);
  nor (_03347_, _03346_, _02683_);
  and (_03348_, _03347_, _03345_);
  and (_03349_, _03348_, _03343_);
  and (_03350_, _02512_, _01566_);
  nor (_03351_, _03041_, _03350_);
  and (_03352_, _03314_, _01717_);
  nor (_03353_, _03352_, _02528_);
  and (_03354_, _03353_, _03351_);
  nor (_03355_, _02926_, _02582_);
  nor (_03356_, _02925_, _02581_);
  and (_03357_, _03356_, _03355_);
  and (_03358_, _03357_, _03354_);
  and (_03359_, _03358_, _03349_);
  and (_03360_, _03359_, _03341_);
  and (_03361_, _03360_, _03332_);
  not (_03362_, _03361_);
  nor (_03363_, _03362_, _01996_);
  and (_03364_, _03363_, _03307_);
  and (_03365_, _03364_, _03305_);
  nor (_03366_, _02049_, _03007_);
  nor (_03367_, _03015_, _02064_);
  and (_03368_, _03367_, _03366_);
  nor (_03369_, _02639_, _02053_);
  nor (_03370_, _02057_, _02042_);
  and (_03371_, _03370_, _03369_);
  nor (_03372_, _03371_, _01952_);
  nor (_03373_, _03372_, _03025_);
  nor (_03374_, _03083_, _02033_);
  and (_03375_, _03374_, _03373_);
  and (_03376_, _03375_, _03368_);
  not (_03377_, _01992_);
  nor (_03378_, _03098_, _03075_);
  and (_03379_, _03378_, _03377_);
  and (_03380_, _03379_, _03068_);
  and (_03381_, _03380_, _03376_);
  and (_03382_, _03381_, _03365_);
  and (_00001_, _39632_, _39026_);
  not (_03383_, _00001_);
  nor (_03384_, _03383_, _03382_);
  not (_03385_, _03384_);
  nor (_03386_, _03385_, _03300_);
  and (_03387_, _03386_, _03101_);
  not (_03388_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_03389_, _02793_, _03388_);
  nand (_03390_, _02793_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_03391_, _03390_, _02939_);
  nand (_03392_, _03391_, _03389_);
  nand (_03393_, _02793_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand (_03394_, _02941_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_03395_, _03394_, _02947_);
  nand (_03396_, _03395_, _03393_);
  nand (_03397_, _03396_, _03392_);
  nand (_03398_, _03397_, _02542_);
  nand (_03399_, _02793_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand (_03400_, _02941_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_03401_, _03400_, _02947_);
  nand (_03402_, _03401_, _03399_);
  nand (_03403_, _02941_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand (_03404_, _02793_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_03405_, _03404_, _02939_);
  nand (_03406_, _03405_, _03403_);
  nand (_03407_, _03406_, _03402_);
  nand (_03408_, _03407_, _02954_);
  nand (_03409_, _03408_, _03398_);
  nand (_03410_, _03409_, _02379_);
  nand (_03411_, _02793_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_03412_, _02941_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_03413_, _03412_, _02947_);
  nand (_03414_, _03413_, _03411_);
  nand (_03415_, _02941_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_03416_, _02793_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_03417_, _03416_, _02939_);
  nand (_03418_, _03417_, _03415_);
  nand (_03419_, _03418_, _03414_);
  nand (_03420_, _03419_, _02542_);
  nand (_03421_, _02793_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_03422_, _02941_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_03423_, _03422_, _02947_);
  nand (_03424_, _03423_, _03421_);
  nand (_03425_, _02941_, \oc8051_golden_model_1.IRAM[12] [3]);
  not (_03426_, \oc8051_golden_model_1.IRAM[13] [3]);
  or (_03427_, _02941_, _03426_);
  and (_03428_, _03427_, _02939_);
  nand (_03429_, _03428_, _03425_);
  nand (_03430_, _03429_, _03424_);
  nand (_03431_, _03430_, _02954_);
  nand (_03432_, _03431_, _03420_);
  nand (_03433_, _03432_, _02971_);
  nand (_03434_, _03433_, _03410_);
  and (_03435_, _03434_, _02683_);
  and (_03436_, _03434_, _03041_);
  and (_03437_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_03438_, _03437_, \oc8051_golden_model_1.SP [2]);
  nor (_03439_, _03438_, \oc8051_golden_model_1.SP [3]);
  and (_03440_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_03441_, _03440_, \oc8051_golden_model_1.SP [3]);
  and (_03442_, _03441_, \oc8051_golden_model_1.SP [0]);
  nor (_03443_, _03442_, _03439_);
  not (_03444_, _03443_);
  nor (_03445_, _03444_, _01750_);
  not (_03446_, _01745_);
  and (_03447_, _03005_, _02118_);
  and (_03448_, _03434_, _02079_);
  nor (_03449_, _03444_, _01747_);
  nor (_03450_, _02078_, \oc8051_golden_model_1.PSW [3]);
  and (_03451_, _03434_, _02078_);
  nor (_03452_, _03451_, _03450_);
  nor (_03453_, _03452_, _02064_);
  and (_03454_, _02064_, _01983_);
  nor (_03455_, _03454_, _02060_);
  not (_03456_, _03455_);
  nor (_03457_, _03456_, _03453_);
  or (_03458_, _03457_, _02079_);
  nor (_03459_, _03458_, _03449_);
  or (_03460_, _03459_, _03007_);
  nor (_03461_, _03460_, _03448_);
  and (_03462_, _03007_, _02120_);
  or (_03463_, _03462_, _03005_);
  nor (_03464_, _03463_, _03461_);
  nor (_03465_, _03464_, _03447_);
  nor (_03466_, _03465_, _03446_);
  nor (_03467_, _03443_, _01745_);
  nor (_03468_, _03467_, _03015_);
  not (_03469_, _03468_);
  nor (_03470_, _03469_, _03466_);
  and (_03471_, _03015_, _02120_);
  nor (_03472_, _03471_, _02582_);
  not (_03473_, _03472_);
  nor (_03474_, _03473_, _03470_);
  and (_03475_, _03434_, _02582_);
  nor (_03476_, _03475_, _03025_);
  not (_03477_, _03476_);
  nor (_03478_, _03477_, _03474_);
  and (_03479_, _03025_, _02120_);
  or (_03480_, _03479_, _03024_);
  nor (_03481_, _03480_, _03478_);
  and (_03482_, _02118_, _03024_);
  nor (_03483_, _03482_, _03481_);
  and (_03484_, _03483_, _03114_);
  and (_03485_, _03443_, _02052_);
  nor (_03486_, _03485_, _03484_);
  nor (_03487_, _03486_, _02049_);
  nor (_03488_, _02050_, _02122_);
  or (_03489_, _03488_, _03487_);
  and (_03490_, _03489_, _01750_);
  or (_03491_, _03490_, _03041_);
  nor (_03492_, _03491_, _03445_);
  or (_03493_, _03492_, _03040_);
  nor (_03494_, _03493_, _03436_);
  not (_03495_, _02118_);
  and (_03496_, _03495_, _03040_);
  nor (_03497_, _03496_, _03494_);
  nor (_03498_, _03497_, _01767_);
  and (_03499_, _03443_, _01767_);
  not (_03500_, _03499_);
  and (_03501_, _03500_, _02040_);
  not (_03502_, _03501_);
  nor (_03503_, _03502_, _03498_);
  nor (_03504_, _02040_, _02120_);
  nor (_03505_, _03504_, _03503_);
  nor (_03506_, _03505_, _02683_);
  or (_03507_, _03506_, _01996_);
  nor (_03508_, _03507_, _03435_);
  nor (_03509_, _01995_, _01984_);
  nor (_03510_, _03509_, _03508_);
  nor (_03511_, _03510_, _01718_);
  and (_03512_, _03443_, _01718_);
  not (_03513_, _03512_);
  and (_03514_, _03513_, _03068_);
  not (_03515_, _03514_);
  nor (_03516_, _03515_, _03511_);
  nor (_03517_, _03068_, _02120_);
  nor (_03518_, _03517_, _01728_);
  not (_03519_, _03518_);
  nor (_03520_, _03519_, _03516_);
  and (_03521_, _03443_, _01728_);
  nor (_03522_, _03521_, _03075_);
  not (_03523_, _03522_);
  nor (_03524_, _03523_, _03520_);
  and (_03525_, _03075_, _01983_);
  nor (_03526_, _03525_, _01726_);
  not (_03527_, _03526_);
  nor (_03528_, _03527_, _03524_);
  and (_03529_, _03443_, _01726_);
  nor (_03530_, _03529_, _03084_);
  not (_03531_, _03530_);
  nor (_03532_, _03531_, _03528_);
  and (_03533_, _03434_, _03084_);
  nor (_03534_, _03533_, _03083_);
  not (_03535_, _03534_);
  nor (_03536_, _03535_, _03532_);
  not (_03537_, _01990_);
  and (_03538_, _03083_, _02120_);
  nor (_03539_, _03538_, _03537_);
  not (_03540_, _03539_);
  nor (_03541_, _03540_, _03536_);
  nor (_03542_, _03443_, _01990_);
  nor (_03543_, _03542_, _01992_);
  not (_03544_, _03543_);
  nor (_03545_, _03544_, _03541_);
  and (_03546_, _01992_, _03495_);
  nor (_03547_, _03546_, _02785_);
  not (_03548_, _03547_);
  nor (_03549_, _03548_, _03545_);
  and (_03550_, _03434_, _02785_);
  nor (_03551_, _03550_, _03098_);
  not (_03552_, _03551_);
  nor (_03553_, _03552_, _03549_);
  nor (_03554_, _02082_, _01984_);
  nor (_03555_, _03554_, _03553_);
  and (_03556_, _03098_, _02453_);
  and (_03557_, _02411_, _01697_);
  nor (_03558_, _03437_, \oc8051_golden_model_1.SP [2]);
  nor (_03559_, _03558_, _03438_);
  and (_03560_, _03559_, _01726_);
  and (_03561_, _02453_, _01996_);
  nor (_03562_, _02040_, _02453_);
  and (_03563_, _03559_, _02052_);
  not (_03564_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_03565_, _02793_, _03564_);
  not (_03566_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_03567_, _02941_, _03566_);
  and (_03568_, _03567_, _02939_);
  nand (_03569_, _03568_, _03565_);
  not (_03570_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_03571_, _02941_, _03570_);
  not (_03572_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_03573_, _02793_, _03572_);
  and (_03574_, _03573_, _02947_);
  nand (_03575_, _03574_, _03571_);
  nand (_03576_, _03575_, _03569_);
  nand (_03577_, _03576_, _02542_);
  not (_03578_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_03579_, _02941_, _03578_);
  not (_03580_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_03581_, _02793_, _03580_);
  and (_03582_, _03581_, _02947_);
  nand (_03583_, _03582_, _03579_);
  not (_03584_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_03585_, _02793_, _03584_);
  not (_03586_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_03587_, _02941_, _03586_);
  and (_03588_, _03587_, _02939_);
  nand (_03589_, _03588_, _03585_);
  nand (_03590_, _03589_, _03583_);
  nand (_03591_, _03590_, _02954_);
  nand (_03592_, _03591_, _03577_);
  nand (_03593_, _03592_, _02379_);
  not (_03594_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_03595_, _02941_, _03594_);
  not (_03596_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_03597_, _02793_, _03596_);
  and (_03598_, _03597_, _02947_);
  nand (_03599_, _03598_, _03595_);
  not (_03600_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_03601_, _02793_, _03600_);
  not (_03602_, \oc8051_golden_model_1.IRAM[9] [2]);
  or (_03603_, _02941_, _03602_);
  and (_03604_, _03603_, _02939_);
  nand (_03605_, _03604_, _03601_);
  nand (_03606_, _03605_, _03599_);
  nand (_03607_, _03606_, _02542_);
  not (_03608_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_03609_, _02941_, _03608_);
  not (_03610_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_03611_, _02793_, _03610_);
  and (_03612_, _03611_, _02947_);
  nand (_03613_, _03612_, _03609_);
  not (_03614_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_03615_, _02793_, _03614_);
  not (_03616_, \oc8051_golden_model_1.IRAM[13] [2]);
  or (_03617_, _02941_, _03616_);
  and (_03618_, _03617_, _02939_);
  nand (_03619_, _03618_, _03615_);
  nand (_03620_, _03619_, _03613_);
  nand (_03621_, _03620_, _02954_);
  nand (_03622_, _03621_, _03607_);
  nand (_03623_, _03622_, _02971_);
  nand (_03624_, _03623_, _03593_);
  not (_03625_, _03624_);
  or (_03626_, _03625_, _02080_);
  nor (_03628_, _03318_, _02064_);
  and (_03630_, _02453_, _02064_);
  or (_03632_, _03630_, _02060_);
  or (_03634_, _03632_, _03628_);
  nor (_03636_, _03559_, _01747_);
  nor (_03638_, _03636_, _02926_);
  and (_03640_, _03638_, _03177_);
  and (_03642_, _03640_, _03634_);
  and (_03644_, _03642_, _03165_);
  and (_03646_, _03644_, _03626_);
  and (_03648_, _03007_, _02453_);
  nor (_03650_, _03648_, _03646_);
  and (_03652_, _03005_, _02410_);
  nor (_03654_, _03652_, _03650_);
  nor (_03656_, _03559_, _01745_);
  nor (_03657_, _03656_, _03015_);
  and (_03658_, _03657_, _03654_);
  and (_03659_, _03015_, _02453_);
  nor (_03660_, _03659_, _03658_);
  and (_03661_, _02129_, _02051_);
  nor (_03662_, _03661_, _03660_);
  and (_03663_, _03624_, _02582_);
  nor (_03664_, _03663_, _03025_);
  and (_03665_, _03664_, _03662_);
  and (_03666_, _03025_, _02453_);
  nor (_03667_, _03666_, _03665_);
  and (_03668_, _02410_, _03024_);
  nor (_03669_, _03668_, _03667_);
  and (_03670_, _03669_, _03114_);
  nor (_03671_, _03670_, _03563_);
  and (_03672_, _02049_, _02410_);
  or (_03673_, _03672_, _03671_);
  nor (_03674_, _03559_, _01750_);
  not (_03675_, _03674_);
  and (_03676_, _03675_, _02136_);
  not (_03677_, _03676_);
  nor (_03678_, _03677_, _03673_);
  and (_03679_, _03624_, _03041_);
  not (_03680_, _03679_);
  and (_03681_, _03680_, _03678_);
  and (_03682_, _02410_, _03040_);
  nor (_03683_, _03682_, _01767_);
  and (_03684_, _03683_, _03681_);
  and (_03685_, _03559_, _01767_);
  nor (_03686_, _03685_, _03684_);
  and (_03688_, _02129_, _01717_);
  or (_03690_, _03688_, _03686_);
  nor (_03692_, _03690_, _03562_);
  and (_03694_, _03624_, _02683_);
  nor (_03696_, _03694_, _01996_);
  and (_03698_, _03696_, _03692_);
  nor (_03700_, _03698_, _03561_);
  nor (_03702_, _03700_, _01718_);
  and (_03704_, _03559_, _01718_);
  nor (_03706_, _03704_, _03702_);
  nor (_03708_, _03068_, _02453_);
  nor (_03710_, _03708_, _01728_);
  not (_03712_, _03710_);
  nor (_03714_, _03712_, _03706_);
  and (_03716_, _03559_, _01728_);
  nor (_03717_, _03716_, _03714_);
  and (_03718_, _03075_, _02452_);
  nor (_03719_, _03718_, _01726_);
  not (_03720_, _03719_);
  nor (_03721_, _03720_, _03717_);
  nor (_03722_, _03721_, _03560_);
  not (_03723_, _02930_);
  and (_03724_, _03275_, _03723_);
  not (_03725_, _03724_);
  nor (_03726_, _03725_, _03722_);
  and (_03727_, _03624_, _03084_);
  nor (_03728_, _03727_, _03083_);
  and (_03729_, _03728_, _03726_);
  and (_03730_, _03083_, _02453_);
  nor (_03731_, _03730_, _03729_);
  nor (_03732_, _03559_, _01990_);
  nor (_03733_, _03732_, _01992_);
  not (_03734_, _03733_);
  nor (_03735_, _03734_, _03731_);
  nor (_03736_, _03735_, _03557_);
  and (_03737_, _02129_, _01731_);
  nor (_03738_, _03737_, _03736_);
  and (_03739_, _03624_, _02785_);
  nor (_03740_, _03739_, _03098_);
  and (_03741_, _03740_, _03738_);
  nor (_03742_, _03741_, _03556_);
  nor (_03743_, _03742_, _03385_);
  not (_03744_, _03743_);
  nor (_03745_, _03744_, _03555_);
  and (_03746_, _03745_, _03387_);
  not (_03747_, _03746_);
  not (_03748_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_03749_, _02793_, _03748_);
  not (_03750_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_03751_, _02941_, _03750_);
  and (_03752_, _03751_, _02939_);
  nand (_03753_, _03752_, _03749_);
  nand (_03754_, _02793_, \oc8051_golden_model_1.IRAM[3] [7]);
  nand (_03755_, _02941_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_03756_, _03755_, _02947_);
  nand (_03757_, _03756_, _03754_);
  nand (_03758_, _03757_, _03753_);
  nand (_03759_, _03758_, _02542_);
  nand (_03760_, _02793_, \oc8051_golden_model_1.IRAM[7] [7]);
  nand (_03761_, _02941_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_03762_, _03761_, _02947_);
  nand (_03763_, _03762_, _03760_);
  nand (_03764_, _02941_, \oc8051_golden_model_1.IRAM[4] [7]);
  nand (_03765_, _02793_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_03766_, _03765_, _02939_);
  nand (_03767_, _03766_, _03764_);
  nand (_03768_, _03767_, _03763_);
  nand (_03769_, _03768_, _02954_);
  nand (_03770_, _03769_, _03759_);
  nand (_03771_, _03770_, _02379_);
  not (_03772_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_03773_, _02941_, _03772_);
  nand (_03774_, _02941_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_03775_, _03774_, _02947_);
  nand (_03776_, _03775_, _03773_);
  nand (_03777_, _02941_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_03778_, _02793_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_03779_, _03778_, _02939_);
  nand (_03780_, _03779_, _03777_);
  nand (_03781_, _03780_, _03776_);
  nand (_03782_, _03781_, _02542_);
  nand (_03783_, _02793_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_03784_, _02941_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_03785_, _03784_, _02947_);
  nand (_03786_, _03785_, _03783_);
  nand (_03787_, _02941_, \oc8051_golden_model_1.IRAM[12] [7]);
  not (_03788_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_03789_, _02941_, _03788_);
  and (_03790_, _03789_, _02939_);
  nand (_03791_, _03790_, _03787_);
  nand (_03792_, _03791_, _03786_);
  nand (_03793_, _03792_, _02954_);
  nand (_03794_, _03793_, _03782_);
  nand (_03795_, _03794_, _02971_);
  nand (_03796_, _03795_, _03771_);
  or (_03797_, _03796_, _01952_);
  and (_03798_, _02118_, _01952_);
  not (_03799_, _02825_);
  and (_03800_, _03799_, _02410_);
  and (_03801_, _03800_, _03798_);
  and (_03802_, _02859_, _02028_);
  and (_03803_, _03802_, _02452_);
  and (_03804_, _03803_, _02120_);
  and (_03805_, _03804_, _03801_);
  and (_03806_, _03805_, \oc8051_golden_model_1.SBUF [7]);
  and (_03807_, _02859_, _02027_);
  and (_03808_, _03807_, _02452_);
  and (_03809_, _03808_, _02120_);
  not (_03810_, _02410_);
  and (_03811_, _02825_, _03810_);
  and (_03812_, _03811_, _03798_);
  and (_03813_, _03812_, _03809_);
  and (_03814_, _03813_, \oc8051_golden_model_1.IE [7]);
  nor (_03815_, _03814_, _03806_);
  and (_03816_, _02452_, _01983_);
  and (_03817_, _03816_, _03807_);
  nor (_03818_, _02825_, _02410_);
  and (_03819_, _03818_, _03798_);
  and (_03820_, _03819_, _03817_);
  and (_03821_, _03820_, \oc8051_golden_model_1.P3 [7]);
  not (_03822_, _03821_);
  and (_03823_, _03798_, _02410_);
  and (_03824_, _03823_, _02825_);
  and (_03825_, _03824_, _01983_);
  nor (_03826_, _02859_, _02027_);
  and (_03827_, _03826_, _02453_);
  and (_03828_, _03827_, _03825_);
  and (_03829_, _03828_, \oc8051_golden_model_1.PCON [7]);
  and (_03830_, _03817_, _03812_);
  and (_03831_, _03830_, \oc8051_golden_model_1.P2 [7]);
  nor (_03832_, _03831_, _03829_);
  and (_03833_, _03832_, _03822_);
  and (_03834_, _03833_, _03815_);
  not (_03835_, _01952_);
  nor (_03836_, _02118_, _03835_);
  and (_03837_, _03836_, _03800_);
  and (_03838_, _03837_, _03817_);
  and (_03839_, _03838_, \oc8051_golden_model_1.PSW [7]);
  and (_03840_, _03836_, _03811_);
  and (_03841_, _03840_, _03817_);
  and (_03842_, _03841_, \oc8051_golden_model_1.ACC [7]);
  nor (_03843_, _03842_, _03839_);
  and (_03844_, _03819_, _03809_);
  and (_03845_, _03844_, \oc8051_golden_model_1.IP [7]);
  and (_03846_, _03818_, _03836_);
  and (_03847_, _03846_, _03817_);
  and (_03848_, _03847_, \oc8051_golden_model_1.B [7]);
  nor (_03849_, _03848_, _03845_);
  and (_03850_, _03849_, _03843_);
  not (_03851_, _03824_);
  nor (_03852_, _02452_, _01983_);
  nand (_03853_, _03852_, _03807_);
  nor (_03854_, _03853_, _03851_);
  and (_03855_, _03854_, \oc8051_golden_model_1.TH0 [7]);
  and (_03856_, _03809_, _03824_);
  and (_03857_, _03856_, \oc8051_golden_model_1.TCON [7]);
  nor (_03858_, _03857_, _03855_);
  and (_03859_, _03817_, _03801_);
  and (_03860_, _03859_, \oc8051_golden_model_1.P1 [7]);
  not (_03861_, _03826_);
  nand (_03862_, _02452_, _02120_);
  or (_03863_, _03862_, _03861_);
  nor (_03864_, _03863_, _03851_);
  and (_03865_, _03864_, \oc8051_golden_model_1.TL1 [7]);
  nor (_03866_, _03865_, _03860_);
  and (_03867_, _03866_, _03858_);
  and (_03868_, _03801_, _03809_);
  and (_03869_, _03868_, \oc8051_golden_model_1.SCON [7]);
  nand (_03870_, _03852_, _03802_);
  nor (_03871_, _03870_, _03851_);
  and (_03872_, _03871_, \oc8051_golden_model_1.TH1 [7]);
  nor (_03873_, _03872_, _03869_);
  nor (_03874_, _02859_, _02028_);
  nor (_03875_, _03862_, _03851_);
  and (_03876_, _03875_, _03874_);
  and (_03877_, _03876_, \oc8051_golden_model_1.TL0 [7]);
  and (_03878_, _03804_, _03824_);
  and (_03879_, _03878_, \oc8051_golden_model_1.TMOD [7]);
  nor (_03880_, _03879_, _03877_);
  and (_03881_, _03880_, _03873_);
  and (_03882_, _03881_, _03867_);
  and (_03883_, _03882_, _03850_);
  and (_03884_, _03883_, _03834_);
  and (_03885_, _03817_, _03824_);
  and (_03886_, _03885_, \oc8051_golden_model_1.P0 [7]);
  not (_03887_, _03886_);
  nand (_03888_, _03816_, _03826_);
  nor (_03889_, _03888_, _03851_);
  and (_03890_, _03889_, \oc8051_golden_model_1.DPH [7]);
  not (_03891_, _03890_);
  nand (_03892_, _03816_, _03802_);
  nor (_03893_, _03892_, _03851_);
  and (_03894_, _03893_, \oc8051_golden_model_1.SP [7]);
  nand (_03895_, _03816_, _03874_);
  nor (_03896_, _03895_, _03851_);
  and (_03897_, _03896_, \oc8051_golden_model_1.DPL [7]);
  nor (_03898_, _03897_, _03894_);
  and (_03899_, _03898_, _03891_);
  and (_03900_, _03899_, _03887_);
  and (_03901_, _03900_, _03884_);
  and (_03902_, _03901_, _03797_);
  not (_03903_, _03902_);
  not (_03904_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_03905_, _02793_, _03904_);
  not (_03906_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_03907_, _02941_, _03906_);
  and (_03908_, _03907_, _02939_);
  nand (_03909_, _03908_, _03905_);
  not (_03910_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_03911_, _02941_, _03910_);
  not (_03912_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_03913_, _02793_, _03912_);
  and (_03914_, _03913_, _02947_);
  nand (_03915_, _03914_, _03911_);
  nand (_03916_, _03915_, _03909_);
  nand (_03917_, _03916_, _02542_);
  not (_03918_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_03919_, _02941_, _03918_);
  not (_03920_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_03921_, _02793_, _03920_);
  and (_03922_, _03921_, _02947_);
  nand (_03923_, _03922_, _03919_);
  not (_03924_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_03925_, _02793_, _03924_);
  not (_03926_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_03927_, _02941_, _03926_);
  and (_03928_, _03927_, _02939_);
  nand (_03929_, _03928_, _03925_);
  nand (_03930_, _03929_, _03923_);
  nand (_03931_, _03930_, _02954_);
  nand (_03932_, _03931_, _03917_);
  nand (_03933_, _03932_, _02379_);
  not (_03934_, \oc8051_golden_model_1.IRAM[11] [6]);
  or (_03935_, _02941_, _03934_);
  not (_03936_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_03937_, _02793_, _03936_);
  and (_03938_, _03937_, _02947_);
  nand (_03939_, _03938_, _03935_);
  not (_03940_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_03941_, _02793_, _03940_);
  not (_03942_, \oc8051_golden_model_1.IRAM[9] [6]);
  or (_03943_, _02941_, _03942_);
  and (_03944_, _03943_, _02939_);
  nand (_03945_, _03944_, _03941_);
  nand (_03946_, _03945_, _03939_);
  nand (_03947_, _03946_, _02542_);
  not (_03948_, \oc8051_golden_model_1.IRAM[15] [6]);
  or (_03949_, _02941_, _03948_);
  not (_03950_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_03951_, _02793_, _03950_);
  and (_03952_, _03951_, _02947_);
  nand (_03953_, _03952_, _03949_);
  not (_03954_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_03955_, _02793_, _03954_);
  not (_03956_, \oc8051_golden_model_1.IRAM[13] [6]);
  or (_03957_, _02941_, _03956_);
  and (_03958_, _03957_, _02939_);
  nand (_03959_, _03958_, _03955_);
  nand (_03960_, _03959_, _03953_);
  nand (_03961_, _03960_, _02954_);
  nand (_03962_, _03961_, _03947_);
  nand (_03963_, _03962_, _02971_);
  nand (_03964_, _03963_, _03933_);
  or (_03965_, _03964_, _01952_);
  and (_03966_, _03805_, \oc8051_golden_model_1.SBUF [6]);
  and (_03967_, _03813_, \oc8051_golden_model_1.IE [6]);
  nor (_03968_, _03967_, _03966_);
  and (_03969_, _03820_, \oc8051_golden_model_1.P3 [6]);
  not (_03970_, _03969_);
  and (_03971_, _03828_, \oc8051_golden_model_1.PCON [6]);
  and (_03972_, _03830_, \oc8051_golden_model_1.P2 [6]);
  nor (_03973_, _03972_, _03971_);
  and (_03974_, _03973_, _03970_);
  and (_03975_, _03974_, _03968_);
  and (_03976_, _03844_, \oc8051_golden_model_1.IP [6]);
  and (_03977_, _03847_, \oc8051_golden_model_1.B [6]);
  nor (_03978_, _03977_, _03976_);
  and (_03979_, _03838_, \oc8051_golden_model_1.PSW [6]);
  and (_03980_, _03841_, \oc8051_golden_model_1.ACC [6]);
  nor (_03981_, _03980_, _03979_);
  and (_03982_, _03981_, _03978_);
  and (_03983_, _03854_, \oc8051_golden_model_1.TH0 [6]);
  and (_03984_, _03856_, \oc8051_golden_model_1.TCON [6]);
  nor (_03985_, _03984_, _03983_);
  and (_03986_, _03859_, \oc8051_golden_model_1.P1 [6]);
  and (_03987_, _03864_, \oc8051_golden_model_1.TL1 [6]);
  nor (_03988_, _03987_, _03986_);
  and (_03989_, _03988_, _03985_);
  and (_03990_, _03868_, \oc8051_golden_model_1.SCON [6]);
  and (_03991_, _03871_, \oc8051_golden_model_1.TH1 [6]);
  nor (_03992_, _03991_, _03990_);
  and (_03993_, _03876_, \oc8051_golden_model_1.TL0 [6]);
  and (_03994_, _03878_, \oc8051_golden_model_1.TMOD [6]);
  nor (_03995_, _03994_, _03993_);
  and (_03996_, _03995_, _03992_);
  and (_03997_, _03996_, _03989_);
  and (_03998_, _03997_, _03982_);
  and (_03999_, _03998_, _03975_);
  and (_04000_, _03885_, \oc8051_golden_model_1.P0 [6]);
  not (_04001_, _04000_);
  and (_04002_, _03889_, \oc8051_golden_model_1.DPH [6]);
  not (_04003_, _04002_);
  and (_04004_, _03893_, \oc8051_golden_model_1.SP [6]);
  and (_04005_, _03896_, \oc8051_golden_model_1.DPL [6]);
  nor (_04006_, _04005_, _04004_);
  and (_04007_, _04006_, _04003_);
  and (_04008_, _04007_, _04001_);
  and (_04009_, _04008_, _03999_);
  and (_04010_, _04009_, _03965_);
  not (_04011_, _04010_);
  nand (_04012_, _02941_, \oc8051_golden_model_1.IRAM[0] [5]);
  nand (_04013_, _02793_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_04014_, _04013_, _02939_);
  nand (_04015_, _04014_, _04012_);
  nand (_04016_, _02793_, \oc8051_golden_model_1.IRAM[3] [5]);
  nand (_04017_, _02941_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_04018_, _04017_, _02947_);
  nand (_04019_, _04018_, _04016_);
  nand (_04020_, _04019_, _04015_);
  nand (_04021_, _04020_, _02542_);
  nand (_04022_, _02793_, \oc8051_golden_model_1.IRAM[7] [5]);
  nand (_04023_, _02941_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_04024_, _04023_, _02947_);
  nand (_04025_, _04024_, _04022_);
  nand (_04026_, _02941_, \oc8051_golden_model_1.IRAM[4] [5]);
  nand (_04027_, _02793_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_04028_, _04027_, _02939_);
  nand (_04029_, _04028_, _04026_);
  nand (_04030_, _04029_, _04025_);
  nand (_04031_, _04030_, _02954_);
  nand (_04032_, _04031_, _04021_);
  nand (_04033_, _04032_, _02379_);
  nand (_04034_, _02793_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_04035_, _02941_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_04036_, _04035_, _02947_);
  nand (_04037_, _04036_, _04034_);
  nand (_04038_, _02941_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_04039_, _02793_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_04040_, _04039_, _02939_);
  nand (_04041_, _04040_, _04038_);
  nand (_04042_, _04041_, _04037_);
  nand (_04043_, _04042_, _02542_);
  nand (_04044_, _02793_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_04045_, _02941_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_04046_, _04045_, _02947_);
  nand (_04047_, _04046_, _04044_);
  nand (_04048_, _02941_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_04049_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_04050_, _02941_, _04049_);
  and (_04051_, _04050_, _02939_);
  nand (_04052_, _04051_, _04048_);
  nand (_04053_, _04052_, _04047_);
  nand (_04054_, _04053_, _02954_);
  nand (_04055_, _04054_, _04043_);
  nand (_04056_, _04055_, _02971_);
  nand (_04057_, _04056_, _04033_);
  or (_04058_, _04057_, _01952_);
  and (_04059_, _03828_, \oc8051_golden_model_1.PCON [5]);
  not (_04060_, _04059_);
  and (_04061_, _03805_, \oc8051_golden_model_1.SBUF [5]);
  and (_04062_, _03813_, \oc8051_golden_model_1.IE [5]);
  nor (_04063_, _04062_, _04061_);
  and (_04064_, _04063_, _04060_);
  and (_04065_, _03830_, \oc8051_golden_model_1.P2 [5]);
  and (_04066_, _03820_, \oc8051_golden_model_1.P3 [5]);
  nor (_04067_, _04066_, _04065_);
  and (_04068_, _04067_, _04064_);
  and (_04069_, _03838_, \oc8051_golden_model_1.PSW [5]);
  and (_04070_, _03847_, \oc8051_golden_model_1.B [5]);
  nor (_04071_, _04070_, _04069_);
  and (_04072_, _03844_, \oc8051_golden_model_1.IP [5]);
  and (_04073_, _03841_, \oc8051_golden_model_1.ACC [5]);
  nor (_04074_, _04073_, _04072_);
  and (_04075_, _04074_, _04071_);
  and (_04076_, _03856_, \oc8051_golden_model_1.TCON [5]);
  and (_04077_, _03854_, \oc8051_golden_model_1.TH0 [5]);
  nor (_04078_, _04077_, _04076_);
  and (_04079_, _03859_, \oc8051_golden_model_1.P1 [5]);
  and (_04080_, _03864_, \oc8051_golden_model_1.TL1 [5]);
  nor (_04081_, _04080_, _04079_);
  and (_04082_, _04081_, _04078_);
  and (_04083_, _03868_, \oc8051_golden_model_1.SCON [5]);
  and (_04084_, _03871_, \oc8051_golden_model_1.TH1 [5]);
  nor (_04085_, _04084_, _04083_);
  and (_04086_, _03878_, \oc8051_golden_model_1.TMOD [5]);
  and (_04087_, _03876_, \oc8051_golden_model_1.TL0 [5]);
  nor (_04088_, _04087_, _04086_);
  and (_04089_, _04088_, _04085_);
  and (_04090_, _04089_, _04082_);
  and (_04091_, _04090_, _04075_);
  and (_04092_, _04091_, _04068_);
  and (_04093_, _03885_, \oc8051_golden_model_1.P0 [5]);
  not (_04094_, _04093_);
  and (_04095_, _03889_, \oc8051_golden_model_1.DPH [5]);
  not (_04096_, _04095_);
  and (_04097_, _03893_, \oc8051_golden_model_1.SP [5]);
  and (_04098_, _03896_, \oc8051_golden_model_1.DPL [5]);
  nor (_04099_, _04098_, _04097_);
  and (_04100_, _04099_, _04096_);
  and (_04101_, _04100_, _04094_);
  and (_04102_, _04101_, _04092_);
  and (_04103_, _04102_, _04058_);
  not (_04104_, _04103_);
  or (_04105_, _03434_, _01952_);
  and (_04106_, _03805_, \oc8051_golden_model_1.SBUF [3]);
  and (_04107_, _03813_, \oc8051_golden_model_1.IE [3]);
  nor (_04108_, _04107_, _04106_);
  and (_04109_, _03820_, \oc8051_golden_model_1.P3 [3]);
  not (_04110_, _04109_);
  and (_04111_, _03828_, \oc8051_golden_model_1.PCON [3]);
  and (_04112_, _03830_, \oc8051_golden_model_1.P2 [3]);
  nor (_04113_, _04112_, _04111_);
  and (_04114_, _04113_, _04110_);
  and (_04115_, _04114_, _04108_);
  and (_04116_, _03838_, \oc8051_golden_model_1.PSW [3]);
  not (_04117_, _04116_);
  and (_04118_, _03844_, \oc8051_golden_model_1.IP [3]);
  not (_04119_, _04118_);
  and (_04120_, _03841_, \oc8051_golden_model_1.ACC [3]);
  and (_04121_, _03847_, \oc8051_golden_model_1.B [3]);
  nor (_04122_, _04121_, _04120_);
  and (_04123_, _04122_, _04119_);
  and (_04124_, _04123_, _04117_);
  and (_04125_, _03854_, \oc8051_golden_model_1.TH0 [3]);
  and (_04126_, _03856_, \oc8051_golden_model_1.TCON [3]);
  nor (_04127_, _04126_, _04125_);
  and (_04128_, _03859_, \oc8051_golden_model_1.P1 [3]);
  and (_04129_, _03864_, \oc8051_golden_model_1.TL1 [3]);
  nor (_04130_, _04129_, _04128_);
  and (_04131_, _04130_, _04127_);
  and (_04132_, _03868_, \oc8051_golden_model_1.SCON [3]);
  and (_04133_, _03871_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04134_, _04133_, _04132_);
  and (_04135_, _03876_, \oc8051_golden_model_1.TL0 [3]);
  and (_04136_, _03878_, \oc8051_golden_model_1.TMOD [3]);
  nor (_04137_, _04136_, _04135_);
  and (_04138_, _04137_, _04134_);
  and (_04139_, _04138_, _04131_);
  and (_04140_, _04139_, _04124_);
  and (_04141_, _04140_, _04115_);
  and (_04142_, _03885_, \oc8051_golden_model_1.P0 [3]);
  not (_04143_, _04142_);
  and (_04144_, _03889_, \oc8051_golden_model_1.DPH [3]);
  not (_04145_, _04144_);
  and (_04146_, _03893_, \oc8051_golden_model_1.SP [3]);
  and (_04147_, _03896_, \oc8051_golden_model_1.DPL [3]);
  nor (_04148_, _04147_, _04146_);
  and (_04149_, _04148_, _04145_);
  and (_04150_, _04149_, _04143_);
  and (_04151_, _04150_, _04141_);
  and (_04152_, _04151_, _04105_);
  not (_04153_, _04152_);
  or (_04154_, _03161_, _01952_);
  and (_04155_, _03838_, \oc8051_golden_model_1.PSW [1]);
  and (_04156_, _03841_, \oc8051_golden_model_1.ACC [1]);
  nor (_04157_, _04156_, _04155_);
  and (_04158_, _03844_, \oc8051_golden_model_1.IP [1]);
  and (_04159_, _03847_, \oc8051_golden_model_1.B [1]);
  nor (_04160_, _04159_, _04158_);
  and (_04161_, _04160_, _04157_);
  and (_04162_, _03808_, _03825_);
  and (_04163_, _04162_, \oc8051_golden_model_1.P0 [1]);
  not (_04164_, _04163_);
  and (_04165_, _03859_, \oc8051_golden_model_1.P1 [1]);
  not (_04166_, _04165_);
  and (_04167_, _03830_, \oc8051_golden_model_1.P2 [1]);
  and (_04168_, _03820_, \oc8051_golden_model_1.P3 [1]);
  nor (_04169_, _04168_, _04167_);
  and (_04170_, _04169_, _04166_);
  and (_04171_, _04170_, _04164_);
  and (_04172_, _04171_, _04161_);
  and (_04173_, _03828_, \oc8051_golden_model_1.PCON [1]);
  not (_04174_, _04173_);
  and (_04175_, _03805_, \oc8051_golden_model_1.SBUF [1]);
  and (_04176_, _03813_, \oc8051_golden_model_1.IE [1]);
  nor (_04177_, _04176_, _04175_);
  and (_04178_, _04177_, _04174_);
  and (_04179_, _03874_, _02452_);
  and (_04180_, _04179_, _03825_);
  and (_04181_, _04180_, \oc8051_golden_model_1.DPL [1]);
  and (_04182_, _03803_, _03825_);
  and (_04183_, _04182_, \oc8051_golden_model_1.SP [1]);
  nor (_04184_, _04183_, _04181_);
  and (_04185_, _04184_, _04178_);
  and (_04186_, _04185_, _04172_);
  and (_04187_, _03876_, \oc8051_golden_model_1.TL0 [1]);
  not (_04188_, _04187_);
  and (_04189_, _03878_, \oc8051_golden_model_1.TMOD [1]);
  and (_04190_, _03868_, \oc8051_golden_model_1.SCON [1]);
  nor (_04191_, _04190_, _04189_);
  and (_04192_, _03856_, \oc8051_golden_model_1.TCON [1]);
  and (_04193_, _03871_, \oc8051_golden_model_1.TH1 [1]);
  nor (_04194_, _04193_, _04192_);
  and (_04195_, _04194_, _04191_);
  and (_04196_, _04195_, _04188_);
  and (_04197_, _03875_, _03826_);
  and (_04198_, _04197_, \oc8051_golden_model_1.TL1 [1]);
  not (_04199_, _04198_);
  and (_04200_, _03854_, \oc8051_golden_model_1.TH0 [1]);
  and (_04201_, _03826_, _02452_);
  and (_04202_, _04201_, _03825_);
  and (_04203_, _04202_, \oc8051_golden_model_1.DPH [1]);
  nor (_04204_, _04203_, _04200_);
  and (_04205_, _04204_, _04199_);
  and (_04206_, _04205_, _04196_);
  and (_04207_, _04206_, _04186_);
  and (_04208_, _04207_, _04154_);
  not (_04209_, _04208_);
  or (_04210_, _03020_, _01952_);
  and (_04211_, _03871_, \oc8051_golden_model_1.TH1 [0]);
  and (_04212_, _03805_, \oc8051_golden_model_1.SBUF [0]);
  nor (_04213_, _04212_, _04211_);
  and (_04214_, _03854_, \oc8051_golden_model_1.TH0 [0]);
  and (_04215_, _03868_, \oc8051_golden_model_1.SCON [0]);
  nor (_04216_, _04215_, _04214_);
  and (_04217_, _04216_, _04213_);
  and (_04218_, _04202_, \oc8051_golden_model_1.DPH [0]);
  not (_04219_, _04218_);
  and (_04220_, _03878_, \oc8051_golden_model_1.TMOD [0]);
  and (_04221_, _03813_, \oc8051_golden_model_1.IE [0]);
  nor (_04222_, _04221_, _04220_);
  and (_04223_, _04222_, _04219_);
  and (_04224_, _03876_, \oc8051_golden_model_1.TL0 [0]);
  and (_04225_, _04197_, \oc8051_golden_model_1.TL1 [0]);
  nor (_04226_, _04225_, _04224_);
  and (_04227_, _04226_, _04223_);
  and (_04228_, _04227_, _04217_);
  and (_04229_, _03828_, \oc8051_golden_model_1.PCON [0]);
  not (_04230_, _04229_);
  and (_04231_, _03856_, \oc8051_golden_model_1.TCON [0]);
  not (_04232_, _04231_);
  and (_04233_, _03844_, \oc8051_golden_model_1.IP [0]);
  and (_04234_, _03847_, \oc8051_golden_model_1.B [0]);
  nor (_04235_, _04234_, _04233_);
  and (_04236_, _03838_, \oc8051_golden_model_1.PSW [0]);
  and (_04237_, _03841_, \oc8051_golden_model_1.ACC [0]);
  nor (_04238_, _04237_, _04236_);
  and (_04239_, _04238_, _04235_);
  and (_04240_, _04239_, _04232_);
  and (_04241_, _04240_, _04230_);
  and (_04242_, _04180_, \oc8051_golden_model_1.DPL [0]);
  and (_04243_, _04182_, \oc8051_golden_model_1.SP [0]);
  nor (_04244_, _04243_, _04242_);
  and (_04245_, _04162_, \oc8051_golden_model_1.P0 [0]);
  not (_04246_, _04245_);
  and (_04247_, _03859_, \oc8051_golden_model_1.P1 [0]);
  not (_04248_, _04247_);
  and (_04249_, _03830_, \oc8051_golden_model_1.P2 [0]);
  and (_04250_, _03820_, \oc8051_golden_model_1.P3 [0]);
  nor (_04251_, _04250_, _04249_);
  and (_04252_, _04251_, _04248_);
  and (_04253_, _04252_, _04246_);
  and (_04254_, _04253_, _04244_);
  and (_04255_, _04254_, _04241_);
  and (_04256_, _04255_, _04228_);
  nand (_04257_, _04256_, _04210_);
  and (_04258_, _04257_, _04209_);
  or (_04259_, _03624_, _01952_);
  and (_04260_, _03854_, \oc8051_golden_model_1.TH0 [2]);
  and (_04261_, _03871_, \oc8051_golden_model_1.TH1 [2]);
  nor (_04262_, _04261_, _04260_);
  and (_04263_, _03878_, \oc8051_golden_model_1.TMOD [2]);
  and (_04264_, _03868_, \oc8051_golden_model_1.SCON [2]);
  nor (_04265_, _04264_, _04263_);
  and (_04266_, _04265_, _04262_);
  and (_04267_, _04197_, \oc8051_golden_model_1.TL1 [2]);
  not (_04268_, _04267_);
  and (_04269_, _03876_, \oc8051_golden_model_1.TL0 [2]);
  and (_04270_, _04202_, \oc8051_golden_model_1.DPH [2]);
  nor (_04271_, _04270_, _04269_);
  and (_04272_, _04271_, _04268_);
  and (_04273_, _04272_, _04266_);
  and (_04274_, _03828_, \oc8051_golden_model_1.PCON [2]);
  not (_04275_, _04274_);
  and (_04276_, _03844_, \oc8051_golden_model_1.IP [2]);
  not (_04277_, _04276_);
  and (_04278_, _03838_, \oc8051_golden_model_1.PSW [2]);
  and (_04279_, _03847_, \oc8051_golden_model_1.B [2]);
  nor (_04280_, _04279_, _04278_);
  and (_04281_, _04280_, _04277_);
  and (_04282_, _03805_, \oc8051_golden_model_1.SBUF [2]);
  not (_04283_, _04282_);
  and (_04284_, _03813_, \oc8051_golden_model_1.IE [2]);
  and (_04285_, _03841_, \oc8051_golden_model_1.ACC [2]);
  nor (_04286_, _04285_, _04284_);
  and (_04287_, _04286_, _04283_);
  and (_04288_, _04287_, _04281_);
  and (_04289_, _04288_, _04275_);
  and (_04290_, _04180_, \oc8051_golden_model_1.DPL [2]);
  not (_04291_, _04290_);
  and (_04292_, _03856_, \oc8051_golden_model_1.TCON [2]);
  and (_04293_, _04182_, \oc8051_golden_model_1.SP [2]);
  nor (_04294_, _04293_, _04292_);
  and (_04295_, _04294_, _04291_);
  and (_04296_, _04162_, \oc8051_golden_model_1.P0 [2]);
  not (_04297_, _04296_);
  and (_04298_, _03859_, \oc8051_golden_model_1.P1 [2]);
  not (_04299_, _04298_);
  and (_04300_, _03830_, \oc8051_golden_model_1.P2 [2]);
  and (_04301_, _03820_, \oc8051_golden_model_1.P3 [2]);
  nor (_04302_, _04301_, _04300_);
  and (_04303_, _04302_, _04299_);
  and (_04304_, _04303_, _04297_);
  and (_04305_, _04304_, _04295_);
  and (_04306_, _04305_, _04289_);
  and (_04307_, _04306_, _04273_);
  and (_04308_, _04307_, _04259_);
  not (_04309_, _04308_);
  and (_04310_, _04309_, _04258_);
  and (_04311_, _04310_, _04153_);
  not (_04312_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_04313_, _02793_, _04312_);
  not (_04314_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_04315_, _02941_, _04314_);
  and (_04316_, _04315_, _02939_);
  nand (_04317_, _04316_, _04313_);
  not (_04318_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_04319_, _02941_, _04318_);
  not (_04320_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_04321_, _02793_, _04320_);
  and (_04322_, _04321_, _02947_);
  nand (_04323_, _04322_, _04319_);
  nand (_04324_, _04323_, _04317_);
  nand (_04325_, _04324_, _02542_);
  not (_04326_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_04327_, _02941_, _04326_);
  not (_04328_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_04329_, _02793_, _04328_);
  and (_04330_, _04329_, _02947_);
  nand (_04331_, _04330_, _04327_);
  not (_04332_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_04333_, _02793_, _04332_);
  not (_04334_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_04335_, _02941_, _04334_);
  and (_04336_, _04335_, _02939_);
  nand (_04337_, _04336_, _04333_);
  nand (_04338_, _04337_, _04331_);
  nand (_04339_, _04338_, _02954_);
  nand (_04340_, _04339_, _04325_);
  nand (_04341_, _04340_, _02379_);
  not (_04342_, \oc8051_golden_model_1.IRAM[11] [4]);
  or (_04343_, _02941_, _04342_);
  not (_04344_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_04345_, _02793_, _04344_);
  and (_04346_, _04345_, _02947_);
  nand (_04347_, _04346_, _04343_);
  not (_04348_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_04349_, _02793_, _04348_);
  not (_04350_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_04351_, _02941_, _04350_);
  and (_04352_, _04351_, _02939_);
  nand (_04353_, _04352_, _04349_);
  nand (_04354_, _04353_, _04347_);
  nand (_04355_, _04354_, _02542_);
  not (_04356_, \oc8051_golden_model_1.IRAM[15] [4]);
  or (_04357_, _02941_, _04356_);
  not (_04358_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_04359_, _02793_, _04358_);
  and (_04360_, _04359_, _02947_);
  nand (_04361_, _04360_, _04357_);
  not (_04362_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_04363_, _02793_, _04362_);
  not (_04364_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_04365_, _02941_, _04364_);
  and (_04366_, _04365_, _02939_);
  nand (_04367_, _04366_, _04363_);
  nand (_04368_, _04367_, _04361_);
  nand (_04369_, _04368_, _02954_);
  nand (_04370_, _04369_, _04355_);
  nand (_04371_, _04370_, _02971_);
  nand (_04372_, _04371_, _04341_);
  or (_04373_, _04372_, _01952_);
  and (_04374_, _03838_, \oc8051_golden_model_1.PSW [4]);
  and (_04375_, _03847_, \oc8051_golden_model_1.B [4]);
  nor (_04376_, _04375_, _04374_);
  and (_04377_, _03844_, \oc8051_golden_model_1.IP [4]);
  and (_04378_, _03841_, \oc8051_golden_model_1.ACC [4]);
  nor (_04379_, _04378_, _04377_);
  and (_04380_, _04379_, _04376_);
  nand (_04381_, _04162_, \oc8051_golden_model_1.P0 [4]);
  and (_04382_, _03859_, \oc8051_golden_model_1.P1 [4]);
  not (_04383_, _04382_);
  and (_04384_, _03830_, \oc8051_golden_model_1.P2 [4]);
  and (_04385_, _03820_, \oc8051_golden_model_1.P3 [4]);
  nor (_04386_, _04385_, _04384_);
  and (_04387_, _04386_, _04383_);
  and (_04388_, _04387_, _04381_);
  and (_04389_, _04388_, _04380_);
  and (_04390_, _03828_, \oc8051_golden_model_1.PCON [4]);
  not (_04391_, _04390_);
  and (_04392_, _03805_, \oc8051_golden_model_1.SBUF [4]);
  and (_04393_, _03813_, \oc8051_golden_model_1.IE [4]);
  nor (_04394_, _04393_, _04392_);
  and (_04395_, _04394_, _04391_);
  and (_04396_, _04180_, \oc8051_golden_model_1.DPL [4]);
  and (_04397_, _04182_, \oc8051_golden_model_1.SP [4]);
  nor (_04398_, _04397_, _04396_);
  and (_04399_, _04398_, _04395_);
  and (_04400_, _04399_, _04389_);
  and (_04401_, _03876_, \oc8051_golden_model_1.TL0 [4]);
  not (_04402_, _04401_);
  and (_04403_, _03878_, \oc8051_golden_model_1.TMOD [4]);
  and (_04404_, _03868_, \oc8051_golden_model_1.SCON [4]);
  nor (_04405_, _04404_, _04403_);
  and (_04406_, _03856_, \oc8051_golden_model_1.TCON [4]);
  and (_04407_, _03871_, \oc8051_golden_model_1.TH1 [4]);
  nor (_04408_, _04407_, _04406_);
  and (_04409_, _04408_, _04405_);
  and (_04410_, _04409_, _04402_);
  and (_04411_, _04197_, \oc8051_golden_model_1.TL1 [4]);
  not (_04412_, _04411_);
  and (_04413_, _03854_, \oc8051_golden_model_1.TH0 [4]);
  and (_04414_, _04202_, \oc8051_golden_model_1.DPH [4]);
  nor (_04415_, _04414_, _04413_);
  and (_04416_, _04415_, _04412_);
  and (_04417_, _04416_, _04410_);
  and (_04418_, _04417_, _04400_);
  and (_04419_, _04418_, _04373_);
  not (_04420_, _04419_);
  and (_04421_, _04420_, _04311_);
  and (_04422_, _04421_, _04104_);
  and (_04423_, _04422_, _04011_);
  nor (_04424_, _04423_, _03903_);
  and (_04425_, _04423_, _03903_);
  nor (_04426_, _04425_, _04424_);
  and (_04427_, _04426_, _03098_);
  and (_04428_, _02319_, _00182_);
  and (_04429_, _02286_, _00195_);
  nor (_04430_, _04429_, _04428_);
  and (_04431_, _02308_, _00134_);
  and (_04432_, _02281_, _00155_);
  nor (_04433_, _04432_, _04431_);
  and (_04434_, _04433_, _04430_);
  and (_04435_, _02301_, _00188_);
  and (_04436_, _02303_, _00191_);
  nor (_04437_, _04436_, _04435_);
  and (_04438_, _02273_, _00217_);
  and (_04439_, _02270_, _00212_);
  nor (_04440_, _04439_, _04438_);
  and (_04441_, _04440_, _04437_);
  and (_04442_, _04441_, _04434_);
  and (_04443_, _02312_, _00165_);
  and (_04444_, _02296_, _00179_);
  nor (_04445_, _04444_, _04443_);
  and (_04446_, _02306_, _00115_);
  and (_04447_, _02277_, _00143_);
  nor (_04448_, _04447_, _04446_);
  and (_04449_, _04448_, _04445_);
  and (_04450_, _02290_, _00199_);
  and (_04451_, _02314_, _00206_);
  nor (_04452_, _04451_, _04450_);
  and (_04453_, _02294_, _00149_);
  and (_04454_, _02317_, _00175_);
  nor (_04455_, _04454_, _04453_);
  and (_04456_, _04455_, _04452_);
  and (_04457_, _04456_, _04449_);
  and (_04458_, _04457_, _04442_);
  nand (_04459_, _04458_, _01996_);
  not (_04460_, _01767_);
  not (_04461_, _03040_);
  not (_04462_, _01984_);
  nor (_04463_, _02826_, _04462_);
  not (_04464_, _02411_);
  and (_04465_, _04464_, _02122_);
  and (_04466_, _04465_, _04463_);
  and (_04467_, _03819_, _04466_);
  and (_04468_, _04467_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_04469_, _02411_, _02122_);
  and (_04470_, _04469_, _04463_);
  and (_04471_, _04470_, _03801_);
  and (_04472_, _04471_, \oc8051_golden_model_1.SCON [7]);
  and (_04473_, _04470_, _03812_);
  and (_04474_, _04473_, \oc8051_golden_model_1.IE [7]);
  nor (_04475_, _04474_, _04472_);
  and (_04476_, _03837_, _04466_);
  and (_04477_, _04476_, \oc8051_golden_model_1.PSW [7]);
  and (_04478_, _03846_, _04466_);
  and (_04479_, _04478_, \oc8051_golden_model_1.B [7]);
  nor (_04480_, _04479_, _04477_);
  and (_04481_, _04470_, _03819_);
  and (_04482_, _04481_, \oc8051_golden_model_1.IP [7]);
  and (_04483_, _03840_, _04466_);
  and (_04484_, _04483_, \oc8051_golden_model_1.ACC [7]);
  nor (_04485_, _04484_, _04482_);
  and (_04486_, _04485_, _04480_);
  and (_04487_, _04470_, _03824_);
  and (_04488_, _04487_, \oc8051_golden_model_1.TCON [7]);
  and (_04489_, _03801_, _04466_);
  and (_04490_, _04489_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_04491_, _04490_, _04488_);
  and (_04492_, _03812_, _04466_);
  and (_04493_, _04492_, \oc8051_golden_model_1.P2INREG [7]);
  and (_04494_, _03825_, \oc8051_golden_model_1.P0INREG [7]);
  nor (_04495_, _04494_, _04493_);
  and (_04496_, _04495_, _04491_);
  and (_04497_, _04496_, _04486_);
  nand (_04498_, _04497_, _04475_);
  nor (_04499_, _04498_, _04468_);
  and (_04500_, _04499_, _03797_);
  nor (_04501_, _04500_, _03827_);
  and (_04502_, _03827_, \oc8051_golden_model_1.PSW [7]);
  nor (_04503_, _04502_, _04501_);
  nor (_04504_, _04503_, _04461_);
  not (_04505_, _03024_);
  and (_04506_, _04467_, \oc8051_golden_model_1.P3 [7]);
  and (_04507_, _04492_, \oc8051_golden_model_1.P2 [7]);
  or (_04508_, _04507_, _04506_);
  nor (_04509_, _04508_, _04488_);
  and (_04510_, _03825_, \oc8051_golden_model_1.P0 [7]);
  and (_04511_, _04489_, \oc8051_golden_model_1.P1 [7]);
  nor (_04512_, _04511_, _04510_);
  and (_04513_, _04512_, _04475_);
  and (_04514_, _04513_, _04486_);
  and (_04515_, _04514_, _04509_);
  and (_04516_, _04515_, _03797_);
  nor (_04517_, _04516_, _03827_);
  or (_04518_, _04517_, _04505_);
  not (_04519_, _03005_);
  not (_04520_, _03827_);
  nand (_04521_, _04516_, _04520_);
  or (_04522_, _04521_, _04519_);
  not (_04523_, _03796_);
  and (_04524_, _04372_, _04057_);
  and (_04525_, _03161_, _03020_);
  and (_04526_, _03624_, _03434_);
  and (_04527_, _04526_, _04525_);
  and (_04528_, _04527_, _04524_);
  and (_04529_, _04528_, _03964_);
  or (_04530_, _04529_, _04523_);
  nand (_04531_, _04529_, _04523_);
  and (_04532_, _04531_, _04530_);
  nor (_04533_, _02926_, _02511_);
  and (_04534_, _04533_, _03177_);
  not (_04535_, _04534_);
  and (_04536_, _04535_, _04532_);
  and (_04537_, _01747_, \oc8051_golden_model_1.ACC [7]);
  and (_04538_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_04539_, _04538_, \oc8051_golden_model_1.PC [6]);
  and (_04540_, _04539_, _01824_);
  nor (_04541_, _04540_, \oc8051_golden_model_1.PC [7]);
  and (_04542_, _04540_, \oc8051_golden_model_1.PC [7]);
  nor (_04543_, _04542_, _04541_);
  not (_04544_, _04543_);
  nor (_04545_, _04544_, _01747_);
  or (_04546_, _04545_, _04537_);
  and (_04547_, _04546_, _04534_);
  or (_04548_, _04547_, _02079_);
  or (_04549_, _04548_, _04536_);
  not (_04550_, _02079_);
  nor (_04551_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04552_, _04551_, _02518_);
  nor (_04553_, _04552_, _02362_);
  nor (_04554_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04555_, _04554_, _02362_);
  and (_04556_, _04555_, _01986_);
  nor (_04557_, _04556_, _04553_);
  nor (_04558_, _04557_, _02520_);
  not (_04559_, _03041_);
  and (_04560_, _03434_, _04559_);
  not (_04561_, _02520_);
  and (_04562_, _03041_, _01983_);
  or (_04563_, _04562_, _04561_);
  nor (_04564_, _04563_, _04560_);
  nor (_04565_, _04564_, _04558_);
  nor (_04566_, _04551_, _02518_);
  nor (_04567_, _04566_, _04552_);
  nor (_04568_, _04567_, _02520_);
  not (_04569_, _04568_);
  nand (_04570_, _03624_, _04559_);
  and (_04571_, _03041_, _02452_);
  nor (_04572_, _04571_, _04561_);
  nand (_04573_, _04572_, _04570_);
  and (_04574_, _04573_, _04569_);
  nor (_04575_, _03161_, _03041_);
  nor (_04576_, _02859_, _04559_);
  or (_04577_, _04576_, _04575_);
  nand (_04578_, _04577_, _02520_);
  nor (_04579_, _03108_, _02520_);
  not (_04580_, _04579_);
  and (_04581_, _04580_, _04578_);
  or (_04582_, _03002_, _03041_);
  and (_04583_, _03041_, _02027_);
  nor (_04584_, _04583_, _04561_);
  nand (_04585_, _04584_, _04582_);
  nor (_04586_, _02520_, \oc8051_golden_model_1.SP [0]);
  not (_04587_, _04586_);
  and (_04588_, _04587_, _04585_);
  or (_04589_, _04588_, _03750_);
  nand (_04590_, _04587_, _04585_);
  or (_04591_, _04590_, _03748_);
  nand (_04592_, _04591_, _04589_);
  and (_04593_, _04592_, _04581_);
  or (_04594_, _04590_, \oc8051_golden_model_1.IRAM[2] [7]);
  nand (_04595_, _04580_, _04578_);
  or (_04596_, _04588_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_04597_, _04596_, _04595_);
  and (_04598_, _04597_, _04594_);
  nor (_04599_, _04598_, _04593_);
  nand (_04600_, _04599_, _04574_);
  not (_04601_, _04574_);
  or (_04602_, _04588_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_04603_, _04590_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_04604_, _04603_, _04581_);
  and (_04605_, _04604_, _04602_);
  or (_04606_, _04590_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_04607_, _04588_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_04608_, _04607_, _04595_);
  and (_04609_, _04608_, _04606_);
  nor (_04610_, _04609_, _04605_);
  nand (_04611_, _04610_, _04601_);
  nand (_04612_, _04611_, _04600_);
  nand (_04613_, _04612_, _04565_);
  not (_04614_, _04565_);
  or (_04615_, _04590_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_04616_, _04588_, \oc8051_golden_model_1.IRAM[9] [7]);
  nand (_04617_, _04616_, _04615_);
  nand (_04618_, _04617_, _04581_);
  or (_04619_, _04590_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_04620_, _04588_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_04621_, _04620_, _04619_);
  nand (_04622_, _04621_, _04595_);
  nand (_04623_, _04622_, _04618_);
  nand (_04624_, _04623_, _04574_);
  or (_04625_, _04590_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_04626_, _04588_, \oc8051_golden_model_1.IRAM[13] [7]);
  nand (_04627_, _04626_, _04625_);
  nand (_04628_, _04627_, _04581_);
  or (_04629_, _04590_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_04630_, _04588_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_04631_, _04630_, _04629_);
  nand (_04632_, _04631_, _04595_);
  nand (_04633_, _04632_, _04628_);
  nand (_04634_, _04633_, _04601_);
  nand (_04635_, _04634_, _04624_);
  nand (_04636_, _04635_, _04614_);
  and (_04637_, _04636_, _04613_);
  or (_04638_, _04637_, _04550_);
  and (_04639_, _04638_, _04549_);
  or (_04640_, _04639_, _03007_);
  and (_04641_, _04419_, _04103_);
  not (_04642_, _04257_);
  and (_04643_, _04642_, _04208_);
  and (_04644_, _04308_, _04152_);
  and (_04645_, _04644_, _04643_);
  and (_04646_, _04645_, _04641_);
  and (_04647_, _04646_, _04010_);
  nor (_04648_, _04647_, _03903_);
  and (_04649_, _04647_, _03903_);
  nor (_04650_, _04649_, _04648_);
  or (_04651_, _04650_, _03165_);
  and (_04652_, _04651_, _04640_);
  or (_04653_, _04652_, _03005_);
  and (_04654_, _04653_, _04522_);
  or (_04655_, _04654_, _03446_);
  nor (_04656_, _04543_, _01745_);
  nor (_04657_, _04656_, _03015_);
  and (_04658_, _04657_, _04655_);
  and (_04659_, _04523_, _03015_);
  or (_04660_, _04659_, _03024_);
  or (_04661_, _04660_, _04658_);
  and (_04662_, _04661_, _04518_);
  or (_04663_, _04662_, _02052_);
  not (_04664_, _03855_);
  and (_04665_, _03880_, _04664_);
  nor (_04666_, _03865_, _03857_);
  and (_04667_, _04666_, _04665_);
  and (_04668_, _03830_, \oc8051_golden_model_1.P2INREG [7]);
  and (_04669_, _03820_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_04670_, _04669_, _04668_);
  and (_04671_, _03859_, \oc8051_golden_model_1.P1INREG [7]);
  and (_04672_, _03885_, \oc8051_golden_model_1.P0INREG [7]);
  nor (_04673_, _04672_, _04671_);
  and (_04674_, _04673_, _04670_);
  and (_04675_, _04674_, _04667_);
  not (_04676_, _03829_);
  and (_04677_, _03873_, _04676_);
  and (_04678_, _04677_, _03815_);
  and (_04679_, _03899_, _03850_);
  and (_04680_, _04679_, _04678_);
  and (_04681_, _04680_, _04675_);
  and (_04682_, _04681_, _03797_);
  nand (_04683_, _04682_, _02052_);
  and (_04684_, _04683_, _02050_);
  and (_04685_, _04684_, _04663_);
  nor (_04686_, _04516_, _04520_);
  not (_04687_, _04686_);
  and (_04688_, _04687_, _04521_);
  and (_04689_, _04688_, _02049_);
  or (_04690_, _04689_, _04685_);
  and (_04691_, _04690_, _01750_);
  or (_04692_, _04544_, _01750_);
  nand (_04693_, _04692_, _02144_);
  or (_04694_, _04693_, _04691_);
  nand (_04695_, _04682_, _02145_);
  and (_04696_, _04695_, _04694_);
  or (_04697_, _04696_, _03041_);
  nand (_04698_, _04636_, _04613_);
  or (_04699_, _04698_, _01952_);
  and (_04700_, _04681_, _03041_);
  nand (_04701_, _04700_, _04699_);
  and (_04702_, _04701_, _04461_);
  and (_04703_, _04702_, _04697_);
  or (_04704_, _04703_, _04504_);
  and (_04705_, _04704_, _04460_);
  and (_04706_, _04543_, _01767_);
  or (_04707_, _04706_, _02035_);
  or (_04708_, _04707_, _04705_);
  nand (_04709_, _03796_, _02035_);
  and (_04710_, _04709_, _04708_);
  or (_04711_, _04710_, _02033_);
  not (_04712_, _02033_);
  or (_04713_, _04637_, _04712_);
  and (_04714_, _04713_, _02039_);
  and (_04715_, _04714_, _04711_);
  not (_04716_, _04458_);
  nor (_04717_, _04716_, _03796_);
  and (_04718_, _02893_, _02679_);
  not (_04719_, _02324_);
  and (_04720_, _02494_, _04719_);
  and (_04721_, _04720_, _04718_);
  and (_04722_, _02319_, _00702_);
  and (_04723_, _02286_, _00671_);
  nor (_04724_, _04723_, _04722_);
  and (_04725_, _02306_, _00664_);
  and (_04726_, _02296_, _00695_);
  nor (_04727_, _04726_, _04725_);
  and (_04728_, _04727_, _04724_);
  and (_04729_, _02273_, _00685_);
  and (_04730_, _02270_, _00687_);
  nor (_04731_, _04730_, _04729_);
  and (_04732_, _02303_, _00666_);
  and (_04733_, _02290_, _00668_);
  nor (_04734_, _04733_, _04732_);
  and (_04735_, _04734_, _04731_);
  and (_04736_, _04735_, _04728_);
  and (_04737_, _02277_, _00706_);
  and (_04738_, _02294_, _00711_);
  nor (_04739_, _04738_, _04737_);
  and (_04740_, _02308_, _00708_);
  and (_04741_, _02281_, _00713_);
  nor (_04742_, _04741_, _04740_);
  and (_04743_, _04742_, _04739_);
  and (_04744_, _02312_, _00697_);
  and (_04745_, _02317_, _00699_);
  nor (_04746_, _04745_, _04744_);
  and (_04747_, _02301_, _00679_);
  and (_04748_, _02314_, _00683_);
  nor (_04749_, _04748_, _04747_);
  and (_04750_, _04749_, _04746_);
  and (_04751_, _04750_, _04743_);
  and (_04752_, _04751_, _04736_);
  and (_04753_, _04752_, _04716_);
  and (_04754_, _02306_, _00567_);
  and (_04755_, _02294_, _00590_);
  nor (_04756_, _04755_, _04754_);
  and (_04757_, _02303_, _00554_);
  and (_04758_, _02290_, _00558_);
  nor (_04759_, _04758_, _04757_);
  and (_04760_, _04759_, _04756_);
  and (_04761_, _02308_, _00564_);
  and (_04762_, _02277_, _00562_);
  nor (_04763_, _04762_, _04761_);
  and (_04764_, _02281_, _00577_);
  and (_04765_, _02296_, _00592_);
  nor (_04766_, _04765_, _04764_);
  and (_04767_, _04766_, _04763_);
  and (_04768_, _04767_, _04760_);
  and (_04769_, _02319_, _00580_);
  and (_04770_, _02301_, _00596_);
  nor (_04771_, _04770_, _04769_);
  and (_04772_, _02314_, _00598_);
  and (_04773_, _02273_, _00600_);
  nor (_04774_, _04773_, _04772_);
  and (_04775_, _04774_, _04771_);
  and (_04776_, _02312_, _00582_);
  and (_04777_, _02317_, _00584_);
  nor (_04778_, _04777_, _04776_);
  and (_04779_, _02286_, _00556_);
  and (_04780_, _02270_, _00602_);
  nor (_04781_, _04780_, _04779_);
  and (_04782_, _04781_, _04778_);
  and (_04783_, _04782_, _04775_);
  and (_04784_, _04783_, _04768_);
  and (_04785_, _02319_, _00635_);
  and (_04786_, _02270_, _00657_);
  nor (_04787_, _04786_, _04785_);
  and (_04788_, _02296_, _00645_);
  and (_04789_, _02286_, _00613_);
  nor (_04790_, _04789_, _04788_);
  and (_04791_, _04790_, _04787_);
  and (_04792_, _02294_, _00617_);
  and (_04793_, _02314_, _00653_);
  nor (_04794_, _04793_, _04792_);
  and (_04795_, _02277_, _00647_);
  and (_04796_, _02281_, _00633_);
  nor (_04797_, _04796_, _04795_);
  and (_04798_, _04797_, _04794_);
  and (_04799_, _04798_, _04791_);
  and (_04800_, _02308_, _00625_);
  and (_04801_, _02273_, _00655_);
  nor (_04802_, _04801_, _04800_);
  and (_04803_, _02317_, _00640_);
  and (_04804_, _02303_, _00609_);
  nor (_04805_, _04804_, _04803_);
  and (_04806_, _04805_, _04802_);
  and (_04807_, _02312_, _00637_);
  and (_04808_, _02301_, _00651_);
  nor (_04809_, _04808_, _04807_);
  and (_04810_, _02306_, _00621_);
  and (_04811_, _02290_, _00611_);
  nor (_04812_, _04811_, _04810_);
  and (_04813_, _04812_, _04809_);
  and (_04814_, _04813_, _04806_);
  and (_04815_, _04814_, _04799_);
  nor (_04816_, _04815_, _04784_);
  and (_04817_, _04816_, _04753_);
  and (_04818_, _04817_, _04721_);
  and (_04819_, _04818_, \oc8051_golden_model_1.IP [7]);
  and (_04820_, _02494_, _02324_);
  and (_04821_, _04820_, _04718_);
  nor (_04822_, _04752_, _04458_);
  and (_04823_, _04822_, _04821_);
  and (_04824_, _04823_, _04816_);
  and (_04825_, _04824_, \oc8051_golden_model_1.B [7]);
  nor (_04826_, _04825_, _04819_);
  not (_04827_, _04815_);
  and (_04828_, _04827_, _04784_);
  and (_04829_, _04828_, _04823_);
  and (_04830_, _04829_, \oc8051_golden_model_1.ACC [7]);
  not (_04831_, _04784_);
  and (_04832_, _04815_, _04831_);
  and (_04833_, _04832_, _04823_);
  and (_04834_, _04833_, \oc8051_golden_model_1.PSW [7]);
  nor (_04835_, _04834_, _04830_);
  and (_04836_, _04835_, _04826_);
  not (_04837_, _02679_);
  and (_04838_, _02893_, _04837_);
  and (_04839_, _04815_, _04784_);
  and (_04840_, _04839_, _04753_);
  nor (_04841_, _02494_, _02324_);
  and (_04842_, _04841_, _04840_);
  and (_04843_, _04842_, _04838_);
  and (_04844_, _04843_, \oc8051_golden_model_1.TH1 [7]);
  not (_04845_, _04844_);
  not (_04846_, _02893_);
  and (_04847_, _04846_, _02679_);
  and (_04848_, _04840_, _04720_);
  and (_04849_, _04848_, _04847_);
  and (_04850_, _04849_, \oc8051_golden_model_1.TL0 [7]);
  and (_04851_, _04840_, _04820_);
  and (_04852_, _04851_, _04838_);
  and (_04853_, _04852_, \oc8051_golden_model_1.SP [7]);
  nor (_04854_, _04853_, _04850_);
  and (_04855_, _04854_, _04845_);
  and (_04856_, _04855_, _04836_);
  and (_04857_, _04842_, _04718_);
  and (_04858_, _04857_, \oc8051_golden_model_1.TH0 [7]);
  nor (_04859_, _02893_, _02679_);
  and (_04860_, _04859_, _04840_);
  and (_04861_, _04860_, _04720_);
  and (_04862_, _04861_, \oc8051_golden_model_1.TL1 [7]);
  nor (_04863_, _04862_, _04858_);
  and (_04864_, _04840_, _04721_);
  and (_04865_, _04864_, \oc8051_golden_model_1.TCON [7]);
  not (_04866_, _02494_);
  and (_04867_, _04866_, _02324_);
  and (_04868_, _04860_, _04867_);
  and (_04869_, _04868_, \oc8051_golden_model_1.PCON [7]);
  nor (_04870_, _04869_, _04865_);
  and (_04871_, _04870_, _04863_);
  and (_04872_, _04851_, _04847_);
  and (_04873_, _04872_, \oc8051_golden_model_1.DPL [7]);
  not (_04874_, _04873_);
  and (_04875_, _04840_, _04821_);
  and (_04876_, _04875_, \oc8051_golden_model_1.P0INREG [7]);
  not (_04877_, _04876_);
  and (_04878_, _04821_, _04816_);
  and (_04879_, _04878_, _04753_);
  nand (_04880_, _04879_, \oc8051_golden_model_1.P3INREG [7]);
  and (_04881_, _04832_, _04753_);
  and (_04882_, _04881_, _04821_);
  and (_04883_, _04882_, \oc8051_golden_model_1.P1INREG [7]);
  and (_04884_, _04828_, _04753_);
  and (_04885_, _04884_, _04821_);
  and (_04886_, _04885_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_04887_, _04886_, _04883_);
  and (_04888_, _04887_, _04880_);
  and (_04889_, _04888_, _04877_);
  and (_04890_, _04889_, _04874_);
  and (_04891_, _04884_, _04721_);
  and (_04892_, _04891_, \oc8051_golden_model_1.IE [7]);
  and (_04893_, _04838_, _04720_);
  and (_04894_, _04893_, _04881_);
  and (_04895_, _04894_, \oc8051_golden_model_1.SBUF [7]);
  and (_04896_, _04881_, _04721_);
  and (_04897_, _04896_, \oc8051_golden_model_1.SCON [7]);
  or (_04898_, _04897_, _04895_);
  nor (_04899_, _04898_, _04892_);
  and (_04900_, _04848_, _04838_);
  and (_04901_, _04900_, \oc8051_golden_model_1.TMOD [7]);
  and (_04902_, _04860_, _04820_);
  and (_04903_, _04902_, \oc8051_golden_model_1.DPH [7]);
  nor (_04904_, _04903_, _04901_);
  and (_04905_, _04904_, _04899_);
  and (_04906_, _04905_, _04890_);
  and (_04907_, _04906_, _04871_);
  and (_04908_, _04907_, _04856_);
  not (_04909_, _04908_);
  nor (_04910_, _04909_, _04717_);
  nor (_04911_, _04910_, _02039_);
  not (_04912_, _02684_);
  nor (_04913_, _03352_, _03344_);
  and (_04914_, _04913_, _04912_);
  and (_04915_, _02138_, _01717_);
  nor (_04916_, _02236_, _02132_);
  nor (_04917_, _04916_, _03333_);
  nor (_04918_, _04917_, _04915_);
  and (_04919_, _04918_, _04914_);
  not (_04920_, _04919_);
  or (_04921_, _04920_, _04911_);
  or (_04922_, _04921_, _04715_);
  or (_04923_, _04919_, _01952_);
  and (_04924_, _04923_, _04922_);
  or (_04925_, _04924_, _01996_);
  and (_04926_, _04925_, _04459_);
  or (_04927_, _04926_, _01718_);
  and (_04928_, _04544_, _01718_);
  nor (_04929_, _04928_, _03060_);
  and (_04930_, _04929_, _04927_);
  nor (_04931_, _04458_, _03902_);
  and (_04932_, _04458_, _03902_);
  nor (_04933_, _04932_, _04931_);
  nor (_04934_, _04933_, _03062_);
  nor (_04935_, _04934_, _03063_);
  or (_04936_, _04935_, _04930_);
  not (_04937_, _03064_);
  not (_04938_, _03062_);
  not (_04939_, \oc8051_golden_model_1.ACC [7]);
  and (_04940_, _03902_, _04939_);
  nor (_04941_, _03902_, _04939_);
  nor (_04942_, _04941_, _04940_);
  or (_04943_, _04942_, _04938_);
  and (_04944_, _04943_, _04937_);
  and (_04945_, _04944_, _04936_);
  and (_04946_, _04931_, _03064_);
  or (_04947_, _04946_, _03066_);
  or (_04948_, _04947_, _04945_);
  not (_04949_, _03066_);
  or (_04950_, _04941_, _04949_);
  and (_04951_, _04950_, _04948_);
  or (_04952_, _04951_, _01728_);
  not (_04953_, _02202_);
  nor (_04954_, _04953_, _01952_);
  and (_04955_, _04544_, _01728_);
  nor (_04956_, _04955_, _04954_);
  and (_04957_, _04956_, _04952_);
  not (_04958_, _02334_);
  nor (_04959_, _04958_, _01952_);
  not (_04960_, _04954_);
  nor (_04961_, _04932_, _04960_);
  or (_04962_, _04961_, _04959_);
  or (_04963_, _04962_, _04957_);
  not (_04964_, _01726_);
  nand (_04965_, _04940_, _04959_);
  and (_04966_, _04965_, _04964_);
  and (_04967_, _04966_, _04963_);
  nand (_04968_, _04543_, _01726_);
  not (_04969_, _01566_);
  nor (_04970_, _02141_, _04969_);
  not (_04971_, _04970_);
  nor (_04972_, _02930_, _02767_);
  and (_04973_, _04972_, _04971_);
  nand (_04974_, _04973_, _04968_);
  or (_04975_, _04974_, _04967_);
  or (_04976_, _04973_, _04532_);
  and (_04977_, _04976_, _03275_);
  and (_04978_, _04977_, _04975_);
  not (_04979_, _03275_);
  and (_04980_, _04532_, _04979_);
  or (_04981_, _04980_, _03084_);
  or (_04982_, _04981_, _04978_);
  not (_04983_, _03083_);
  not (_04984_, _03084_);
  or (_04985_, _04588_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_04986_, _04590_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_04987_, _04986_, _04581_);
  and (_04988_, _04987_, _04985_);
  or (_04989_, _04590_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_04990_, _04588_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_04991_, _04990_, _04595_);
  and (_04992_, _04991_, _04989_);
  nor (_04993_, _04992_, _04988_);
  nand (_04994_, _04993_, _04574_);
  or (_04995_, _04588_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_04996_, _04590_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_04997_, _04996_, _04581_);
  and (_04998_, _04997_, _04995_);
  or (_04999_, _04590_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_05000_, _04588_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_05001_, _05000_, _04595_);
  and (_05002_, _05001_, _04999_);
  nor (_05003_, _05002_, _04998_);
  nand (_05004_, _05003_, _04601_);
  nand (_05005_, _05004_, _04994_);
  nand (_05006_, _05005_, _04565_);
  or (_05007_, _04590_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_05008_, _04588_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_05009_, _05008_, _05007_);
  nand (_05010_, _05009_, _04581_);
  or (_05011_, _04590_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_05012_, _04588_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05013_, _05012_, _05011_);
  nand (_05014_, _05013_, _04595_);
  nand (_05015_, _05014_, _05010_);
  nand (_05016_, _05015_, _04574_);
  or (_05017_, _04590_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_05018_, _04588_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_05019_, _05018_, _05017_);
  nand (_05020_, _05019_, _04581_);
  or (_05021_, _04590_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_05022_, _04588_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_05023_, _05022_, _05021_);
  nand (_05024_, _05023_, _04595_);
  nand (_05025_, _05024_, _05020_);
  nand (_05026_, _05025_, _04601_);
  nand (_05027_, _05026_, _05016_);
  nand (_05028_, _05027_, _04614_);
  and (_05029_, _05028_, _05006_);
  not (_05030_, _05029_);
  or (_05031_, _04588_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_05032_, _04590_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_05033_, _05032_, _04581_);
  and (_05034_, _05033_, _05031_);
  or (_05035_, _04590_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_05036_, _04588_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_05037_, _05036_, _04595_);
  and (_05038_, _05037_, _05035_);
  nor (_05039_, _05038_, _05034_);
  nand (_05040_, _05039_, _04574_);
  or (_05041_, _04588_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_05042_, _04590_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_05043_, _05042_, _04581_);
  and (_05044_, _05043_, _05041_);
  or (_05045_, _04590_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_05046_, _04588_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_05047_, _05046_, _04595_);
  and (_05048_, _05047_, _05045_);
  nor (_05049_, _05048_, _05044_);
  nand (_05050_, _05049_, _04601_);
  nand (_05051_, _05050_, _05040_);
  nand (_05052_, _05051_, _04565_);
  or (_05053_, _04590_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_05054_, _04588_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_05055_, _05054_, _05053_);
  nand (_05056_, _05055_, _04581_);
  or (_05057_, _04590_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_05058_, _04588_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_05059_, _05058_, _05057_);
  nand (_05060_, _05059_, _04595_);
  nand (_05061_, _05060_, _05056_);
  nand (_05062_, _05061_, _04574_);
  or (_05063_, _04590_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_05064_, _04588_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_05065_, _05064_, _05063_);
  nand (_05066_, _05065_, _04581_);
  or (_05067_, _04590_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_05068_, _04588_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_05069_, _05068_, _05067_);
  nand (_05070_, _05069_, _04595_);
  nand (_05071_, _05070_, _05066_);
  nand (_05072_, _05071_, _04601_);
  nand (_05073_, _05072_, _05062_);
  nand (_05074_, _05073_, _04614_);
  and (_05075_, _05074_, _05052_);
  or (_05076_, _04588_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_05077_, _04590_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_05078_, _05077_, _04581_);
  and (_05079_, _05078_, _05076_);
  or (_05080_, _04590_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_05081_, _04588_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_05082_, _05081_, _04595_);
  and (_05083_, _05082_, _05080_);
  nor (_05084_, _05083_, _05079_);
  nand (_05085_, _05084_, _04574_);
  or (_05086_, _04588_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_05087_, _04590_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_05088_, _05087_, _04581_);
  and (_05089_, _05088_, _05086_);
  or (_05090_, _04590_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_05091_, _04588_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_05092_, _05091_, _04595_);
  and (_05093_, _05092_, _05090_);
  nor (_05094_, _05093_, _05089_);
  nand (_05095_, _05094_, _04601_);
  nand (_05096_, _05095_, _05085_);
  nand (_05097_, _05096_, _04565_);
  or (_05098_, _04590_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_05099_, _04588_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_05100_, _05099_, _05098_);
  nand (_05101_, _05100_, _04581_);
  or (_05102_, _04590_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_05103_, _04588_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_05104_, _05103_, _05102_);
  nand (_05105_, _05104_, _04595_);
  nand (_05106_, _05105_, _05101_);
  nand (_05107_, _05106_, _04574_);
  or (_05108_, _04590_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_05109_, _04588_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_05110_, _05109_, _05108_);
  nand (_05111_, _05110_, _04581_);
  or (_05112_, _04590_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_05113_, _04588_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_05114_, _05113_, _05112_);
  nand (_05115_, _05114_, _04595_);
  nand (_05116_, _05115_, _05111_);
  nand (_05117_, _05116_, _04601_);
  nand (_05118_, _05117_, _05107_);
  nand (_05119_, _05118_, _04614_);
  and (_05120_, _05119_, _05097_);
  nor (_05121_, _05120_, _05075_);
  or (_05122_, _04588_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_05123_, _04590_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_05124_, _05123_, _04581_);
  and (_05125_, _05124_, _05122_);
  or (_05126_, _04590_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_05127_, _04588_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_05128_, _05127_, _04595_);
  and (_05129_, _05128_, _05126_);
  nor (_05130_, _05129_, _05125_);
  nand (_05131_, _05130_, _04574_);
  or (_05132_, _04588_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_05133_, _04590_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_05134_, _05133_, _04581_);
  and (_05135_, _05134_, _05132_);
  or (_05136_, _04590_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_05137_, _04588_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_05138_, _05137_, _04595_);
  and (_05139_, _05138_, _05136_);
  nor (_05140_, _05139_, _05135_);
  nand (_05141_, _05140_, _04601_);
  nand (_05142_, _05141_, _05131_);
  nand (_05143_, _05142_, _04565_);
  or (_05144_, _04590_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_05145_, _04588_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_05146_, _05145_, _05144_);
  nand (_05147_, _05146_, _04581_);
  or (_05148_, _04590_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_05149_, _04588_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_05150_, _05149_, _05148_);
  nand (_05151_, _05150_, _04595_);
  nand (_05152_, _05151_, _05147_);
  nand (_05153_, _05152_, _04574_);
  or (_05154_, _04590_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_05155_, _04588_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_05156_, _05155_, _05154_);
  nand (_05157_, _05156_, _04581_);
  or (_05158_, _04590_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_05159_, _04588_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_05160_, _05159_, _05158_);
  nand (_05161_, _05160_, _04595_);
  nand (_05162_, _05161_, _05157_);
  nand (_05163_, _05162_, _04601_);
  nand (_05164_, _05163_, _05153_);
  nand (_05165_, _05164_, _04614_);
  and (_05166_, _05165_, _05143_);
  or (_05167_, _04588_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_05168_, _04590_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_05169_, _05168_, _04581_);
  and (_05170_, _05169_, _05167_);
  or (_05171_, _04590_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05172_, _04588_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_05173_, _05172_, _04595_);
  and (_05174_, _05173_, _05171_);
  nor (_05175_, _05174_, _05170_);
  nand (_05176_, _05175_, _04574_);
  or (_05177_, _04588_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_05178_, _04590_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_05179_, _05178_, _04581_);
  and (_05180_, _05179_, _05177_);
  or (_05181_, _04590_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_05182_, _04588_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_05183_, _05182_, _04595_);
  and (_05184_, _05183_, _05181_);
  nor (_05185_, _05184_, _05180_);
  nand (_05186_, _05185_, _04601_);
  nand (_05187_, _05186_, _05176_);
  nand (_05188_, _05187_, _04565_);
  or (_05189_, _04590_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_05190_, _04588_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_05191_, _05190_, _05189_);
  nand (_05192_, _05191_, _04581_);
  or (_05193_, _04590_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_05194_, _04588_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_05195_, _05194_, _05193_);
  nand (_05196_, _05195_, _04595_);
  nand (_05197_, _05196_, _05192_);
  nand (_05198_, _05197_, _04574_);
  or (_05199_, _04590_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_05200_, _04588_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_05201_, _05200_, _05199_);
  nand (_05202_, _05201_, _04581_);
  or (_05203_, _04590_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_05204_, _04588_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_05205_, _05204_, _05203_);
  nand (_05206_, _05205_, _04595_);
  nand (_05207_, _05206_, _05202_);
  nand (_05208_, _05207_, _04601_);
  nand (_05209_, _05208_, _05198_);
  nand (_05210_, _05209_, _04614_);
  and (_05211_, _05210_, _05188_);
  nor (_05212_, _05211_, _05166_);
  and (_05213_, _05212_, _05121_);
  or (_05214_, _04588_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05215_, _04590_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_05216_, _05215_, _04581_);
  and (_05217_, _05216_, _05214_);
  or (_05218_, _04590_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05219_, _04588_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_05220_, _05219_, _04595_);
  and (_05221_, _05220_, _05218_);
  nor (_05222_, _05221_, _05217_);
  nand (_05223_, _05222_, _04574_);
  or (_05224_, _04588_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_05225_, _04590_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_05226_, _05225_, _04581_);
  and (_05227_, _05226_, _05224_);
  or (_05228_, _04590_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_05229_, _04588_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_05230_, _05229_, _04595_);
  and (_05231_, _05230_, _05228_);
  nor (_05232_, _05231_, _05227_);
  nand (_05233_, _05232_, _04601_);
  nand (_05234_, _05233_, _05223_);
  nand (_05235_, _05234_, _04565_);
  or (_05236_, _04590_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_05237_, _04588_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_05238_, _05237_, _05236_);
  nand (_05239_, _05238_, _04581_);
  or (_05240_, _04590_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_05241_, _04588_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_05242_, _05241_, _05240_);
  nand (_05243_, _05242_, _04595_);
  nand (_05244_, _05243_, _05239_);
  nand (_05245_, _05244_, _04574_);
  or (_05246_, _04590_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_05247_, _04588_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_05248_, _05247_, _05246_);
  nand (_05249_, _05248_, _04581_);
  or (_05250_, _04590_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_05251_, _04588_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_05252_, _05251_, _05250_);
  nand (_05253_, _05252_, _04595_);
  nand (_05254_, _05253_, _05249_);
  nand (_05255_, _05254_, _04601_);
  nand (_05256_, _05255_, _05245_);
  nand (_05257_, _05256_, _04614_);
  and (_05258_, _05257_, _05235_);
  or (_05259_, _04588_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05260_, _04590_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_05261_, _05260_, _04581_);
  and (_05262_, _05261_, _05259_);
  or (_05263_, _04590_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05264_, _04588_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_05265_, _05264_, _04595_);
  and (_05266_, _05265_, _05263_);
  nor (_05267_, _05266_, _05262_);
  nand (_05268_, _05267_, _04574_);
  or (_05269_, _04588_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05270_, _04590_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_05271_, _05270_, _04581_);
  and (_05272_, _05271_, _05269_);
  or (_05273_, _04590_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05274_, _04588_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_05275_, _05274_, _04595_);
  and (_05276_, _05275_, _05273_);
  nor (_05277_, _05276_, _05272_);
  nand (_05278_, _05277_, _04601_);
  nand (_05279_, _05278_, _05268_);
  nand (_05280_, _05279_, _04565_);
  or (_05281_, _04590_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_05282_, _04588_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_05283_, _05282_, _05281_);
  nand (_05284_, _05283_, _04581_);
  or (_05285_, _04590_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05286_, _04588_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_05287_, _05286_, _05285_);
  nand (_05288_, _05287_, _04595_);
  nand (_05289_, _05288_, _05284_);
  nand (_05290_, _05289_, _04574_);
  or (_05291_, _04590_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_05292_, _04588_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_05293_, _05292_, _05291_);
  nand (_05294_, _05293_, _04581_);
  or (_05295_, _04590_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05296_, _04588_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_05297_, _05296_, _05295_);
  nand (_05298_, _05297_, _04595_);
  nand (_05299_, _05298_, _05294_);
  nand (_05300_, _05299_, _04601_);
  nand (_05301_, _05300_, _05290_);
  nand (_05302_, _05301_, _04614_);
  and (_05303_, _05302_, _05280_);
  nor (_05304_, _05303_, _05258_);
  and (_05305_, _05304_, _05213_);
  and (_05306_, _05305_, _05030_);
  nor (_05307_, _05306_, _04698_);
  and (_05308_, _05306_, _04698_);
  or (_05309_, _05308_, _05307_);
  or (_05310_, _05309_, _04984_);
  and (_05311_, _05310_, _04983_);
  and (_05312_, _05311_, _04982_);
  and (_05313_, _04650_, _03083_);
  or (_05314_, _05313_, _01989_);
  or (_05315_, _05314_, _05312_);
  and (_05316_, _01443_, \oc8051_golden_model_1.PC [2]);
  and (_05317_, _05316_, \oc8051_golden_model_1.PC [3]);
  and (_05318_, _05317_, _04539_);
  nor (_05319_, _05318_, \oc8051_golden_model_1.PC [7]);
  and (_05320_, _04539_, \oc8051_golden_model_1.PC [7]);
  and (_05321_, _05317_, _05320_);
  nor (_05322_, _05321_, _05319_);
  not (_05323_, _05322_);
  nand (_05325_, _05323_, _01989_);
  and (_05326_, _05325_, _05315_);
  or (_05327_, _05326_, _01733_);
  and (_05328_, _04544_, _01733_);
  nor (_05329_, _05328_, _01992_);
  and (_05330_, _05329_, _05327_);
  and (_05331_, _04501_, _01992_);
  not (_05332_, _01631_);
  and (_05333_, _02527_, _05332_);
  not (_05334_, _05333_);
  and (_05335_, _02138_, _01731_);
  nor (_05336_, _02925_, _05335_);
  and (_05337_, _05336_, _05334_);
  not (_05338_, _05337_);
  nor (_05339_, _05338_, _05331_);
  not (_05340_, _05339_);
  nor (_05341_, _05340_, _05330_);
  not (_05342_, _04057_);
  not (_05343_, _04372_);
  nor (_05344_, _03161_, _03020_);
  nor (_05345_, _03624_, _03434_);
  and (_05346_, _05345_, _05344_);
  and (_05347_, _05346_, _05343_);
  and (_05348_, _05347_, _05342_);
  and (_05349_, _03964_, _03796_);
  nor (_05350_, _03964_, _03796_);
  nor (_05351_, _05350_, _05349_);
  and (_05352_, _05351_, _05348_);
  nor (_05353_, _05348_, _03796_);
  nor (_05354_, _05353_, _05352_);
  and (_05355_, _05354_, _05338_);
  nor (_05356_, _05355_, _03293_);
  not (_05357_, _05356_);
  nor (_05358_, _05357_, _05341_);
  nor (_05359_, _05354_, _03292_);
  nor (_05360_, _05359_, _02785_);
  not (_05361_, _05360_);
  nor (_05362_, _05361_, _05358_);
  not (_05363_, _02785_);
  and (_05364_, _05120_, _05075_);
  and (_05365_, _05211_, _05166_);
  and (_05366_, _05365_, _05364_);
  and (_05367_, _05303_, _05258_);
  and (_05368_, _05367_, _05366_);
  and (_05369_, _05368_, _05029_);
  nor (_05370_, _05369_, _04698_);
  and (_05371_, _05369_, _04698_);
  or (_05372_, _05371_, _05370_);
  nor (_05373_, _05372_, _05363_);
  nor (_05374_, _05373_, _03098_);
  not (_05375_, _05374_);
  nor (_05376_, _05375_, _05362_);
  nor (_05377_, _05376_, _04427_);
  nor (_05378_, _05377_, _03385_);
  or (_05379_, _05378_, _03747_);
  or (_05380_, _03746_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_05381_, _05380_, _05379_);
  not (_05382_, _03105_);
  and (_05383_, _03441_, _01986_);
  and (_05384_, _03440_, _01986_);
  nor (_05385_, _05384_, _03443_);
  nor (_05386_, _05385_, _05383_);
  nor (_05387_, _03559_, _03106_);
  nor (_05388_, _05387_, _05384_);
  and (_05389_, _03313_, _01990_);
  nor (_05390_, _05389_, _03383_);
  and (_05391_, _05390_, _05388_);
  nand (_05392_, _05391_, _05386_);
  or (_05393_, _05392_, _05382_);
  and (_05394_, _05393_, _05381_);
  not (_05395_, _01989_);
  and (_05396_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_05397_, _05396_, \oc8051_golden_model_1.PC [10]);
  and (_05398_, _05397_, _05321_);
  and (_05399_, _05398_, \oc8051_golden_model_1.PC [11]);
  and (_05400_, _05399_, \oc8051_golden_model_1.PC [12]);
  and (_05401_, _05400_, \oc8051_golden_model_1.PC [13]);
  and (_05402_, _05401_, \oc8051_golden_model_1.PC [14]);
  nor (_05403_, _05402_, \oc8051_golden_model_1.PC [15]);
  and (_05404_, _05321_, \oc8051_golden_model_1.PC [8]);
  and (_05405_, _05404_, \oc8051_golden_model_1.PC [9]);
  and (_05406_, _05405_, \oc8051_golden_model_1.PC [10]);
  and (_05407_, _05406_, \oc8051_golden_model_1.PC [11]);
  and (_05408_, _05407_, \oc8051_golden_model_1.PC [12]);
  and (_05409_, _05408_, \oc8051_golden_model_1.PC [13]);
  and (_05410_, _05409_, \oc8051_golden_model_1.PC [14]);
  and (_05411_, _05410_, \oc8051_golden_model_1.PC [15]);
  nor (_05412_, _05411_, _05403_);
  or (_05413_, _05412_, _05395_);
  and (_05414_, _05397_, _04542_);
  and (_05415_, _05414_, \oc8051_golden_model_1.PC [11]);
  and (_05416_, _05415_, \oc8051_golden_model_1.PC [12]);
  and (_05417_, _05416_, \oc8051_golden_model_1.PC [13]);
  and (_05418_, _05417_, \oc8051_golden_model_1.PC [14]);
  nor (_05419_, _05418_, \oc8051_golden_model_1.PC [15]);
  and (_05420_, _04542_, \oc8051_golden_model_1.PC [8]);
  and (_05421_, _05420_, \oc8051_golden_model_1.PC [9]);
  and (_05422_, _05421_, \oc8051_golden_model_1.PC [10]);
  and (_05423_, _05422_, \oc8051_golden_model_1.PC [11]);
  and (_05424_, _05423_, \oc8051_golden_model_1.PC [12]);
  and (_05425_, _05424_, \oc8051_golden_model_1.PC [13]);
  and (_05426_, _05425_, \oc8051_golden_model_1.PC [14]);
  and (_05427_, _05426_, \oc8051_golden_model_1.PC [15]);
  nor (_05428_, _05427_, _05419_);
  or (_05429_, _05428_, _01989_);
  and (_05430_, _05429_, _05413_);
  and (_05431_, _05430_, _05390_);
  nor (_05432_, _05431_, _05393_);
  nor (_38581_, _05432_, _05394_);
  not (_05433_, \oc8051_golden_model_1.B [7]);
  nor (_05434_, _39632_, _05433_);
  nor (_05435_, _03847_, _05433_);
  and (_05436_, _04942_, _03847_);
  or (_05437_, _05436_, _05435_);
  and (_05438_, _05437_, _02331_);
  not (_05439_, _03847_);
  nor (_05440_, _05439_, _03796_);
  or (_05441_, _05440_, _05435_);
  nor (_05442_, _03314_, _02137_);
  nor (_05443_, _05442_, _01772_);
  nor (_05444_, _05443_, _02644_);
  or (_05445_, _05444_, _05441_);
  nor (_05446_, _04478_, _05433_);
  and (_05447_, _04517_, _04478_);
  or (_05448_, _05447_, _05446_);
  and (_05449_, _05448_, _02053_);
  and (_05450_, _04650_, _03847_);
  or (_05451_, _05450_, _05435_);
  and (_05452_, _05451_, _02158_);
  nor (_05453_, _02062_, _05433_);
  and (_05454_, _03847_, \oc8051_golden_model_1.ACC [7]);
  or (_05455_, _05454_, _05435_);
  and (_05456_, _05455_, _02062_);
  or (_05457_, _05456_, _05453_);
  and (_05458_, _05457_, _03006_);
  or (_05459_, _05458_, _02057_);
  or (_05460_, _05459_, _05452_);
  and (_05461_, _04521_, _04478_);
  or (_05462_, _05461_, _05446_);
  or (_05463_, _05462_, _02058_);
  and (_05464_, _05463_, _02519_);
  and (_05465_, _05464_, _05460_);
  and (_05466_, _05441_, _02155_);
  or (_05467_, _05466_, _02153_);
  or (_05468_, _05467_, _05465_);
  or (_05469_, _05455_, _02549_);
  and (_05470_, _05469_, _02054_);
  and (_05471_, _05470_, _05468_);
  or (_05472_, _05471_, _05449_);
  and (_05473_, _05472_, _02047_);
  and (_05474_, _02245_, _02128_);
  or (_05475_, _05446_, _04687_);
  and (_05476_, _05475_, _02046_);
  and (_05477_, _05476_, _05462_);
  or (_05478_, _05477_, _05474_);
  or (_05479_, _05478_, _05473_);
  and (_05480_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_05481_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_05482_, _05481_, _05480_);
  and (_05483_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_05484_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_05485_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_05486_, _05485_, _05484_);
  nor (_05487_, _05486_, _05482_);
  and (_05488_, _05487_, _05483_);
  nor (_05489_, _05488_, _05482_);
  and (_05490_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_05491_, _05490_, _05485_);
  and (_05492_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_05493_, _05492_, _05480_);
  nor (_05494_, _05493_, _05491_);
  not (_05495_, _05494_);
  nor (_05496_, _05495_, _05489_);
  and (_05497_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_05498_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_05499_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_05500_, _05499_, _05498_);
  nor (_05501_, _05499_, _05498_);
  nor (_05502_, _05501_, _05500_);
  and (_05503_, _05502_, _05497_);
  nor (_05504_, _05502_, _05497_);
  nor (_05505_, _05504_, _05503_);
  and (_05506_, _05495_, _05489_);
  nor (_05507_, _05506_, _05496_);
  and (_05508_, _05507_, _05505_);
  nor (_05509_, _05508_, _05496_);
  not (_05510_, _05485_);
  and (_05511_, _05490_, _05510_);
  and (_05512_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_05513_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_05514_, _05513_, _05498_);
  and (_05515_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_05516_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_05517_, _05516_, _05515_);
  nor (_05518_, _05517_, _05514_);
  and (_05519_, _05518_, _05512_);
  nor (_05520_, _05518_, _05512_);
  nor (_05521_, _05520_, _05519_);
  and (_05522_, _05521_, _05511_);
  nor (_05523_, _05521_, _05511_);
  nor (_05524_, _05523_, _05522_);
  not (_05525_, _05524_);
  nor (_05526_, _05525_, _05509_);
  and (_05527_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_05528_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_05529_, _05528_, _05527_);
  nor (_05530_, _05503_, _05500_);
  and (_05531_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_05532_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_05533_, _05532_, _05531_);
  nor (_05534_, _05532_, _05531_);
  nor (_05535_, _05534_, _05533_);
  not (_05536_, _05535_);
  nor (_05537_, _05536_, _05530_);
  and (_05538_, _05536_, _05530_);
  nor (_05539_, _05538_, _05537_);
  and (_05540_, _05539_, _05529_);
  nor (_05541_, _05539_, _05529_);
  nor (_05542_, _05541_, _05540_);
  and (_05543_, _05525_, _05509_);
  nor (_05544_, _05543_, _05526_);
  and (_05545_, _05544_, _05542_);
  nor (_05546_, _05545_, _05526_);
  nor (_05547_, _05519_, _05514_);
  and (_05548_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_05549_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_05550_, _05549_, _05548_);
  nor (_05551_, _05549_, _05548_);
  nor (_05552_, _05551_, _05550_);
  not (_05553_, _05552_);
  nor (_05554_, _05553_, _05547_);
  and (_05555_, _05553_, _05547_);
  nor (_05556_, _05555_, _05554_);
  and (_05557_, _05556_, _05533_);
  nor (_05558_, _05556_, _05533_);
  nor (_05559_, _05558_, _05557_);
  nor (_05560_, _05522_, _05491_);
  and (_05561_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_05562_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_05563_, _05562_, _05513_);
  nor (_05564_, _05562_, _05513_);
  nor (_05565_, _05564_, _05563_);
  and (_05566_, _05565_, _05561_);
  nor (_05567_, _05565_, _05561_);
  nor (_05568_, _05567_, _05566_);
  not (_05569_, _05568_);
  nor (_05570_, _05569_, _05560_);
  and (_05571_, _05569_, _05560_);
  nor (_05572_, _05571_, _05570_);
  and (_05573_, _05572_, _05559_);
  nor (_05574_, _05572_, _05559_);
  nor (_05575_, _05574_, _05573_);
  not (_05576_, _05575_);
  nor (_05577_, _05576_, _05546_);
  nor (_05578_, _05540_, _05537_);
  not (_05579_, _05578_);
  and (_05580_, _05576_, _05546_);
  nor (_05581_, _05580_, _05577_);
  and (_05582_, _05581_, _05579_);
  nor (_05583_, _05582_, _05577_);
  nor (_05584_, _05557_, _05554_);
  not (_05585_, _05584_);
  nor (_05586_, _05573_, _05570_);
  not (_05588_, _05586_);
  and (_05590_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_05592_, _05590_, _05513_);
  and (_05594_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_05596_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_05598_, _05596_, _05594_);
  nor (_05600_, _05598_, _05592_);
  nor (_05602_, _05566_, _05563_);
  and (_05604_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_05606_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_05608_, _05606_, _05604_);
  nor (_05610_, _05606_, _05604_);
  nor (_05612_, _05610_, _05608_);
  not (_05614_, _05612_);
  nor (_05616_, _05614_, _05602_);
  and (_05618_, _05614_, _05602_);
  nor (_05620_, _05618_, _05616_);
  and (_05622_, _05620_, _05550_);
  nor (_05624_, _05620_, _05550_);
  nor (_05626_, _05624_, _05622_);
  and (_05628_, _05626_, _05600_);
  nor (_05630_, _05626_, _05600_);
  nor (_05632_, _05630_, _05628_);
  and (_05634_, _05632_, _05588_);
  nor (_05636_, _05632_, _05588_);
  nor (_05638_, _05636_, _05634_);
  and (_05640_, _05638_, _05585_);
  nor (_05642_, _05638_, _05585_);
  nor (_05644_, _05642_, _05640_);
  not (_05646_, _05644_);
  nor (_05648_, _05646_, _05583_);
  nor (_05649_, _05640_, _05634_);
  nor (_05651_, _05622_, _05616_);
  not (_05652_, _05651_);
  and (_05654_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_05655_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_05657_, _05655_, _05654_);
  nor (_05659_, _05655_, _05654_);
  nor (_05660_, _05659_, _05657_);
  and (_05662_, _05660_, _05592_);
  nor (_05663_, _05660_, _05592_);
  nor (_05665_, _05663_, _05662_);
  and (_05666_, _05665_, _05608_);
  nor (_05668_, _05665_, _05608_);
  nor (_05669_, _05668_, _05666_);
  and (_05671_, _05669_, _05590_);
  nor (_05672_, _05669_, _05590_);
  nor (_05674_, _05672_, _05671_);
  and (_05675_, _05674_, _05628_);
  nor (_05677_, _05674_, _05628_);
  nor (_05678_, _05677_, _05675_);
  and (_05680_, _05678_, _05652_);
  nor (_05682_, _05678_, _05652_);
  nor (_05684_, _05682_, _05680_);
  not (_05686_, _05684_);
  nor (_05688_, _05686_, _05649_);
  and (_05690_, _05686_, _05649_);
  nor (_05692_, _05690_, _05688_);
  and (_05694_, _05692_, _05648_);
  nor (_05696_, _05680_, _05675_);
  nor (_05698_, _05666_, _05662_);
  not (_05700_, _05698_);
  and (_05702_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_05704_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_05706_, _05704_, _05702_);
  nor (_05708_, _05704_, _05702_);
  nor (_05710_, _05708_, _05706_);
  and (_05712_, _05710_, _05657_);
  nor (_05714_, _05710_, _05657_);
  nor (_05716_, _05714_, _05712_);
  and (_05718_, _05716_, _05671_);
  nor (_05720_, _05716_, _05671_);
  nor (_05722_, _05720_, _05718_);
  and (_05724_, _05722_, _05700_);
  nor (_05726_, _05722_, _05700_);
  nor (_05728_, _05726_, _05724_);
  not (_05730_, _05728_);
  nor (_05732_, _05730_, _05696_);
  and (_05734_, _05730_, _05696_);
  nor (_05736_, _05734_, _05732_);
  and (_05738_, _05736_, _05688_);
  nor (_05740_, _05736_, _05688_);
  nor (_05742_, _05740_, _05738_);
  and (_05744_, _05742_, _05694_);
  nor (_05746_, _05742_, _05694_);
  and (_05748_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_05750_, _05748_, _05485_);
  and (_05752_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_05754_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_05756_, _05754_, _05481_);
  nor (_05758_, _05756_, _05750_);
  and (_05760_, _05758_, _05752_);
  nor (_05762_, _05760_, _05750_);
  not (_05764_, _05762_);
  nor (_05766_, _05487_, _05483_);
  nor (_05768_, _05766_, _05488_);
  and (_05770_, _05768_, _05764_);
  and (_05772_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_05774_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_05776_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_05778_, _05776_, _05774_);
  nor (_05780_, _05776_, _05774_);
  nor (_05782_, _05780_, _05778_);
  and (_05784_, _05782_, _05772_);
  nor (_05786_, _05782_, _05772_);
  nor (_05788_, _05786_, _05784_);
  nor (_05790_, _05768_, _05764_);
  nor (_05792_, _05790_, _05770_);
  and (_05794_, _05792_, _05788_);
  nor (_05796_, _05794_, _05770_);
  nor (_05798_, _05507_, _05505_);
  nor (_05800_, _05798_, _05508_);
  not (_05802_, _05800_);
  nor (_05804_, _05802_, _05796_);
  and (_05806_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_05808_, _05806_, _05528_);
  nor (_05810_, _05784_, _05778_);
  nor (_05812_, _05528_, _05527_);
  nor (_05814_, _05812_, _05529_);
  not (_05816_, _05814_);
  nor (_05818_, _05816_, _05810_);
  and (_05820_, _05816_, _05810_);
  nor (_05822_, _05820_, _05818_);
  and (_05824_, _05822_, _05808_);
  nor (_05826_, _05822_, _05808_);
  nor (_05828_, _05826_, _05824_);
  and (_05830_, _05802_, _05796_);
  nor (_05832_, _05830_, _05804_);
  and (_05834_, _05832_, _05828_);
  nor (_05836_, _05834_, _05804_);
  nor (_05838_, _05544_, _05542_);
  nor (_05840_, _05838_, _05545_);
  not (_05842_, _05840_);
  nor (_05844_, _05842_, _05836_);
  nor (_05846_, _05824_, _05818_);
  not (_05848_, _05846_);
  and (_05850_, _05842_, _05836_);
  nor (_05852_, _05850_, _05844_);
  and (_05854_, _05852_, _05848_);
  nor (_05856_, _05854_, _05844_);
  nor (_05858_, _05581_, _05579_);
  nor (_05860_, _05858_, _05582_);
  not (_05862_, _05860_);
  nor (_05864_, _05862_, _05856_);
  and (_05866_, _05646_, _05583_);
  nor (_05868_, _05866_, _05648_);
  and (_05870_, _05868_, _05864_);
  nor (_05872_, _05692_, _05648_);
  nor (_05874_, _05872_, _05694_);
  and (_05876_, _05874_, _05870_);
  and (_05878_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_05880_, _05878_, _05748_);
  and (_05882_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_05884_, _05878_, _05748_);
  nor (_05886_, _05884_, _05880_);
  and (_05888_, _05886_, _05882_);
  nor (_05890_, _05888_, _05880_);
  not (_05892_, _05890_);
  nor (_05894_, _05758_, _05752_);
  nor (_05896_, _05894_, _05760_);
  and (_05898_, _05896_, _05892_);
  and (_05900_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_05902_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_05904_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_05906_, _05904_, _05902_);
  nor (_05908_, _05904_, _05902_);
  nor (_05910_, _05908_, _05906_);
  and (_05912_, _05910_, _05900_);
  nor (_05914_, _05910_, _05900_);
  nor (_05916_, _05914_, _05912_);
  nor (_05918_, _05896_, _05892_);
  nor (_05920_, _05918_, _05898_);
  and (_05922_, _05920_, _05916_);
  nor (_05924_, _05922_, _05898_);
  not (_05926_, _05924_);
  nor (_05928_, _05792_, _05788_);
  nor (_05930_, _05928_, _05794_);
  and (_05932_, _05930_, _05926_);
  nor (_05934_, _05912_, _05906_);
  and (_05936_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_05938_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_05940_, _05938_, _05936_);
  nor (_05942_, _05940_, _05808_);
  not (_05944_, _05942_);
  nor (_05946_, _05944_, _05934_);
  and (_05948_, _05944_, _05934_);
  nor (_05950_, _05948_, _05946_);
  nor (_05952_, _05930_, _05926_);
  nor (_05954_, _05952_, _05932_);
  and (_05956_, _05954_, _05950_);
  nor (_05958_, _05956_, _05932_);
  nor (_05960_, _05832_, _05828_);
  nor (_05962_, _05960_, _05834_);
  not (_05964_, _05962_);
  nor (_05966_, _05964_, _05958_);
  and (_05968_, _05964_, _05958_);
  nor (_05970_, _05968_, _05966_);
  and (_05972_, _05970_, _05946_);
  nor (_05974_, _05972_, _05966_);
  nor (_05976_, _05852_, _05848_);
  nor (_05978_, _05976_, _05854_);
  not (_05980_, _05978_);
  nor (_05982_, _05980_, _05974_);
  and (_05984_, _05862_, _05856_);
  nor (_05985_, _05984_, _05864_);
  and (_05986_, _05985_, _05982_);
  nor (_05987_, _05868_, _05864_);
  nor (_05988_, _05987_, _05870_);
  and (_05989_, _05988_, _05986_);
  nor (_05990_, _05988_, _05986_);
  nor (_05991_, _05990_, _05989_);
  and (_05992_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_05993_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_05994_, _05993_, _05992_);
  and (_05995_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_05996_, _05993_, _05992_);
  nor (_05997_, _05996_, _05994_);
  and (_05998_, _05997_, _05995_);
  nor (_05999_, _05998_, _05994_);
  not (_06000_, _05999_);
  nor (_06001_, _05886_, _05882_);
  nor (_06002_, _06001_, _05888_);
  and (_06003_, _06002_, _06000_);
  and (_06004_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_06005_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_06006_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_06007_, _06006_, _06005_);
  nor (_06008_, _06006_, _06005_);
  nor (_06009_, _06008_, _06007_);
  and (_06010_, _06009_, _06004_);
  nor (_06011_, _06009_, _06004_);
  nor (_06012_, _06011_, _06010_);
  nor (_06013_, _06002_, _06000_);
  nor (_06014_, _06013_, _06003_);
  and (_06015_, _06014_, _06012_);
  nor (_06016_, _06015_, _06003_);
  not (_06017_, _06016_);
  nor (_06018_, _05920_, _05916_);
  nor (_06019_, _06018_, _05922_);
  and (_06020_, _06019_, _06017_);
  not (_06021_, _05806_);
  nor (_06022_, _06010_, _06007_);
  nor (_06023_, _06022_, _06021_);
  and (_06024_, _06022_, _06021_);
  nor (_06025_, _06024_, _06023_);
  nor (_06026_, _06019_, _06017_);
  nor (_06027_, _06026_, _06020_);
  and (_06028_, _06027_, _06025_);
  nor (_06029_, _06028_, _06020_);
  not (_06030_, _06029_);
  nor (_06031_, _05954_, _05950_);
  nor (_06032_, _06031_, _05956_);
  and (_06033_, _06032_, _06030_);
  nor (_06034_, _06032_, _06030_);
  nor (_06035_, _06034_, _06033_);
  and (_06036_, _06035_, _06023_);
  nor (_06037_, _06036_, _06033_);
  nor (_06038_, _05970_, _05946_);
  nor (_06039_, _06038_, _05972_);
  not (_06040_, _06039_);
  nor (_06041_, _06040_, _06037_);
  and (_06042_, _05980_, _05974_);
  nor (_06043_, _06042_, _05982_);
  and (_06044_, _06043_, _06041_);
  nor (_06045_, _05985_, _05982_);
  nor (_06046_, _06045_, _05986_);
  and (_06047_, _06046_, _06044_);
  nor (_06048_, _06046_, _06044_);
  nor (_06049_, _06048_, _06047_);
  and (_06050_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_06051_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_06052_, _06051_, _06050_);
  and (_06053_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06054_, _06051_, _06050_);
  nor (_06055_, _06054_, _06052_);
  and (_06056_, _06055_, _06053_);
  nor (_06057_, _06056_, _06052_);
  not (_06058_, _06057_);
  nor (_06059_, _05997_, _05995_);
  nor (_06060_, _06059_, _05998_);
  and (_06061_, _06060_, _06058_);
  and (_06062_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_06063_, _06062_, _06006_);
  and (_06064_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_06065_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_06066_, _06065_, _06064_);
  nor (_06067_, _06066_, _06063_);
  nor (_06068_, _06060_, _06058_);
  nor (_06069_, _06068_, _06061_);
  and (_06070_, _06069_, _06067_);
  nor (_06071_, _06070_, _06061_);
  not (_06072_, _06071_);
  nor (_06073_, _06014_, _06012_);
  nor (_06074_, _06073_, _06015_);
  and (_06075_, _06074_, _06072_);
  nor (_06076_, _06074_, _06072_);
  nor (_06077_, _06076_, _06075_);
  and (_06078_, _06077_, _06063_);
  nor (_06079_, _06078_, _06075_);
  not (_06080_, _06079_);
  nor (_06081_, _06027_, _06025_);
  nor (_06082_, _06081_, _06028_);
  and (_06083_, _06082_, _06080_);
  nor (_06084_, _06035_, _06023_);
  nor (_06085_, _06084_, _06036_);
  and (_06086_, _06085_, _06083_);
  and (_06087_, _06040_, _06037_);
  nor (_06088_, _06087_, _06041_);
  and (_06089_, _06088_, _06086_);
  nor (_06090_, _06043_, _06041_);
  nor (_06091_, _06090_, _06044_);
  and (_06092_, _06091_, _06089_);
  nor (_06093_, _06091_, _06089_);
  nor (_06094_, _06093_, _06092_);
  and (_06095_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_06096_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_06097_, _06096_, _06095_);
  and (_06098_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_06099_, _06096_, _06095_);
  nor (_06100_, _06099_, _06097_);
  and (_06101_, _06100_, _06098_);
  nor (_06102_, _06101_, _06097_);
  not (_06103_, _06102_);
  nor (_06104_, _06055_, _06053_);
  nor (_06105_, _06104_, _06056_);
  and (_06106_, _06105_, _06103_);
  nor (_06107_, _06105_, _06103_);
  nor (_06108_, _06107_, _06106_);
  and (_06109_, _06108_, _06062_);
  nor (_06110_, _06109_, _06106_);
  not (_06111_, _06110_);
  nor (_06112_, _06069_, _06067_);
  nor (_06113_, _06112_, _06070_);
  and (_06114_, _06113_, _06111_);
  nor (_06115_, _06077_, _06063_);
  nor (_06116_, _06115_, _06078_);
  and (_06117_, _06116_, _06114_);
  nor (_06118_, _06082_, _06080_);
  nor (_06119_, _06118_, _06083_);
  and (_06120_, _06119_, _06117_);
  nor (_06121_, _06085_, _06083_);
  nor (_06122_, _06121_, _06086_);
  and (_06123_, _06122_, _06120_);
  nor (_06124_, _06088_, _06086_);
  nor (_06125_, _06124_, _06089_);
  and (_06126_, _06125_, _06123_);
  and (_06127_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_06128_, _06127_, _06096_);
  nor (_06129_, _06100_, _06098_);
  nor (_06130_, _06129_, _06101_);
  and (_06131_, _06130_, _06128_);
  nor (_06132_, _06108_, _06062_);
  nor (_06133_, _06132_, _06109_);
  and (_06134_, _06133_, _06131_);
  nor (_06135_, _06113_, _06111_);
  nor (_06136_, _06135_, _06114_);
  and (_06137_, _06136_, _06134_);
  nor (_06138_, _06116_, _06114_);
  nor (_06139_, _06138_, _06117_);
  and (_06140_, _06139_, _06137_);
  nor (_06141_, _06119_, _06117_);
  nor (_06142_, _06141_, _06120_);
  and (_06143_, _06142_, _06140_);
  nor (_06144_, _06122_, _06120_);
  nor (_06145_, _06144_, _06123_);
  and (_06146_, _06145_, _06143_);
  nor (_06147_, _06125_, _06123_);
  nor (_06148_, _06147_, _06126_);
  and (_06149_, _06148_, _06146_);
  nor (_06150_, _06149_, _06126_);
  not (_06151_, _06150_);
  and (_06152_, _06151_, _06094_);
  nor (_06153_, _06152_, _06092_);
  not (_06154_, _06153_);
  and (_06155_, _06154_, _06049_);
  nor (_06156_, _06155_, _06047_);
  not (_06157_, _06156_);
  and (_06158_, _06157_, _05991_);
  nor (_06159_, _06158_, _05989_);
  not (_06160_, _06159_);
  nor (_06161_, _05874_, _05870_);
  nor (_06162_, _06161_, _05876_);
  and (_06163_, _06162_, _06160_);
  nor (_06164_, _06163_, _05876_);
  nor (_06165_, _06164_, _05746_);
  or (_06166_, _06165_, _05744_);
  and (_06167_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_06168_, _06167_);
  nor (_06169_, _06168_, _05655_);
  nor (_06170_, _06169_, _05712_);
  nor (_06171_, _05724_, _05718_);
  nor (_06172_, _06171_, _06170_);
  and (_06173_, _06171_, _06170_);
  nor (_06174_, _06173_, _06172_);
  not (_06175_, _06174_);
  nor (_06176_, _05738_, _05732_);
  and (_06177_, _06176_, _06175_);
  nor (_06178_, _06176_, _06175_);
  nor (_06179_, _06178_, _06177_);
  and (_06180_, _06179_, _06166_);
  not (_06181_, _05474_);
  or (_06182_, _05706_, _06181_);
  or (_06183_, _06182_, _06172_);
  or (_06184_, _06183_, _06178_);
  or (_06185_, _06184_, _06180_);
  and (_06186_, _06185_, _02043_);
  and (_06187_, _06186_, _05479_);
  not (_06188_, _05444_);
  not (_06189_, _04478_);
  nor (_06190_, _04503_, _06189_);
  or (_06191_, _06190_, _05446_);
  and (_06192_, _06191_, _02042_);
  or (_06193_, _06192_, _06188_);
  or (_06194_, _06193_, _06187_);
  and (_06195_, _06194_, _05445_);
  or (_06196_, _06195_, _02031_);
  and (_06197_, _04637_, _03847_);
  or (_06198_, _05435_, _02032_);
  or (_06199_, _06198_, _06197_);
  and (_06200_, _06199_, _02037_);
  and (_06201_, _06200_, _06196_);
  and (_06202_, _02245_, _01710_);
  nor (_06203_, _04910_, _05439_);
  or (_06204_, _06203_, _05435_);
  and (_06205_, _06204_, _01765_);
  or (_06206_, _06205_, _06202_);
  or (_06207_, _06206_, _06201_);
  not (_06208_, \oc8051_golden_model_1.B [1]);
  nor (_06209_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_06210_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_06211_, _06210_, _06209_);
  and (_06212_, _06211_, _06208_);
  nor (_06213_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not (_06214_, \oc8051_golden_model_1.B [0]);
  and (_06215_, _06214_, \oc8051_golden_model_1.ACC [7]);
  and (_06216_, _06215_, _06213_);
  and (_06217_, _06216_, _06212_);
  or (_06218_, _06214_, \oc8051_golden_model_1.ACC [7]);
  and (_06219_, _06218_, _06213_);
  and (_06220_, _06219_, _06212_);
  or (_06221_, _06220_, _04939_);
  not (_06222_, \oc8051_golden_model_1.B [2]);
  not (_06223_, \oc8051_golden_model_1.B [3]);
  not (_06224_, \oc8051_golden_model_1.B [4]);
  not (_06225_, \oc8051_golden_model_1.B [5]);
  nor (_06226_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_06227_, _06226_, _06225_);
  and (_06228_, _06227_, _06224_);
  and (_06229_, _06228_, _06223_);
  and (_06230_, _06229_, _06222_);
  not (_06231_, \oc8051_golden_model_1.ACC [6]);
  and (_06232_, \oc8051_golden_model_1.B [0], _06231_);
  nor (_06233_, _06232_, _04939_);
  nor (_06234_, _06233_, _06208_);
  not (_06235_, _06234_);
  and (_06236_, _06235_, _06230_);
  nor (_06237_, _06236_, _06221_);
  nor (_06238_, _06237_, _06217_);
  and (_06239_, _06236_, \oc8051_golden_model_1.B [0]);
  nor (_06240_, _06239_, _06231_);
  and (_06241_, _06240_, _06208_);
  nor (_06242_, _06240_, _06208_);
  nor (_06243_, _06242_, _06241_);
  nor (_06244_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_06245_, _06244_, _05748_);
  nor (_06246_, _06245_, \oc8051_golden_model_1.ACC [4]);
  nor (_06247_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_06248_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_06249_, _06248_, _06214_);
  nor (_06250_, _06249_, _06247_);
  nor (_06251_, _06250_, _06246_);
  not (_06252_, _06251_);
  and (_06253_, _06252_, _06243_);
  nor (_06254_, _06238_, \oc8051_golden_model_1.B [2]);
  nor (_06255_, _06254_, _06241_);
  not (_06256_, _06255_);
  nor (_06257_, _06256_, _06253_);
  and (_06258_, \oc8051_golden_model_1.B [2], _04939_);
  nor (_06259_, _06258_, \oc8051_golden_model_1.B [7]);
  and (_06260_, _06259_, _06211_);
  not (_06261_, _06260_);
  nor (_06262_, _06261_, _06257_);
  nor (_06263_, _06262_, _06238_);
  nor (_06264_, _06263_, _06217_);
  and (_06265_, _06228_, \oc8051_golden_model_1.ACC [7]);
  nor (_06266_, _06265_, _06229_);
  nor (_06267_, _06252_, _06243_);
  nor (_06268_, _06267_, _06253_);
  not (_06269_, _06268_);
  and (_06270_, _06269_, _06262_);
  nor (_06271_, _06262_, _06240_);
  nor (_06272_, _06271_, _06270_);
  and (_06273_, _06272_, _06222_);
  nor (_06274_, _06272_, _06222_);
  nor (_06275_, _06274_, _06273_);
  not (_06276_, _06275_);
  not (_06277_, \oc8051_golden_model_1.ACC [5]);
  nor (_06278_, _06262_, _06277_);
  and (_06279_, _06262_, _06245_);
  or (_06280_, _06279_, _06278_);
  and (_06281_, _06280_, _06208_);
  nor (_06282_, _06280_, _06208_);
  not (_06283_, \oc8051_golden_model_1.ACC [4]);
  and (_06284_, \oc8051_golden_model_1.B [0], _06283_);
  nor (_06285_, _06284_, _06282_);
  nor (_06286_, _06285_, _06281_);
  nor (_06287_, _06286_, _06276_);
  nor (_06288_, _06264_, \oc8051_golden_model_1.B [3]);
  nor (_06289_, _06288_, _06273_);
  not (_06290_, _06289_);
  nor (_06291_, _06290_, _06287_);
  nor (_06292_, _06291_, _06266_);
  nor (_06293_, _06292_, _06264_);
  nor (_06294_, _06293_, _06217_);
  not (_06295_, _06292_);
  and (_06296_, _06286_, _06276_);
  nor (_06297_, _06296_, _06287_);
  nor (_06298_, _06297_, _06295_);
  nor (_06299_, _06292_, _06272_);
  nor (_06300_, _06299_, _06298_);
  and (_06301_, _06300_, _06223_);
  nor (_06302_, _06300_, _06223_);
  nor (_06303_, _06302_, _06301_);
  not (_06304_, _06303_);
  nor (_06305_, _06292_, _06280_);
  nor (_06306_, _06282_, _06281_);
  and (_06307_, _06306_, _06284_);
  nor (_06308_, _06306_, _06284_);
  nor (_06309_, _06308_, _06307_);
  and (_06310_, _06309_, _06292_);
  or (_06311_, _06310_, _06305_);
  nor (_06312_, _06311_, \oc8051_golden_model_1.B [2]);
  and (_06313_, _06311_, \oc8051_golden_model_1.B [2]);
  nor (_06314_, _06292_, _06283_);
  nor (_06315_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_06316_, _06315_, _05992_);
  and (_06317_, _06292_, _06316_);
  or (_06318_, _06317_, _06314_);
  and (_06319_, _06318_, _06208_);
  nor (_06320_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_06321_, _06320_, _06050_);
  nor (_06322_, _06321_, \oc8051_golden_model_1.ACC [2]);
  nor (_06323_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_06324_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_06325_, _06324_, _06214_);
  nor (_06326_, _06325_, _06323_);
  nor (_06327_, _06326_, _06322_);
  not (_06328_, _06327_);
  nor (_06329_, _06318_, _06208_);
  nor (_06330_, _06329_, _06319_);
  and (_06331_, _06330_, _06328_);
  nor (_06332_, _06331_, _06319_);
  nor (_06333_, _06332_, _06313_);
  nor (_06334_, _06333_, _06312_);
  nor (_06335_, _06334_, _06304_);
  nor (_06336_, _06294_, \oc8051_golden_model_1.B [4]);
  nor (_06337_, _06336_, _06301_);
  not (_06338_, _06337_);
  nor (_06339_, _06338_, _06335_);
  not (_06340_, _06227_);
  and (_06341_, \oc8051_golden_model_1.B [4], _04939_);
  nor (_06342_, _06341_, _06340_);
  not (_06343_, _06342_);
  nor (_06344_, _06343_, _06339_);
  nor (_06345_, _06344_, _06294_);
  nor (_06346_, _06345_, _06217_);
  and (_06347_, _06226_, \oc8051_golden_model_1.ACC [7]);
  nor (_06348_, _06347_, _06227_);
  nor (_06349_, _06346_, \oc8051_golden_model_1.B [5]);
  and (_06350_, _06334_, _06304_);
  nor (_06351_, _06350_, _06335_);
  not (_06352_, _06351_);
  and (_06353_, _06352_, _06344_);
  nor (_06354_, _06344_, _06300_);
  nor (_06355_, _06354_, _06353_);
  and (_06356_, _06355_, _06224_);
  nor (_06357_, _06355_, _06224_);
  nor (_06358_, _06357_, _06356_);
  not (_06359_, _06358_);
  nor (_06360_, _06344_, _06311_);
  nor (_06361_, _06313_, _06312_);
  and (_06362_, _06361_, _06332_);
  nor (_06363_, _06361_, _06332_);
  nor (_06364_, _06363_, _06362_);
  not (_06365_, _06364_);
  and (_06366_, _06365_, _06344_);
  nor (_06367_, _06366_, _06360_);
  nor (_06368_, _06367_, \oc8051_golden_model_1.B [3]);
  and (_06369_, _06367_, \oc8051_golden_model_1.B [3]);
  nor (_06370_, _06330_, _06328_);
  nor (_06371_, _06370_, _06331_);
  not (_06372_, _06371_);
  and (_06373_, _06372_, _06344_);
  nor (_06374_, _06344_, _06318_);
  nor (_06375_, _06374_, _06373_);
  and (_06376_, _06375_, _06222_);
  not (_06377_, \oc8051_golden_model_1.ACC [3]);
  nor (_06378_, _06344_, _06377_);
  and (_06379_, _06344_, _06321_);
  or (_06380_, _06379_, _06378_);
  and (_06381_, _06380_, _06208_);
  nor (_06382_, _06380_, _06208_);
  not (_06383_, \oc8051_golden_model_1.ACC [2]);
  and (_06384_, \oc8051_golden_model_1.B [0], _06383_);
  nor (_06385_, _06384_, _06382_);
  nor (_06386_, _06385_, _06381_);
  nor (_06387_, _06375_, _06222_);
  nor (_06389_, _06387_, _06376_);
  not (_06390_, _06389_);
  nor (_06391_, _06390_, _06386_);
  nor (_06392_, _06391_, _06376_);
  nor (_06393_, _06392_, _06369_);
  nor (_06394_, _06393_, _06368_);
  nor (_06395_, _06394_, _06359_);
  or (_06396_, _06395_, _06356_);
  nor (_06397_, _06396_, _06349_);
  nor (_06398_, _06397_, _06348_);
  nor (_06400_, _06398_, _06346_);
  not (_06401_, _06398_);
  and (_06402_, _06394_, _06359_);
  nor (_06403_, _06402_, _06395_);
  nor (_06404_, _06403_, _06401_);
  nor (_06405_, _06398_, _06355_);
  nor (_06406_, _06405_, _06404_);
  and (_06407_, _06406_, _06225_);
  nor (_06408_, _06406_, _06225_);
  nor (_06409_, _06408_, _06407_);
  not (_06411_, _06409_);
  nor (_06412_, _06398_, _06367_);
  nor (_06413_, _06369_, _06368_);
  nor (_06414_, _06413_, _06392_);
  and (_06415_, _06413_, _06392_);
  or (_06416_, _06415_, _06414_);
  and (_06417_, _06416_, _06398_);
  or (_06418_, _06417_, _06412_);
  and (_06419_, _06418_, _06224_);
  nor (_06420_, _06418_, _06224_);
  and (_06422_, _06390_, _06386_);
  nor (_06423_, _06422_, _06391_);
  nor (_06424_, _06423_, _06401_);
  nor (_06425_, _06398_, _06375_);
  nor (_06426_, _06425_, _06424_);
  and (_06427_, _06426_, _06223_);
  nor (_06428_, _06382_, _06381_);
  nor (_06429_, _06428_, _06384_);
  and (_06430_, _06428_, _06384_);
  or (_06431_, _06430_, _06429_);
  nor (_06433_, _06431_, _06401_);
  nor (_06434_, _06398_, _06380_);
  nor (_06435_, _06434_, _06433_);
  and (_06436_, _06435_, _06222_);
  nor (_06437_, _06435_, _06222_);
  nor (_06438_, _06398_, _06383_);
  nor (_06439_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_06440_, _06439_, _06095_);
  and (_06441_, _06398_, _06440_);
  or (_06442_, _06441_, _06438_);
  and (_06444_, _06442_, _06208_);
  and (_06445_, \oc8051_golden_model_1.B [0], _01804_);
  not (_06446_, _06445_);
  nor (_06447_, _06442_, _06208_);
  nor (_06448_, _06447_, _06444_);
  and (_06449_, _06448_, _06446_);
  nor (_06450_, _06449_, _06444_);
  nor (_06451_, _06450_, _06437_);
  nor (_06452_, _06451_, _06436_);
  nor (_06453_, _06426_, _06223_);
  nor (_06454_, _06453_, _06427_);
  not (_06455_, _06454_);
  nor (_06456_, _06455_, _06452_);
  nor (_06457_, _06456_, _06427_);
  nor (_06458_, _06457_, _06420_);
  nor (_06459_, _06458_, _06419_);
  nor (_06460_, _06459_, _06411_);
  nor (_06461_, _06460_, _06407_);
  and (_06462_, _05433_, \oc8051_golden_model_1.ACC [7]);
  nor (_06463_, _06462_, _06226_);
  nor (_06464_, _06463_, _06461_);
  not (_06465_, _06226_);
  nor (_06466_, _06400_, _06217_);
  nor (_06467_, _06466_, _06465_);
  nor (_06468_, _06467_, _06464_);
  and (_06469_, _06468_, _06400_);
  nor (_06470_, _06469_, _06217_);
  and (_06471_, _06470_, \oc8051_golden_model_1.B [7]);
  and (_06472_, _06470_, _05433_);
  nor (_06473_, _06472_, _06167_);
  not (_06474_, _06473_);
  not (_06475_, \oc8051_golden_model_1.B [6]);
  and (_06476_, _06459_, _06411_);
  nor (_06477_, _06476_, _06460_);
  nor (_06478_, _06477_, _06468_);
  not (_06479_, _06468_);
  nor (_06480_, _06479_, _06406_);
  nor (_06481_, _06480_, _06478_);
  nor (_06482_, _06481_, _06475_);
  and (_06483_, _06481_, _06475_);
  nor (_06484_, _06420_, _06419_);
  nor (_06485_, _06484_, _06457_);
  and (_06486_, _06484_, _06457_);
  or (_06487_, _06486_, _06485_);
  nor (_06488_, _06487_, _06468_);
  nor (_06489_, _06479_, _06418_);
  nor (_06490_, _06489_, _06488_);
  nor (_06491_, _06490_, _06225_);
  and (_06492_, _06490_, _06225_);
  not (_06493_, _06492_);
  and (_06494_, _06455_, _06452_);
  nor (_06495_, _06494_, _06456_);
  nor (_06496_, _06495_, _06468_);
  nor (_06497_, _06479_, _06426_);
  nor (_06498_, _06497_, _06496_);
  nor (_06499_, _06498_, _06224_);
  and (_06500_, _06468_, _06435_);
  nor (_06501_, _06437_, _06436_);
  and (_06502_, _06501_, _06450_);
  nor (_06503_, _06501_, _06450_);
  nor (_06504_, _06503_, _06502_);
  nor (_06505_, _06504_, _06468_);
  or (_06506_, _06505_, _06500_);
  and (_06507_, _06506_, _06223_);
  nor (_06508_, _06506_, _06223_);
  nor (_06509_, _06508_, _06507_);
  nor (_06510_, _06448_, _06446_);
  nor (_06511_, _06510_, _06449_);
  nor (_06512_, _06511_, _06468_);
  nor (_06513_, _06479_, _06442_);
  nor (_06514_, _06513_, _06512_);
  nor (_06515_, _06514_, _06222_);
  and (_06516_, _06514_, _06222_);
  nor (_06517_, _06516_, _06515_);
  and (_06518_, _06517_, _06509_);
  and (_06519_, _06468_, _01804_);
  and (_06520_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_06521_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_06522_, _06521_, _06520_);
  nor (_06523_, _06468_, _06522_);
  nor (_06524_, _06523_, _06519_);
  and (_06525_, _06524_, _06208_);
  nor (_06526_, _06524_, _06208_);
  and (_06527_, _06214_, \oc8051_golden_model_1.ACC [0]);
  not (_06528_, _06527_);
  nor (_06529_, _06528_, _06526_);
  nor (_06530_, _06529_, _06525_);
  and (_06531_, _06530_, _06518_);
  and (_06532_, _06515_, _06509_);
  nor (_06533_, _06532_, _06508_);
  not (_06534_, _06533_);
  nor (_06535_, _06534_, _06531_);
  and (_06536_, _06498_, _06224_);
  nor (_06537_, _06536_, _06535_);
  or (_06538_, _06537_, _06499_);
  and (_06539_, _06538_, _06493_);
  nor (_06540_, _06539_, _06491_);
  nor (_06541_, _06540_, _06483_);
  or (_06542_, _06541_, _06482_);
  and (_06543_, _06542_, _06474_);
  nor (_06544_, _06543_, _06471_);
  nor (_06545_, _06483_, _06482_);
  and (_06546_, _06545_, _06474_);
  nor (_06547_, _06536_, _06499_);
  nor (_06548_, _06492_, _06491_);
  and (_06549_, _06548_, _06547_);
  and (_06550_, _06549_, _06546_);
  and (_06551_, \oc8051_golden_model_1.B [0], _01887_);
  not (_06552_, _06551_);
  nor (_06553_, _06526_, _06525_);
  and (_06554_, _06553_, _06552_);
  and (_06555_, _06554_, _06528_);
  and (_06556_, _06555_, _06518_);
  and (_06557_, _06556_, _06550_);
  nor (_06558_, _06557_, _06544_);
  and (_06559_, _06558_, _06469_);
  not (_06560_, _06202_);
  or (_06561_, _06217_, _06560_);
  or (_06562_, _06561_, _06559_);
  and (_06563_, _06562_, _01995_);
  and (_06564_, _06563_, _06207_);
  and (_06565_, _04716_, _03847_);
  or (_06566_, _06565_, _05435_);
  and (_06567_, _06566_, _01994_);
  or (_06568_, _06567_, _02210_);
  or (_06569_, _06568_, _06564_);
  and (_06570_, _04933_, _03847_);
  or (_06571_, _05435_, _03059_);
  or (_06572_, _06571_, _06570_);
  and (_06573_, _06572_, _03061_);
  and (_06574_, _06573_, _06569_);
  or (_06575_, _06574_, _05438_);
  and (_06576_, _06575_, _02208_);
  or (_06577_, _05435_, _03903_);
  and (_06578_, _06566_, _02206_);
  and (_06579_, _06578_, _06577_);
  or (_06580_, _06579_, _06576_);
  and (_06581_, _06580_, _03065_);
  and (_06582_, _05455_, _02342_);
  and (_06583_, _06582_, _06577_);
  or (_06584_, _06583_, _02202_);
  or (_06585_, _06584_, _06581_);
  nor (_06586_, _04932_, _05439_);
  or (_06587_, _05435_, _04953_);
  or (_06588_, _06587_, _06586_);
  and (_06589_, _06588_, _04958_);
  and (_06590_, _06589_, _06585_);
  nor (_06591_, _04940_, _05439_);
  or (_06592_, _06591_, _05435_);
  and (_06593_, _06592_, _02334_);
  or (_06594_, _06593_, _02366_);
  or (_06595_, _06594_, _06590_);
  or (_06596_, _05451_, _02778_);
  and (_06597_, _06596_, _01698_);
  and (_06598_, _06597_, _06595_);
  and (_06599_, _05448_, _01697_);
  or (_06600_, _06599_, _02081_);
  or (_06601_, _06600_, _06598_);
  and (_06602_, _04426_, _03847_);
  or (_06603_, _05435_, _02082_);
  or (_06604_, _06603_, _06602_);
  and (_06605_, _06604_, _39632_);
  and (_06606_, _06605_, _06601_);
  or (_06607_, _06606_, _05434_);
  and (_38582_, _06607_, _39026_);
  nor (_06608_, _39632_, _04939_);
  and (_06609_, _02030_, _01737_);
  nor (_06610_, _02141_, _02499_);
  nor (_06611_, _02134_, _02499_);
  or (_06612_, _02914_, _02753_);
  or (_06613_, _06612_, _06611_);
  nor (_06614_, _06613_, _06610_);
  and (_06615_, _03796_, _04939_);
  nor (_06616_, _03796_, _04939_);
  nor (_06617_, _06616_, _06615_);
  nor (_06618_, _03964_, _06231_);
  and (_06619_, _03964_, _06231_);
  nor (_06620_, _06619_, _06618_);
  nor (_06621_, _04057_, _06277_);
  and (_06622_, _04057_, _06277_);
  nor (_06623_, _04372_, _06283_);
  and (_06624_, _04372_, _06283_);
  nor (_06625_, _06624_, _06623_);
  not (_06626_, _06625_);
  nor (_06627_, _03434_, _06377_);
  not (_06628_, _06627_);
  and (_06629_, _03434_, _06377_);
  nor (_06630_, _03624_, _06383_);
  and (_06631_, _03624_, _06383_);
  nor (_06632_, _06631_, _06630_);
  not (_06633_, _06632_);
  nor (_06634_, _03161_, _01804_);
  and (_06635_, _03161_, _01804_);
  nor (_06636_, _06635_, _06634_);
  and (_06637_, _03002_, \oc8051_golden_model_1.ACC [0]);
  and (_06638_, _06637_, _06636_);
  nor (_06639_, _06638_, _06634_);
  nor (_06640_, _06639_, _06633_);
  nor (_06641_, _06640_, _06630_);
  or (_06642_, _06641_, _06629_);
  and (_06643_, _06642_, _06628_);
  nor (_06644_, _06643_, _06626_);
  nor (_06645_, _06644_, _06623_);
  nor (_06646_, _06645_, _06622_);
  or (_06647_, _06646_, _06621_);
  and (_06648_, _06647_, _06620_);
  nor (_06649_, _06648_, _06618_);
  nor (_06650_, _06649_, _06617_);
  and (_06651_, _06649_, _06617_);
  or (_06652_, _06651_, _06650_);
  or (_06653_, _06652_, _06614_);
  and (_06654_, _02030_, _01725_);
  not (_06655_, _03964_);
  and (_06656_, _05348_, \oc8051_golden_model_1.PSW [7]);
  and (_06657_, _06656_, _06655_);
  nor (_06658_, _06657_, _03796_);
  and (_06659_, _06657_, _03796_);
  nor (_06660_, _06659_, _06658_);
  and (_06661_, _06660_, \oc8051_golden_model_1.ACC [7]);
  nor (_06662_, _06660_, \oc8051_golden_model_1.ACC [7]);
  nor (_06663_, _06662_, _06661_);
  nor (_06664_, _06656_, _06655_);
  nor (_06665_, _06664_, _06657_);
  and (_06666_, _06665_, \oc8051_golden_model_1.ACC [6]);
  nor (_06667_, _06665_, _06231_);
  and (_06668_, _06665_, _06231_);
  nor (_06669_, _06668_, _06667_);
  and (_06670_, _05347_, \oc8051_golden_model_1.PSW [7]);
  nor (_06671_, _06670_, _05342_);
  nor (_06672_, _06671_, _06656_);
  and (_06673_, _06672_, \oc8051_golden_model_1.ACC [5]);
  and (_06674_, _06672_, _06277_);
  nor (_06675_, _06672_, _06277_);
  nor (_06676_, _06675_, _06674_);
  and (_06677_, _05344_, \oc8051_golden_model_1.PSW [7]);
  and (_06678_, _06677_, _05345_);
  nor (_06679_, _06678_, _05343_);
  nor (_06680_, _06679_, _06670_);
  and (_06681_, _06680_, \oc8051_golden_model_1.ACC [4]);
  nor (_06682_, _06680_, _06283_);
  and (_06683_, _06680_, _06283_);
  nor (_06684_, _06683_, _06682_);
  not (_06685_, _03434_);
  and (_06686_, _05344_, _03625_);
  and (_06687_, _06686_, \oc8051_golden_model_1.PSW [7]);
  nor (_06688_, _06687_, _06685_);
  nor (_06689_, _06688_, _06678_);
  and (_06690_, _06689_, \oc8051_golden_model_1.ACC [3]);
  nor (_06691_, _06689_, _06377_);
  and (_06692_, _06689_, _06377_);
  nor (_06693_, _06692_, _06691_);
  nor (_06694_, _06677_, _03625_);
  nor (_06695_, _06694_, _06687_);
  and (_06696_, _06695_, \oc8051_golden_model_1.ACC [2]);
  nor (_06697_, _06695_, _06383_);
  and (_06698_, _06695_, _06383_);
  nor (_06699_, _06698_, _06697_);
  and (_06700_, _03002_, \oc8051_golden_model_1.PSW [7]);
  nor (_06701_, _06700_, _03163_);
  nor (_06702_, _06701_, _06677_);
  and (_06703_, _06702_, \oc8051_golden_model_1.ACC [1]);
  and (_06704_, _06702_, _01804_);
  nor (_06705_, _06702_, _01804_);
  nor (_06706_, _06705_, _06704_);
  not (_06707_, \oc8051_golden_model_1.PSW [7]);
  and (_06708_, _03020_, _06707_);
  nor (_06709_, _06708_, _06700_);
  and (_06710_, _06709_, \oc8051_golden_model_1.ACC [0]);
  not (_06711_, _06710_);
  nor (_06712_, _06711_, _06706_);
  nor (_06713_, _06712_, _06703_);
  nor (_06714_, _06713_, _06699_);
  nor (_06715_, _06714_, _06696_);
  nor (_06716_, _06715_, _06693_);
  nor (_06717_, _06716_, _06690_);
  nor (_06718_, _06717_, _06684_);
  nor (_06719_, _06718_, _06681_);
  nor (_06720_, _06719_, _06676_);
  nor (_06721_, _06720_, _06673_);
  nor (_06722_, _06721_, _06669_);
  nor (_06723_, _06722_, _06666_);
  nor (_06724_, _06723_, _06663_);
  and (_06725_, _06723_, _06663_);
  nor (_06726_, _06725_, _06724_);
  and (_06727_, _02132_, _01725_);
  not (_06728_, _06727_);
  or (_06729_, _05442_, _02729_);
  and (_06730_, _06729_, _06728_);
  or (_06731_, _06730_, _06726_);
  and (_06732_, _02137_, _01735_);
  nand (_06733_, _06732_, _06615_);
  and (_06734_, _02245_, _01721_);
  nor (_06735_, _03841_, _04939_);
  not (_06736_, _03841_);
  nor (_06737_, _06736_, _03796_);
  nor (_06738_, _06737_, _06735_);
  nand (_06739_, _06738_, _06188_);
  and (_06740_, _02245_, _01766_);
  not (_06741_, _06740_);
  and (_06742_, _03826_, \oc8051_golden_model_1.PSW [7]);
  and (_06743_, _06742_, _03852_);
  and (_06744_, _06743_, _03818_);
  and (_06745_, _06744_, _03495_);
  nor (_06746_, _06745_, _03835_);
  and (_06747_, _06744_, _02119_);
  nor (_06748_, _06747_, _06746_);
  and (_06749_, _06748_, \oc8051_golden_model_1.ACC [7]);
  nor (_06750_, _06748_, \oc8051_golden_model_1.ACC [7]);
  nor (_06751_, _06750_, _06749_);
  not (_06752_, _06751_);
  nor (_06753_, _06744_, _03495_);
  nor (_06754_, _06753_, _06745_);
  nor (_06755_, _06754_, _06231_);
  and (_06756_, _06754_, _06231_);
  nor (_06757_, _06755_, _06756_);
  and (_06758_, _06743_, _03799_);
  nor (_06759_, _06758_, _03810_);
  nor (_06760_, _06759_, _06744_);
  nor (_06761_, _06760_, _06277_);
  and (_06762_, _06760_, _06277_);
  nor (_06763_, _06762_, _06761_);
  nor (_06764_, _06743_, _03799_);
  nor (_06765_, _06764_, _06758_);
  nor (_06766_, _06765_, _06283_);
  and (_06767_, _06765_, _06283_);
  nor (_06768_, _06767_, _06766_);
  and (_06769_, _06768_, _06763_);
  nor (_06770_, _04502_, _02120_);
  nor (_06771_, _06770_, _06743_);
  nor (_06772_, _06771_, _06377_);
  and (_06773_, _06771_, _06377_);
  nor (_06774_, _06773_, _06772_);
  nor (_06775_, _06742_, _02453_);
  nor (_06776_, _06775_, _04502_);
  nor (_06777_, _06776_, _06383_);
  and (_06778_, _06776_, _06383_);
  nor (_06779_, _06778_, _06777_);
  and (_06780_, _06779_, _06774_);
  nor (_06781_, _02027_, _06707_);
  nor (_06782_, _06781_, _02860_);
  nor (_06783_, _06782_, _06742_);
  nor (_06784_, _06783_, _01804_);
  and (_06785_, _06783_, _01804_);
  nor (_06786_, _06785_, _06784_);
  nor (_06787_, _02027_, \oc8051_golden_model_1.PSW [7]);
  and (_06788_, _02027_, \oc8051_golden_model_1.PSW [7]);
  nor (_06789_, _06788_, _06787_);
  nor (_06790_, _06789_, _01887_);
  and (_06791_, _06789_, _01887_);
  or (_06792_, _06791_, _06790_);
  and (_06793_, _06792_, _06786_);
  and (_06794_, _06793_, _06780_);
  and (_06795_, _06789_, \oc8051_golden_model_1.ACC [0]);
  nor (_06796_, _06795_, _06784_);
  or (_06797_, _06796_, _06785_);
  and (_06798_, _06797_, _06780_);
  not (_06799_, _06798_);
  and (_06800_, _06778_, _06774_);
  nor (_06801_, _06800_, _06773_);
  and (_06802_, _06801_, _06799_);
  nor (_06803_, _06802_, _06794_);
  not (_06804_, _06803_);
  and (_06805_, _06804_, _06769_);
  nor (_06806_, _06766_, _06761_);
  nor (_06807_, _06806_, _06762_);
  or (_06808_, _06807_, _06805_);
  and (_06809_, _06808_, _06757_);
  or (_06810_, _06809_, _06755_);
  and (_06811_, _06810_, _06752_);
  nor (_06812_, _06810_, _06752_);
  or (_06813_, _06812_, _06811_);
  or (_06814_, _06813_, _06741_);
  and (_06815_, _02030_, _01766_);
  nand (_06816_, _01766_, _01693_);
  not (_06817_, _06816_);
  nor (_06818_, _02590_, _02528_);
  nor (_06819_, _03315_, _02581_);
  and (_06820_, _06819_, _06818_);
  not (_06821_, _06820_);
  nand (_06822_, _06821_, _03796_);
  and (_06823_, _02245_, _02056_);
  nor (_06824_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06825_, _06824_, _06377_);
  and (_06826_, _06825_, _06248_);
  and (_06827_, _06826_, \oc8051_golden_model_1.ACC [6]);
  and (_06828_, _06827_, \oc8051_golden_model_1.ACC [7]);
  nor (_06829_, _06827_, \oc8051_golden_model_1.ACC [7]);
  nor (_06830_, _06829_, _06828_);
  and (_06831_, _06825_, \oc8051_golden_model_1.ACC [4]);
  nor (_06832_, _06831_, \oc8051_golden_model_1.ACC [5]);
  nor (_06833_, _06832_, _06826_);
  nor (_06834_, _06826_, \oc8051_golden_model_1.ACC [6]);
  nor (_06835_, _06834_, _06827_);
  nor (_06836_, _06835_, _06833_);
  not (_06837_, _06836_);
  and (_06838_, _06837_, _06830_);
  nor (_06839_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_06840_, _06839_, _06836_);
  nor (_06841_, _06840_, _06830_);
  nor (_06842_, _06841_, _06838_);
  not (_06843_, _06842_);
  nand (_06844_, _06843_, _06823_);
  and (_06845_, _02245_, _02159_);
  nor (_06846_, _06845_, _02158_);
  not (_06847_, _02160_);
  nor (_06848_, _04682_, _06847_);
  not (_06849_, _02552_);
  or (_06850_, _04637_, _06849_);
  nor (_06851_, _05442_, _01751_);
  nor (_06852_, _06851_, _02560_);
  not (_06853_, _06852_);
  nand (_06854_, _06853_, _03796_);
  and (_06855_, _02245_, _02061_);
  nor (_06856_, _06855_, _04939_);
  and (_06857_, _06855_, _04939_);
  nor (_06858_, _06857_, _06856_);
  and (_06859_, _06852_, _06849_);
  nand (_06860_, _06859_, _06858_);
  and (_06861_, _06860_, _06854_);
  and (_06862_, _06861_, _06847_);
  and (_06863_, _06862_, _06850_);
  or (_06864_, _06863_, _06848_);
  and (_06865_, _06864_, _06846_);
  and (_06866_, _04650_, _03841_);
  nor (_06867_, _06866_, _06735_);
  nor (_06868_, _06867_, _03006_);
  or (_06869_, _06868_, _06823_);
  or (_06870_, _06869_, _06865_);
  and (_06871_, _06870_, _06844_);
  or (_06872_, _06871_, _02057_);
  nor (_06873_, _04483_, _04939_);
  and (_06874_, _04521_, _04483_);
  nor (_06875_, _06874_, _06873_);
  nand (_06876_, _06875_, _02057_);
  and (_06877_, _06876_, _02519_);
  and (_06878_, _06877_, _06872_);
  nor (_06879_, _06738_, _02519_);
  or (_06880_, _06879_, _06821_);
  or (_06881_, _06880_, _06878_);
  and (_06882_, _06881_, _06822_);
  or (_06883_, _06882_, _02582_);
  not (_06884_, _02582_);
  or (_06885_, _04637_, _06884_);
  and (_06886_, _06885_, _02549_);
  and (_06887_, _06886_, _06883_);
  and (_06888_, _02245_, _02051_);
  nor (_06889_, _04682_, _02549_);
  or (_06890_, _06889_, _06888_);
  or (_06891_, _06890_, _06887_);
  nand (_06892_, _06888_, _06377_);
  and (_06893_, _06892_, _06891_);
  or (_06894_, _06893_, _02053_);
  and (_06895_, _04517_, _04483_);
  nor (_06896_, _06895_, _06873_);
  nand (_06897_, _06896_, _02053_);
  and (_06898_, _06897_, _02047_);
  and (_06899_, _06898_, _06894_);
  and (_06900_, _06874_, _04687_);
  nor (_06901_, _06900_, _06873_);
  nor (_06902_, _06901_, _02047_);
  or (_06903_, _06902_, _05474_);
  or (_06904_, _06903_, _06899_);
  nor (_06905_, _06145_, _06143_);
  nor (_06906_, _06905_, _06146_);
  or (_06907_, _06906_, _06181_);
  and (_06908_, _06907_, _06904_);
  or (_06909_, _06908_, _06817_);
  not (_06910_, _06663_);
  and (_06911_, _06684_, _06676_);
  not (_06912_, _06911_);
  and (_06913_, _06699_, _06693_);
  nor (_06914_, _06709_, _01887_);
  nor (_06915_, _06914_, _06705_);
  nor (_06916_, _06915_, _06704_);
  not (_06917_, _06916_);
  and (_06918_, _06917_, _06913_);
  not (_06919_, _06918_);
  and (_06920_, _06698_, _06693_);
  nor (_06921_, _06920_, _06692_);
  and (_06922_, _06921_, _06919_);
  and (_06923_, _06709_, _01887_);
  nor (_06924_, _06914_, _06923_);
  and (_06925_, _06924_, _06706_);
  and (_06926_, _06925_, _06913_);
  nor (_06927_, _06926_, _06922_);
  nor (_06928_, _06927_, _06912_);
  not (_06929_, _06928_);
  and (_06930_, _06682_, _06676_);
  nor (_06931_, _06930_, _06675_);
  and (_06932_, _06931_, _06929_);
  nor (_06933_, _06932_, _06668_);
  or (_06934_, _06933_, _06667_);
  and (_06935_, _06934_, _06910_);
  nor (_06936_, _06934_, _06910_);
  or (_06937_, _06936_, _06935_);
  or (_06938_, _06937_, _06816_);
  and (_06939_, _06938_, _06909_);
  or (_06940_, _06939_, _06815_);
  not (_06941_, _06815_);
  and (_06942_, _05369_, \oc8051_golden_model_1.PSW [7]);
  nor (_06943_, _06942_, _04698_);
  and (_06944_, _06942_, _04698_);
  nor (_06945_, _06944_, _06943_);
  and (_06946_, _06945_, \oc8051_golden_model_1.ACC [7]);
  nor (_06947_, _06945_, \oc8051_golden_model_1.ACC [7]);
  nor (_06948_, _06947_, _06946_);
  and (_06949_, _05368_, \oc8051_golden_model_1.PSW [7]);
  nor (_06950_, _06949_, _05029_);
  nor (_06951_, _06950_, _06942_);
  nor (_06952_, _06951_, _06231_);
  and (_06953_, _06951_, _06231_);
  and (_06954_, _05366_, _05303_);
  and (_06955_, _06954_, \oc8051_golden_model_1.PSW [7]);
  nor (_06956_, _06955_, _05258_);
  nor (_06957_, _06956_, _06949_);
  and (_06958_, _06957_, _06277_);
  nor (_06959_, _06957_, _06277_);
  and (_06960_, _05364_, \oc8051_golden_model_1.PSW [7]);
  and (_06961_, _06960_, _05365_);
  nor (_06962_, _06961_, _05303_);
  nor (_06963_, _06962_, _06955_);
  nor (_06964_, _06963_, _06283_);
  nor (_06965_, _06964_, _06959_);
  nor (_06966_, _06965_, _06958_);
  nor (_06967_, _06959_, _06958_);
  and (_06968_, _06963_, _06283_);
  nor (_06969_, _06968_, _06964_);
  and (_06970_, _06969_, _06967_);
  not (_06971_, _06970_);
  and (_06972_, _05364_, _05211_);
  and (_06973_, _06972_, \oc8051_golden_model_1.PSW [7]);
  nor (_06974_, _06973_, _05166_);
  nor (_06975_, _06974_, _06961_);
  nor (_06976_, _06975_, _06377_);
  and (_06977_, _06975_, _06377_);
  nor (_06978_, _06977_, _06976_);
  nor (_06979_, _06960_, _05211_);
  nor (_06980_, _06979_, _06973_);
  nor (_06981_, _06980_, _06383_);
  and (_06982_, _06980_, _06383_);
  nor (_06983_, _06982_, _06981_);
  and (_06984_, _06983_, _06978_);
  and (_06985_, _05120_, \oc8051_golden_model_1.PSW [7]);
  nor (_06986_, _06985_, _05075_);
  nor (_06987_, _06986_, _06960_);
  and (_06988_, _06987_, _01804_);
  nor (_06989_, _06987_, _01804_);
  nor (_06990_, _05120_, \oc8051_golden_model_1.PSW [7]);
  nor (_06991_, _06990_, _06985_);
  nor (_06992_, _06991_, _01887_);
  nor (_06993_, _06992_, _06989_);
  or (_06994_, _06993_, _06988_);
  and (_06995_, _06994_, _06984_);
  not (_06996_, _06995_);
  and (_06997_, _06982_, _06978_);
  nor (_06998_, _06997_, _06977_);
  and (_06999_, _06998_, _06996_);
  nor (_07000_, _06989_, _06988_);
  and (_07001_, _06991_, _01887_);
  nor (_07002_, _06992_, _07001_);
  and (_07003_, _07002_, _07000_);
  and (_07004_, _07003_, _06984_);
  nor (_07005_, _07004_, _06999_);
  nor (_07006_, _07005_, _06971_);
  nor (_07007_, _07006_, _06966_);
  nor (_07008_, _07007_, _06953_);
  or (_07009_, _07008_, _06952_);
  or (_07010_, _07009_, _06948_);
  nand (_07011_, _07009_, _06948_);
  and (_07012_, _07011_, _07010_);
  or (_07013_, _07012_, _06941_);
  and (_07014_, _07013_, _02191_);
  and (_07015_, _07014_, _06940_);
  nor (_07016_, _06740_, _02186_);
  not (_07017_, _07016_);
  not (_07018_, _03984_);
  nor (_07019_, _03987_, _03983_);
  and (_07020_, _07019_, _03995_);
  and (_07021_, _07020_, _07018_);
  and (_07022_, _07021_, _04007_);
  not (_07023_, _03971_);
  and (_07024_, _03992_, _07023_);
  and (_07025_, _07024_, _03968_);
  and (_07026_, _03830_, \oc8051_golden_model_1.P2INREG [6]);
  and (_07027_, _03820_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_07028_, _07027_, _07026_);
  and (_07029_, _03859_, \oc8051_golden_model_1.P1INREG [6]);
  and (_07030_, _03885_, \oc8051_golden_model_1.P0INREG [6]);
  nor (_07031_, _07030_, _07029_);
  and (_07032_, _07031_, _07028_);
  and (_07033_, _07032_, _03982_);
  and (_07034_, _07033_, _07025_);
  and (_07035_, _07034_, _07022_);
  and (_07036_, _07035_, _03965_);
  not (_07037_, _07036_);
  not (_07038_, _04126_);
  nor (_07039_, _04129_, _04125_);
  and (_07040_, _07039_, _04137_);
  and (_07041_, _07040_, _07038_);
  and (_07042_, _07041_, _04149_);
  not (_07043_, _04111_);
  and (_07044_, _04108_, _07043_);
  and (_07045_, _07044_, _04134_);
  and (_07046_, _03830_, \oc8051_golden_model_1.P2INREG [3]);
  and (_07047_, _03820_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_07048_, _07047_, _07046_);
  and (_07049_, _03859_, \oc8051_golden_model_1.P1INREG [3]);
  and (_07050_, _03885_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_07051_, _07050_, _07049_);
  and (_07052_, _07051_, _07048_);
  and (_07053_, _07052_, _04124_);
  and (_07054_, _07053_, _07045_);
  and (_07055_, _07054_, _07042_);
  and (_07056_, _07055_, _04105_);
  not (_07057_, _07056_);
  and (_07058_, _03830_, \oc8051_golden_model_1.P2INREG [2]);
  and (_07059_, _03820_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_07060_, _07059_, _07058_);
  and (_07061_, _03859_, \oc8051_golden_model_1.P1INREG [2]);
  and (_07062_, _03885_, \oc8051_golden_model_1.P0INREG [2]);
  nor (_07063_, _07062_, _07061_);
  and (_07064_, _07063_, _07060_);
  and (_07065_, _07064_, _04295_);
  and (_07066_, _07065_, _04289_);
  and (_07067_, _07066_, _04273_);
  and (_07068_, _07067_, _04259_);
  not (_07069_, _07068_);
  and (_07070_, _04162_, \oc8051_golden_model_1.P0INREG [1]);
  not (_07071_, _07070_);
  and (_07072_, _03859_, \oc8051_golden_model_1.P1INREG [1]);
  not (_07073_, _07072_);
  and (_07074_, _03830_, \oc8051_golden_model_1.P2INREG [1]);
  and (_07075_, _03820_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_07076_, _07075_, _07074_);
  and (_07077_, _07076_, _07073_);
  and (_07078_, _07077_, _04161_);
  and (_07079_, _07078_, _07071_);
  and (_07080_, _07079_, _04185_);
  and (_07081_, _07080_, _04206_);
  and (_07082_, _07081_, _04154_);
  not (_07083_, _07082_);
  and (_07084_, _03830_, \oc8051_golden_model_1.P2INREG [0]);
  and (_07085_, _03820_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_07086_, _07085_, _07084_);
  and (_07087_, _03859_, \oc8051_golden_model_1.P1INREG [0]);
  and (_07088_, _03885_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_07089_, _07088_, _07087_);
  and (_07090_, _07089_, _07086_);
  and (_07091_, _07090_, _04244_);
  and (_07092_, _07091_, _04241_);
  and (_07093_, _07092_, _04228_);
  and (_07094_, _07093_, _04210_);
  nor (_07095_, _07094_, _06707_);
  and (_07096_, _07095_, _07083_);
  and (_07097_, _07096_, _07069_);
  and (_07098_, _07097_, _07057_);
  not (_07099_, _04076_);
  nor (_07100_, _04080_, _04077_);
  and (_07101_, _07100_, _04088_);
  and (_07102_, _07101_, _07099_);
  and (_07103_, _07102_, _04100_);
  and (_07104_, _04085_, _04064_);
  and (_07105_, _03830_, \oc8051_golden_model_1.P2INREG [5]);
  and (_07106_, _03820_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_07107_, _07106_, _07105_);
  and (_07108_, _03859_, \oc8051_golden_model_1.P1INREG [5]);
  and (_07109_, _03885_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_07110_, _07109_, _07108_);
  and (_07111_, _07110_, _07107_);
  and (_07112_, _07111_, _04075_);
  and (_07113_, _07112_, _07104_);
  and (_07114_, _07113_, _07103_);
  and (_07115_, _07114_, _04058_);
  and (_07116_, _03830_, \oc8051_golden_model_1.P2INREG [4]);
  and (_07117_, _03820_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_07118_, _07117_, _07116_);
  and (_07119_, _03859_, \oc8051_golden_model_1.P1INREG [4]);
  and (_07120_, _03885_, \oc8051_golden_model_1.P0INREG [4]);
  nor (_07121_, _07120_, _07119_);
  and (_07122_, _07121_, _07118_);
  and (_07123_, _07122_, _04380_);
  and (_07124_, _07123_, _04399_);
  and (_07125_, _07124_, _04417_);
  and (_07126_, _07125_, _04373_);
  nor (_07127_, _07126_, _07115_);
  and (_07128_, _07127_, _07098_);
  and (_07129_, _07128_, _07037_);
  nor (_07130_, _07129_, _04682_);
  and (_07131_, _07129_, _04682_);
  nor (_07132_, _07131_, _07130_);
  and (_07133_, _07132_, \oc8051_golden_model_1.ACC [7]);
  nor (_07134_, _07132_, \oc8051_golden_model_1.ACC [7]);
  nor (_07135_, _07134_, _07133_);
  not (_07136_, _07135_);
  nor (_07137_, _07128_, _07037_);
  nor (_07138_, _07137_, _07129_);
  nor (_07139_, _07138_, _06231_);
  and (_07140_, _07138_, _06231_);
  not (_07141_, _07115_);
  not (_07142_, _07126_);
  and (_07143_, _07098_, _07142_);
  nor (_07144_, _07143_, _07141_);
  nor (_07145_, _07144_, _07128_);
  and (_07146_, _07145_, _06277_);
  nor (_07147_, _07145_, _06277_);
  nor (_07148_, _07098_, _07142_);
  nor (_07149_, _07148_, _07143_);
  nor (_07150_, _07149_, _06283_);
  nor (_07151_, _07150_, _07147_);
  nor (_07152_, _07151_, _07146_);
  nor (_07153_, _07147_, _07146_);
  and (_07154_, _07149_, _06283_);
  nor (_07155_, _07154_, _07150_);
  and (_07156_, _07155_, _07153_);
  not (_07157_, _07156_);
  nor (_07158_, _07097_, _07057_);
  nor (_07159_, _07158_, _07098_);
  nor (_07160_, _07159_, _06377_);
  and (_07161_, _07159_, _06377_);
  nor (_07162_, _07161_, _07160_);
  nor (_07164_, _07096_, _07069_);
  nor (_07165_, _07164_, _07097_);
  nor (_07166_, _07165_, _06383_);
  and (_07167_, _07165_, _06383_);
  nor (_07168_, _07167_, _07166_);
  and (_07169_, _07168_, _07162_);
  not (_07170_, _07169_);
  nor (_07171_, _07095_, _07083_);
  nor (_07172_, _07171_, _07096_);
  and (_07173_, _07172_, _01804_);
  nor (_07174_, _07172_, _01804_);
  and (_07175_, _07094_, _06707_);
  nor (_07176_, _07175_, _07095_);
  nor (_07177_, _07176_, _01887_);
  nor (_07178_, _07177_, _07174_);
  nor (_07179_, _07178_, _07173_);
  nor (_07180_, _07179_, _07170_);
  and (_07181_, _07167_, _07162_);
  nor (_07182_, _07181_, _07161_);
  not (_07183_, _07182_);
  nor (_07184_, _07183_, _07180_);
  and (_07185_, _07176_, _01887_);
  nor (_07186_, _07177_, _07185_);
  nor (_07187_, _07082_, \oc8051_golden_model_1.ACC [1]);
  and (_07188_, _07082_, \oc8051_golden_model_1.ACC [1]);
  nor (_07189_, _07188_, _07187_);
  and (_07190_, \oc8051_golden_model_1.PSW [7], _01887_);
  and (_07191_, _06707_, \oc8051_golden_model_1.ACC [0]);
  nor (_07192_, _07094_, _07191_);
  nor (_07193_, _07192_, _07190_);
  and (_07194_, _07193_, _07189_);
  nor (_07195_, _07193_, _07189_);
  or (_07196_, _07195_, _07194_);
  nand (_07197_, _07196_, _07186_);
  nor (_07198_, _07197_, _07170_);
  nor (_07199_, _07198_, _07184_);
  nor (_07200_, _07199_, _07157_);
  nor (_07201_, _07200_, _07152_);
  nor (_07202_, _07201_, _07140_);
  or (_07203_, _07202_, _07139_);
  and (_07204_, _07203_, _07136_);
  nor (_07205_, _07203_, _07136_);
  nor (_07206_, _07205_, _07204_);
  nand (_07207_, _07206_, _06741_);
  and (_07208_, _07207_, _07017_);
  or (_07209_, _07208_, _07015_);
  and (_07210_, _07209_, _06814_);
  or (_07211_, _07210_, _01876_);
  or (_07212_, _01952_, _01778_);
  and (_07213_, _07212_, _02043_);
  and (_07214_, _07213_, _07211_);
  not (_07215_, _04483_);
  nor (_07216_, _04503_, _07215_);
  nor (_07217_, _07216_, _06873_);
  nor (_07218_, _07217_, _02043_);
  or (_07219_, _07218_, _06188_);
  or (_07220_, _07219_, _07214_);
  and (_07221_, _07220_, _06739_);
  or (_07222_, _07221_, _02031_);
  and (_07223_, _04637_, _03841_);
  or (_07224_, _07223_, _06735_);
  or (_07225_, _07224_, _02032_);
  and (_07226_, _07225_, _02037_);
  and (_07227_, _07226_, _07222_);
  nor (_07228_, _04910_, _06736_);
  nor (_07229_, _07228_, _06735_);
  nor (_07230_, _07229_, _02037_);
  or (_07231_, _07230_, _06202_);
  or (_07232_, _07231_, _07227_);
  or (_07233_, _06220_, _06560_);
  and (_07234_, _07233_, _07232_);
  or (_07235_, _07234_, _01775_);
  or (_07236_, _01952_, _01776_);
  and (_07237_, _07236_, _07235_);
  or (_07238_, _07237_, _01994_);
  and (_07239_, _02245_, _01717_);
  not (_07240_, _07239_);
  and (_07241_, _04716_, _03841_);
  nor (_07242_, _07241_, _06735_);
  nand (_07243_, _07242_, _01994_);
  and (_07244_, _07243_, _07240_);
  and (_07245_, _07244_, _07238_);
  and (_07246_, _07239_, _01952_);
  not (_07247_, _01721_);
  nor (_07248_, _02141_, _07247_);
  or (_07249_, _07248_, _07246_);
  or (_07250_, _07249_, _07245_);
  not (_07251_, _07248_);
  or (_07252_, _07251_, _06617_);
  nor (_07253_, _02902_, _02693_);
  and (_07254_, _07253_, _07252_);
  and (_07255_, _07254_, _07250_);
  not (_07256_, _07253_);
  and (_07257_, _07256_, _06617_);
  and (_07258_, _02133_, _01721_);
  and (_07259_, _02691_, _01630_);
  or (_07260_, _07259_, _07258_);
  or (_07261_, _07260_, _07257_);
  or (_07262_, _07261_, _07255_);
  and (_07263_, _02030_, _01721_);
  not (_07264_, _07263_);
  not (_07265_, _06617_);
  nand (_07266_, _07260_, _07265_);
  and (_07267_, _07266_, _07264_);
  and (_07268_, _07267_, _07262_);
  and (_07269_, _04698_, _04939_);
  and (_07270_, _04637_, \oc8051_golden_model_1.ACC [7]);
  nor (_07271_, _07270_, _07269_);
  and (_07272_, _07271_, _07263_);
  or (_07273_, _07272_, _02329_);
  or (_07274_, _07273_, _07268_);
  or (_07275_, _04942_, _02330_);
  and (_07276_, _07275_, _07274_);
  or (_07277_, _07276_, _06734_);
  nor (_07278_, _01952_, \oc8051_golden_model_1.ACC [7]);
  and (_07279_, _01952_, \oc8051_golden_model_1.ACC [7]);
  nor (_07280_, _07279_, _07278_);
  not (_07281_, _06734_);
  or (_07282_, _07281_, _07280_);
  and (_07283_, _07282_, _07277_);
  or (_07284_, _07283_, _02210_);
  and (_07285_, _04933_, _03841_);
  nor (_07286_, _07285_, _06735_);
  nand (_07287_, _07286_, _02210_);
  and (_07288_, _07287_, _03061_);
  and (_07289_, _07288_, _07284_);
  and (_07290_, _06735_, _02331_);
  not (_07291_, _01727_);
  nor (_07292_, _02141_, _07291_);
  or (_07293_, _07292_, _07290_);
  or (_07294_, _07293_, _07289_);
  not (_07295_, _07292_);
  nor (_07296_, _07295_, _06616_);
  nor (_07297_, _03314_, _02138_);
  nor (_07298_, _07297_, _07291_);
  nor (_07299_, _07298_, _07296_);
  and (_07300_, _07299_, _07294_);
  and (_07301_, _07298_, _06616_);
  or (_07302_, _07301_, _02702_);
  or (_07303_, _07302_, _07300_);
  and (_07304_, _02030_, _01727_);
  not (_07305_, _07304_);
  or (_07306_, _06616_, _02703_);
  and (_07307_, _07306_, _07305_);
  and (_07308_, _07307_, _07303_);
  and (_07309_, _07270_, _07304_);
  or (_07310_, _07309_, _02340_);
  or (_07311_, _07310_, _07308_);
  and (_07312_, _02245_, _01727_);
  not (_07313_, _07312_);
  or (_07314_, _04941_, _02341_);
  and (_07315_, _07314_, _07313_);
  and (_07316_, _07315_, _07311_);
  and (_07317_, _07312_, _07279_);
  or (_07318_, _07317_, _07316_);
  and (_07319_, _07318_, _02208_);
  or (_07320_, _07242_, _04940_);
  nor (_07321_, _07320_, _02208_);
  or (_07322_, _07321_, _06732_);
  or (_07323_, _07322_, _07319_);
  and (_07324_, _07323_, _06733_);
  and (_07325_, _03314_, _01735_);
  or (_07326_, _07325_, _07324_);
  not (_07327_, _02719_);
  nand (_07328_, _07325_, _06615_);
  and (_07329_, _07328_, _07327_);
  and (_07330_, _07329_, _07326_);
  and (_07331_, _02030_, _01735_);
  nor (_07332_, _06615_, _07327_);
  or (_07333_, _07332_, _07331_);
  or (_07334_, _07333_, _07330_);
  nand (_07335_, _07269_, _07331_);
  and (_07336_, _07335_, _02337_);
  and (_07337_, _07336_, _07334_);
  and (_07338_, _02245_, _01735_);
  nor (_07339_, _07338_, _02336_);
  not (_07340_, _07339_);
  not (_07341_, _07338_);
  nand (_07342_, _07341_, _04940_);
  and (_07343_, _07342_, _07340_);
  or (_07344_, _07343_, _07337_);
  nand (_07345_, _07338_, _07278_);
  and (_07346_, _07345_, _04953_);
  and (_07347_, _07346_, _07344_);
  not (_07348_, _06730_);
  nor (_07349_, _04932_, _06736_);
  nor (_07350_, _07349_, _06735_);
  nor (_07351_, _07350_, _04953_);
  or (_07352_, _07351_, _07348_);
  or (_07353_, _07352_, _07347_);
  and (_07354_, _07353_, _06731_);
  or (_07355_, _07354_, _06654_);
  not (_07356_, _06654_);
  and (_07357_, _06951_, \oc8051_golden_model_1.ACC [6]);
  nor (_07358_, _06952_, _06953_);
  and (_07359_, _06957_, \oc8051_golden_model_1.ACC [5]);
  and (_07360_, _06963_, \oc8051_golden_model_1.ACC [4]);
  and (_07361_, _06975_, \oc8051_golden_model_1.ACC [3]);
  and (_07362_, _06980_, \oc8051_golden_model_1.ACC [2]);
  and (_07363_, _06987_, \oc8051_golden_model_1.ACC [1]);
  and (_07364_, _06991_, \oc8051_golden_model_1.ACC [0]);
  not (_07365_, _07364_);
  nor (_07366_, _07365_, _07000_);
  nor (_07367_, _07366_, _07363_);
  nor (_07368_, _07367_, _06983_);
  nor (_07369_, _07368_, _07362_);
  nor (_07370_, _07369_, _06978_);
  nor (_07371_, _07370_, _07361_);
  nor (_07372_, _07371_, _06969_);
  nor (_07373_, _07372_, _07360_);
  nor (_07374_, _07373_, _06967_);
  nor (_07375_, _07374_, _07359_);
  nor (_07376_, _07375_, _07358_);
  nor (_07377_, _07376_, _07357_);
  nor (_07378_, _07377_, _06948_);
  and (_07379_, _07377_, _06948_);
  nor (_07380_, _07379_, _07378_);
  or (_07381_, _07380_, _07356_);
  and (_07382_, _07381_, _02346_);
  and (_07383_, _07382_, _07355_);
  and (_07384_, _02245_, _01725_);
  nor (_07385_, _07384_, _02345_);
  not (_07386_, _07385_);
  and (_07387_, _07138_, \oc8051_golden_model_1.ACC [6]);
  nor (_07388_, _07139_, _07140_);
  and (_07389_, _07145_, \oc8051_golden_model_1.ACC [5]);
  and (_07390_, _07149_, \oc8051_golden_model_1.ACC [4]);
  and (_07391_, _07159_, \oc8051_golden_model_1.ACC [3]);
  and (_07392_, _07165_, \oc8051_golden_model_1.ACC [2]);
  and (_07393_, _07172_, \oc8051_golden_model_1.ACC [1]);
  nor (_07394_, _07174_, _07173_);
  and (_07395_, _07176_, \oc8051_golden_model_1.ACC [0]);
  not (_07396_, _07395_);
  nor (_07397_, _07396_, _07394_);
  nor (_07398_, _07397_, _07393_);
  nor (_07399_, _07398_, _07168_);
  nor (_07400_, _07399_, _07392_);
  nor (_07401_, _07400_, _07162_);
  nor (_07402_, _07401_, _07391_);
  nor (_07403_, _07402_, _07155_);
  nor (_07404_, _07403_, _07390_);
  nor (_07405_, _07404_, _07153_);
  nor (_07406_, _07405_, _07389_);
  nor (_07407_, _07406_, _07388_);
  nor (_07408_, _07407_, _07387_);
  nor (_07409_, _07408_, _07135_);
  and (_07410_, _07408_, _07135_);
  nor (_07411_, _07410_, _07409_);
  or (_07412_, _07411_, _07384_);
  and (_07413_, _07412_, _07386_);
  or (_07414_, _07413_, _07383_);
  and (_07415_, _02201_, _01725_);
  not (_07416_, _07415_);
  not (_07417_, _07384_);
  and (_07418_, _06754_, \oc8051_golden_model_1.ACC [6]);
  and (_07419_, _06760_, \oc8051_golden_model_1.ACC [5]);
  and (_07420_, _06765_, \oc8051_golden_model_1.ACC [4]);
  and (_07421_, _06771_, \oc8051_golden_model_1.ACC [3]);
  and (_07422_, _06776_, \oc8051_golden_model_1.ACC [2]);
  and (_07423_, _06783_, \oc8051_golden_model_1.ACC [1]);
  not (_07424_, _06790_);
  nor (_07425_, _07424_, _06786_);
  nor (_07426_, _07425_, _07423_);
  nor (_07427_, _07426_, _06779_);
  nor (_07428_, _07427_, _07422_);
  nor (_07429_, _07428_, _06774_);
  nor (_07430_, _07429_, _07421_);
  nor (_07431_, _07430_, _06768_);
  nor (_07432_, _07431_, _07420_);
  nor (_07433_, _07432_, _06763_);
  nor (_07434_, _07433_, _07419_);
  nor (_07435_, _07434_, _06757_);
  nor (_07436_, _07435_, _07418_);
  nor (_07437_, _07436_, _06751_);
  and (_07438_, _07436_, _06751_);
  nor (_07439_, _07438_, _07437_);
  or (_07440_, _07439_, _07417_);
  and (_07441_, _07440_, _07416_);
  and (_07442_, _07441_, _07414_);
  nand (_07443_, _07415_, \oc8051_golden_model_1.ACC [6]);
  nand (_07444_, _06614_, _07443_);
  or (_07445_, _07444_, _07442_);
  and (_07446_, _07445_, _06653_);
  or (_07447_, _07446_, _06609_);
  not (_07448_, _06609_);
  and (_07449_, _05029_, \oc8051_golden_model_1.ACC [6]);
  nor (_07450_, _05029_, \oc8051_golden_model_1.ACC [6]);
  nor (_07451_, _07449_, _07450_);
  and (_07452_, _05258_, \oc8051_golden_model_1.ACC [5]);
  nor (_07453_, _05258_, \oc8051_golden_model_1.ACC [5]);
  and (_07454_, _05303_, \oc8051_golden_model_1.ACC [4]);
  nor (_07455_, _05303_, \oc8051_golden_model_1.ACC [4]);
  nor (_07456_, _07454_, _07455_);
  nor (_07457_, _05166_, \oc8051_golden_model_1.ACC [3]);
  not (_07458_, _07457_);
  and (_07459_, _05166_, \oc8051_golden_model_1.ACC [3]);
  not (_07460_, _07459_);
  and (_07461_, _05211_, \oc8051_golden_model_1.ACC [2]);
  nor (_07462_, _05211_, \oc8051_golden_model_1.ACC [2]);
  nor (_07463_, _07461_, _07462_);
  not (_07464_, _07463_);
  and (_07465_, _05075_, \oc8051_golden_model_1.ACC [1]);
  nor (_07466_, _05075_, \oc8051_golden_model_1.ACC [1]);
  nor (_07467_, _07465_, _07466_);
  and (_07468_, _05120_, \oc8051_golden_model_1.ACC [0]);
  and (_07469_, _07468_, _07467_);
  nor (_07470_, _07469_, _07465_);
  nor (_07471_, _07470_, _07464_);
  nor (_07472_, _07471_, _07461_);
  nand (_07473_, _07472_, _07460_);
  and (_07474_, _07473_, _07458_);
  and (_07475_, _07474_, _07456_);
  nor (_07476_, _07475_, _07454_);
  nor (_07477_, _07476_, _07453_);
  or (_07478_, _07477_, _07452_);
  and (_07479_, _07478_, _07451_);
  nor (_07480_, _07479_, _07449_);
  nor (_07481_, _07480_, _07271_);
  and (_07482_, _07480_, _07271_);
  or (_07483_, _07482_, _07481_);
  or (_07484_, _07483_, _07448_);
  and (_07485_, _07484_, _02087_);
  and (_07486_, _07485_, _07447_);
  and (_07487_, _02245_, _01737_);
  nor (_07488_, _07487_, _02085_);
  not (_07489_, _07488_);
  and (_07490_, _04682_, _04939_);
  nor (_07491_, _04682_, _04939_);
  nor (_07492_, _07491_, _07490_);
  nor (_07493_, _07036_, _06231_);
  and (_07494_, _07036_, \oc8051_golden_model_1.ACC [6]);
  nor (_07495_, _07036_, \oc8051_golden_model_1.ACC [6]);
  nor (_07496_, _07495_, _07494_);
  nor (_07497_, _07115_, _06277_);
  nor (_07498_, _07115_, \oc8051_golden_model_1.ACC [5]);
  and (_07499_, _07115_, \oc8051_golden_model_1.ACC [5]);
  nor (_07500_, _07499_, _07498_);
  nor (_07501_, _07126_, _06283_);
  and (_07502_, _07126_, \oc8051_golden_model_1.ACC [4]);
  nor (_07503_, _07126_, \oc8051_golden_model_1.ACC [4]);
  nor (_07504_, _07503_, _07502_);
  not (_07505_, _07504_);
  nor (_07506_, _07068_, _06383_);
  and (_07507_, _07068_, \oc8051_golden_model_1.ACC [2]);
  nor (_07508_, _07068_, \oc8051_golden_model_1.ACC [2]);
  nor (_07509_, _07508_, _07507_);
  nor (_07510_, _07082_, _01804_);
  nor (_07511_, _07094_, _01887_);
  not (_07512_, _07511_);
  nor (_07513_, _07512_, _07189_);
  nor (_07514_, _07513_, _07510_);
  nor (_07515_, _07514_, _07509_);
  nor (_07516_, _07515_, _07506_);
  nor (_07517_, _07516_, _07056_);
  or (_07518_, _07517_, \oc8051_golden_model_1.ACC [3]);
  nand (_07519_, _07516_, _07056_);
  and (_07520_, _07519_, _07518_);
  and (_07521_, _07520_, _07505_);
  nor (_07522_, _07521_, _07501_);
  nor (_07523_, _07522_, _07500_);
  nor (_07524_, _07523_, _07497_);
  nor (_07525_, _07524_, _07496_);
  nor (_07526_, _07525_, _07493_);
  nor (_07527_, _07526_, _07492_);
  and (_07528_, _07526_, _07492_);
  or (_07529_, _07528_, _07527_);
  or (_07530_, _07529_, _07487_);
  and (_07531_, _07530_, _07489_);
  or (_07532_, _07531_, _07486_);
  and (_07533_, _02201_, _01737_);
  not (_07534_, _07533_);
  nor (_07535_, _02118_, _06231_);
  and (_07536_, _02118_, _06231_);
  nor (_07537_, _07536_, _07535_);
  nor (_07538_, _02410_, _06277_);
  and (_07539_, _02410_, _06277_);
  or (_07540_, _07539_, _07538_);
  nor (_07541_, _02825_, _06283_);
  and (_07542_, _02825_, _06283_);
  nor (_07543_, _07542_, _07541_);
  nor (_07544_, _01983_, _06377_);
  and (_07545_, _01983_, _06377_);
  nor (_07546_, _02452_, _06383_);
  and (_07547_, _02452_, _06383_);
  nor (_07548_, _07547_, _07546_);
  not (_07549_, _07548_);
  nor (_07550_, _02859_, _01804_);
  and (_07551_, _02859_, _01804_);
  nor (_07552_, _07551_, _07550_);
  nor (_07553_, _02027_, _01887_);
  and (_07554_, _07553_, _07552_);
  nor (_07555_, _07554_, _07550_);
  nor (_07556_, _07555_, _07549_);
  nor (_07557_, _07556_, _07546_);
  nor (_07558_, _07557_, _07545_);
  or (_07559_, _07558_, _07544_);
  and (_07560_, _07559_, _07543_);
  nor (_07561_, _07560_, _07541_);
  nor (_07562_, _07561_, _07540_);
  or (_07563_, _07562_, _07538_);
  and (_07564_, _07563_, _07537_);
  nor (_07565_, _07564_, _07535_);
  nor (_07566_, _07565_, _07280_);
  and (_07567_, _07565_, _07280_);
  nor (_07568_, _07567_, _07566_);
  nand (_07569_, _07568_, _07487_);
  and (_07570_, _07569_, _07534_);
  and (_07571_, _07570_, _07532_);
  and (_07572_, _07533_, \oc8051_golden_model_1.ACC [6]);
  or (_07573_, _07572_, _02366_);
  or (_07574_, _07573_, _07571_);
  and (_07575_, _02245_, _01566_);
  not (_07576_, _07575_);
  nand (_07577_, _06867_, _02366_);
  and (_07578_, _07577_, _07576_);
  and (_07579_, _07578_, _07574_);
  and (_07580_, _02201_, _01566_);
  nor (_07581_, _07580_, _07575_);
  nor (_07582_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_07583_, _07582_, _06323_);
  and (_07584_, _07583_, _06247_);
  and (_07585_, _07584_, _06231_);
  nor (_07586_, _07585_, _04939_);
  and (_07587_, _07585_, _04939_);
  nor (_07588_, _07587_, _07586_);
  not (_07589_, _07588_);
  nor (_07590_, _07589_, _07580_);
  nor (_07591_, _07590_, _07581_);
  or (_07592_, _07591_, _07579_);
  nand (_07593_, _07580_, _06707_);
  and (_07594_, _07593_, _01698_);
  and (_07595_, _07594_, _07592_);
  nor (_07596_, _06896_, _01698_);
  or (_07597_, _07596_, _02081_);
  or (_07598_, _07597_, _07595_);
  and (_07599_, _02245_, _01731_);
  not (_07600_, _07599_);
  and (_07601_, _04426_, _03841_);
  nor (_07602_, _07601_, _06735_);
  nand (_07603_, _07602_, _02081_);
  and (_07604_, _07603_, _07600_);
  and (_07605_, _07604_, _07598_);
  and (_07606_, _02201_, _01731_);
  and (_07607_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_07608_, _07607_, _06324_);
  nor (_07609_, _07608_, _06283_);
  and (_07610_, _07609_, \oc8051_golden_model_1.ACC [5]);
  and (_07611_, _07610_, \oc8051_golden_model_1.ACC [6]);
  nor (_07612_, _07611_, \oc8051_golden_model_1.ACC [7]);
  and (_07613_, _07611_, \oc8051_golden_model_1.ACC [7]);
  nor (_07614_, _07613_, _07612_);
  and (_07615_, _07614_, _07599_);
  or (_07616_, _07615_, _07606_);
  or (_07617_, _07616_, _07605_);
  nand (_07618_, _07606_, _01887_);
  and (_07619_, _07618_, _39632_);
  and (_07620_, _07619_, _07617_);
  or (_07621_, _07620_, _06608_);
  and (_38583_, _07621_, _39026_);
  not (_07622_, \oc8051_golden_model_1.DPL [7]);
  nor (_07623_, _39632_, _07622_);
  nor (_07624_, _04180_, _07622_);
  not (_07625_, _04180_);
  nor (_07626_, _04940_, _07625_);
  or (_07627_, _07626_, _07624_);
  and (_07628_, _07627_, _02334_);
  not (_07629_, _02212_);
  nor (_07630_, _07625_, _03796_);
  or (_07631_, _07630_, _07624_);
  or (_07632_, _07631_, _05444_);
  not (_07633_, _02218_);
  and (_07634_, _04650_, _04180_);
  or (_07635_, _07634_, _07624_);
  or (_07636_, _07635_, _03006_);
  and (_07637_, _03896_, \oc8051_golden_model_1.ACC [7]);
  or (_07638_, _07637_, _07624_);
  and (_07639_, _07638_, _02062_);
  nor (_07640_, _02062_, _07622_);
  or (_07641_, _07640_, _02158_);
  or (_07642_, _07641_, _07639_);
  and (_07643_, _07642_, _02519_);
  and (_07644_, _07643_, _07636_);
  and (_07645_, _07631_, _02155_);
  or (_07646_, _07645_, _02153_);
  or (_07647_, _07646_, _07644_);
  nor (_07648_, _01774_, _01754_);
  not (_07649_, _07648_);
  or (_07650_, _07638_, _02549_);
  and (_07651_, _07650_, _07649_);
  and (_07652_, _07651_, _07647_);
  and (_07653_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_07654_, _07653_, \oc8051_golden_model_1.DPL [2]);
  and (_07655_, _07654_, \oc8051_golden_model_1.DPL [3]);
  and (_07656_, _07655_, \oc8051_golden_model_1.DPL [4]);
  and (_07657_, _07656_, \oc8051_golden_model_1.DPL [5]);
  and (_07658_, _07657_, \oc8051_golden_model_1.DPL [6]);
  nor (_07659_, _07658_, \oc8051_golden_model_1.DPL [7]);
  and (_07660_, _07658_, \oc8051_golden_model_1.DPL [7]);
  nor (_07661_, _07660_, _07659_);
  and (_07662_, _07661_, _07648_);
  or (_07663_, _07662_, _07652_);
  and (_07664_, _07663_, _07633_);
  nor (_07665_, _04458_, _07633_);
  or (_07666_, _07665_, _06188_);
  or (_07667_, _07666_, _07664_);
  and (_07668_, _07667_, _07632_);
  or (_07669_, _07668_, _02031_);
  or (_07670_, _07624_, _02032_);
  and (_07671_, _04637_, _03896_);
  or (_07672_, _07671_, _07670_);
  and (_07673_, _07672_, _02037_);
  and (_07674_, _07673_, _07669_);
  not (_07675_, _03896_);
  nor (_07676_, _04910_, _07675_);
  or (_07677_, _07676_, _07624_);
  and (_07678_, _07677_, _01765_);
  or (_07679_, _07678_, _07674_);
  or (_07680_, _07679_, _07629_);
  and (_07681_, _04933_, _04180_);
  or (_07682_, _07624_, _03059_);
  or (_07683_, _07682_, _07681_);
  and (_07684_, _04716_, _03896_);
  or (_07685_, _07684_, _07624_);
  or (_07686_, _07685_, _01995_);
  and (_07687_, _07686_, _03061_);
  and (_07688_, _07687_, _07683_);
  and (_07689_, _07688_, _07680_);
  and (_07690_, _04942_, _04180_);
  or (_07691_, _07690_, _07624_);
  and (_07692_, _07691_, _02331_);
  or (_07693_, _07692_, _07689_);
  and (_07694_, _07693_, _02208_);
  or (_07695_, _07624_, _03903_);
  and (_07696_, _07685_, _02206_);
  and (_07697_, _07696_, _07695_);
  or (_07698_, _07697_, _07694_);
  and (_07699_, _07698_, _03065_);
  and (_07700_, _07638_, _02342_);
  and (_07701_, _07700_, _07695_);
  or (_07702_, _07701_, _02202_);
  or (_07703_, _07702_, _07699_);
  nor (_07704_, _04932_, _07625_);
  or (_07705_, _07624_, _04953_);
  or (_07706_, _07705_, _07704_);
  and (_07707_, _07706_, _04958_);
  and (_07708_, _07707_, _07703_);
  or (_07709_, _07708_, _07628_);
  and (_07710_, _07709_, _02778_);
  and (_07711_, _07635_, _02366_);
  or (_07712_, _07711_, _02081_);
  or (_07713_, _07712_, _07710_);
  and (_07714_, _04426_, _04180_);
  or (_07715_, _07624_, _02082_);
  or (_07716_, _07715_, _07714_);
  and (_07717_, _07716_, _39632_);
  and (_07718_, _07717_, _07713_);
  or (_07719_, _07718_, _07623_);
  and (_38584_, _07719_, _39026_);
  not (_07720_, \oc8051_golden_model_1.DPH [7]);
  nor (_07721_, _39632_, _07720_);
  nor (_07722_, _04202_, _07720_);
  not (_07723_, _04202_);
  nor (_07724_, _04940_, _07723_);
  or (_07725_, _07724_, _07722_);
  and (_07726_, _07725_, _02334_);
  nor (_07727_, _07723_, _03796_);
  or (_07728_, _07727_, _07722_);
  or (_07729_, _07728_, _05444_);
  and (_07730_, _04650_, _04202_);
  or (_07731_, _07730_, _07722_);
  or (_07732_, _07731_, _03006_);
  and (_07733_, _03889_, \oc8051_golden_model_1.ACC [7]);
  or (_07734_, _07733_, _07722_);
  and (_07735_, _07734_, _02062_);
  nor (_07736_, _02062_, _07720_);
  or (_07737_, _07736_, _02158_);
  or (_07738_, _07737_, _07735_);
  and (_07739_, _07738_, _02519_);
  and (_07740_, _07739_, _07732_);
  and (_07741_, _07728_, _02155_);
  or (_07742_, _07741_, _02153_);
  or (_07743_, _07742_, _07740_);
  or (_07744_, _07734_, _02549_);
  and (_07745_, _07744_, _07649_);
  and (_07746_, _07745_, _07743_);
  not (_07747_, \oc8051_golden_model_1.DPH [2]);
  and (_07748_, _07660_, \oc8051_golden_model_1.DPH [0]);
  nand (_07749_, _07748_, \oc8051_golden_model_1.DPH [1]);
  nor (_07750_, _07749_, _07747_);
  and (_07751_, _07750_, \oc8051_golden_model_1.DPH [3]);
  and (_07752_, _07751_, \oc8051_golden_model_1.DPH [4]);
  and (_07753_, _07752_, \oc8051_golden_model_1.DPH [5]);
  and (_07754_, _07753_, \oc8051_golden_model_1.DPH [6]);
  nor (_07755_, _07754_, _07720_);
  and (_07756_, _07754_, _07720_);
  or (_07757_, _07756_, _07755_);
  and (_07758_, _07757_, _07648_);
  or (_07759_, _07758_, _07746_);
  and (_07760_, _07759_, _07633_);
  and (_07761_, _02218_, _01952_);
  or (_07762_, _07761_, _06188_);
  or (_07763_, _07762_, _07760_);
  and (_07764_, _07763_, _07729_);
  or (_07765_, _07764_, _02031_);
  or (_07766_, _07722_, _02032_);
  and (_07767_, _04637_, _03889_);
  or (_07768_, _07767_, _07766_);
  and (_07769_, _07768_, _02037_);
  and (_07770_, _07769_, _07765_);
  not (_07771_, _03889_);
  nor (_07772_, _04910_, _07771_);
  or (_07773_, _07772_, _07722_);
  and (_07774_, _07773_, _01765_);
  or (_07775_, _07774_, _07770_);
  or (_07776_, _07775_, _07629_);
  and (_07777_, _04933_, _04202_);
  or (_07778_, _07722_, _03059_);
  or (_07779_, _07778_, _07777_);
  and (_07780_, _04716_, _03889_);
  or (_07781_, _07780_, _07722_);
  or (_07782_, _07781_, _01995_);
  and (_07783_, _07782_, _03061_);
  and (_07784_, _07783_, _07779_);
  and (_07785_, _07784_, _07776_);
  and (_07786_, _04942_, _04202_);
  or (_07787_, _07786_, _07722_);
  and (_07788_, _07787_, _02331_);
  or (_07789_, _07788_, _07785_);
  and (_07790_, _07789_, _02208_);
  or (_07791_, _07722_, _03903_);
  and (_07792_, _07781_, _02206_);
  and (_07793_, _07792_, _07791_);
  or (_07794_, _07793_, _07790_);
  and (_07795_, _07794_, _03065_);
  and (_07796_, _07734_, _02342_);
  and (_07797_, _07796_, _07791_);
  or (_07798_, _07797_, _02202_);
  or (_07799_, _07798_, _07795_);
  nor (_07800_, _04932_, _07723_);
  or (_07801_, _07722_, _04953_);
  or (_07802_, _07801_, _07800_);
  and (_07803_, _07802_, _04958_);
  and (_07804_, _07803_, _07799_);
  or (_07805_, _07804_, _07726_);
  and (_07806_, _07805_, _02778_);
  and (_07807_, _07731_, _02366_);
  or (_07808_, _07807_, _02081_);
  or (_07809_, _07808_, _07806_);
  and (_07810_, _04426_, _04202_);
  or (_07811_, _07722_, _02082_);
  or (_07812_, _07811_, _07810_);
  and (_07813_, _07812_, _39632_);
  and (_07814_, _07813_, _07809_);
  or (_07815_, _07814_, _07721_);
  and (_38586_, _07815_, _39026_);
  not (_07816_, \oc8051_golden_model_1.IE [7]);
  nor (_07817_, _03813_, _07816_);
  not (_07818_, _03813_);
  nor (_07819_, _07818_, _03796_);
  nor (_07820_, _07819_, _07817_);
  and (_07821_, _07820_, _06188_);
  nor (_07822_, _04473_, _07816_);
  and (_07823_, _04517_, _04473_);
  nor (_07824_, _07823_, _07822_);
  nor (_07825_, _07824_, _02054_);
  and (_07826_, _03813_, \oc8051_golden_model_1.ACC [7]);
  nor (_07827_, _07826_, _07817_);
  nor (_07828_, _07827_, _02063_);
  nor (_07829_, _02062_, _07816_);
  or (_07830_, _07829_, _07828_);
  and (_07831_, _07830_, _03006_);
  and (_07832_, _04650_, _03813_);
  nor (_07833_, _07832_, _07817_);
  nor (_07834_, _07833_, _03006_);
  or (_07835_, _07834_, _07831_);
  and (_07836_, _07835_, _02058_);
  and (_07837_, _04521_, _04473_);
  nor (_07838_, _07837_, _07822_);
  nor (_07839_, _07838_, _02058_);
  or (_07840_, _07839_, _07836_);
  and (_07841_, _07840_, _02519_);
  nor (_07842_, _07820_, _02519_);
  or (_07843_, _07842_, _07841_);
  and (_07844_, _07843_, _02549_);
  nor (_07845_, _07827_, _02549_);
  or (_07846_, _07845_, _07844_);
  and (_07847_, _07846_, _02054_);
  nor (_07848_, _07847_, _07825_);
  nor (_07849_, _07848_, _02046_);
  nor (_07850_, _07822_, _04687_);
  or (_07851_, _07838_, _02047_);
  nor (_07852_, _07851_, _07850_);
  nor (_07853_, _07852_, _07849_);
  nor (_07854_, _07853_, _02042_);
  not (_07855_, _04473_);
  nor (_07856_, _04503_, _07855_);
  nor (_07857_, _07856_, _07822_);
  nor (_07858_, _07857_, _02043_);
  nor (_07859_, _07858_, _06188_);
  not (_07860_, _07859_);
  nor (_07861_, _07860_, _07854_);
  nor (_07862_, _07861_, _07821_);
  nor (_07863_, _07862_, _02031_);
  and (_07864_, _04637_, _03813_);
  nor (_07865_, _07817_, _02032_);
  not (_07866_, _07865_);
  nor (_07867_, _07866_, _07864_);
  nor (_07868_, _07867_, _01765_);
  not (_07869_, _07868_);
  nor (_07870_, _07869_, _07863_);
  nor (_07871_, _04910_, _07818_);
  nor (_07872_, _07871_, _07817_);
  nor (_07873_, _07872_, _02037_);
  or (_07874_, _07873_, _07629_);
  or (_07875_, _07874_, _07870_);
  and (_07876_, _04933_, _03813_);
  or (_07877_, _07817_, _03059_);
  or (_07878_, _07877_, _07876_);
  and (_07879_, _04716_, _03813_);
  nor (_07880_, _07879_, _07817_);
  and (_07881_, _07880_, _01994_);
  nor (_07882_, _07881_, _02331_);
  and (_07883_, _07882_, _07878_);
  and (_07884_, _07883_, _07875_);
  and (_07885_, _04942_, _03813_);
  nor (_07886_, _07885_, _07817_);
  nor (_07887_, _07886_, _03061_);
  nor (_07888_, _07887_, _07884_);
  nor (_07889_, _07888_, _02206_);
  nor (_07890_, _07817_, _03903_);
  not (_07891_, _07890_);
  nor (_07892_, _07880_, _02208_);
  and (_07893_, _07892_, _07891_);
  nor (_07894_, _07893_, _07889_);
  nor (_07895_, _07894_, _02342_);
  or (_07896_, _07890_, _03065_);
  nor (_07897_, _07896_, _07827_);
  or (_07898_, _07897_, _02202_);
  nor (_07899_, _07898_, _07895_);
  nor (_07900_, _04932_, _07818_);
  or (_07901_, _07817_, _04953_);
  nor (_07902_, _07901_, _07900_);
  or (_07903_, _07902_, _02334_);
  nor (_07904_, _07903_, _07899_);
  nor (_07905_, _04940_, _07818_);
  nor (_07906_, _07905_, _07817_);
  nor (_07907_, _07906_, _04958_);
  or (_07908_, _07907_, _07904_);
  and (_07909_, _07908_, _02778_);
  nor (_07910_, _07833_, _02778_);
  or (_07911_, _07910_, _07909_);
  and (_07912_, _07911_, _01698_);
  nor (_07913_, _07824_, _01698_);
  or (_07914_, _07913_, _07912_);
  and (_07915_, _07914_, _02082_);
  and (_07916_, _04426_, _03813_);
  nor (_07917_, _07916_, _07817_);
  nor (_07918_, _07917_, _02082_);
  or (_07919_, _07918_, _07915_);
  or (_07920_, _07919_, _39633_);
  or (_07921_, _39632_, \oc8051_golden_model_1.IE [7]);
  and (_07922_, _07921_, _39026_);
  and (_38587_, _07922_, _07920_);
  not (_07923_, \oc8051_golden_model_1.IP [7]);
  nor (_07924_, _03844_, _07923_);
  not (_07925_, _03844_);
  nor (_07926_, _07925_, _03796_);
  nor (_07927_, _07926_, _07924_);
  and (_07928_, _07927_, _06188_);
  and (_07929_, _03844_, \oc8051_golden_model_1.ACC [7]);
  nor (_07930_, _07929_, _07924_);
  nor (_07931_, _07930_, _02063_);
  nor (_07932_, _02062_, _07923_);
  or (_07933_, _07932_, _07931_);
  and (_07934_, _07933_, _03006_);
  and (_07935_, _04650_, _03844_);
  nor (_07936_, _07935_, _07924_);
  nor (_07937_, _07936_, _03006_);
  or (_07938_, _07937_, _07934_);
  and (_07939_, _07938_, _02058_);
  nor (_07940_, _04481_, _07923_);
  and (_07941_, _04521_, _04481_);
  nor (_07942_, _07941_, _07940_);
  nor (_07943_, _07942_, _02058_);
  or (_07944_, _07943_, _07939_);
  and (_07945_, _07944_, _02519_);
  nor (_07946_, _07927_, _02519_);
  or (_07947_, _07946_, _07945_);
  and (_07948_, _07947_, _02549_);
  nor (_07949_, _07930_, _02549_);
  or (_07950_, _07949_, _07948_);
  and (_07951_, _07950_, _02054_);
  and (_07952_, _04517_, _04481_);
  nor (_07953_, _07952_, _07940_);
  nor (_07954_, _07953_, _02054_);
  nor (_07955_, _07954_, _07951_);
  nor (_07956_, _07955_, _02046_);
  nor (_07957_, _07940_, _04687_);
  or (_07958_, _07942_, _02047_);
  nor (_07959_, _07958_, _07957_);
  nor (_07960_, _07959_, _07956_);
  nor (_07961_, _07960_, _02042_);
  not (_07962_, _04481_);
  nor (_07963_, _04503_, _07962_);
  nor (_07964_, _07963_, _07940_);
  nor (_07965_, _07964_, _02043_);
  nor (_07966_, _07965_, _06188_);
  not (_07967_, _07966_);
  nor (_07968_, _07967_, _07961_);
  nor (_07969_, _07968_, _07928_);
  nor (_07970_, _07969_, _02031_);
  and (_07971_, _04637_, _03844_);
  nor (_07972_, _07924_, _02032_);
  not (_07973_, _07972_);
  nor (_07974_, _07973_, _07971_);
  nor (_07975_, _07974_, _01765_);
  not (_07976_, _07975_);
  nor (_07977_, _07976_, _07970_);
  nor (_07978_, _04910_, _07925_);
  nor (_07979_, _07978_, _07924_);
  nor (_07980_, _07979_, _02037_);
  or (_07981_, _07980_, _07629_);
  or (_07982_, _07981_, _07977_);
  and (_07983_, _04933_, _03844_);
  or (_07984_, _07924_, _03059_);
  or (_07985_, _07984_, _07983_);
  and (_07986_, _04716_, _03844_);
  nor (_07987_, _07986_, _07924_);
  and (_07988_, _07987_, _01994_);
  nor (_07989_, _07988_, _02331_);
  and (_07990_, _07989_, _07985_);
  and (_07991_, _07990_, _07982_);
  and (_07992_, _04942_, _03844_);
  nor (_07993_, _07992_, _07924_);
  nor (_07994_, _07993_, _03061_);
  nor (_07995_, _07994_, _07991_);
  nor (_07996_, _07995_, _02206_);
  nor (_07997_, _07924_, _03903_);
  not (_07998_, _07997_);
  nor (_07999_, _07987_, _02208_);
  and (_08000_, _07999_, _07998_);
  nor (_08001_, _08000_, _07996_);
  nor (_08002_, _08001_, _02342_);
  or (_08003_, _07997_, _03065_);
  nor (_08004_, _08003_, _07930_);
  or (_08005_, _08004_, _02202_);
  nor (_08006_, _08005_, _08002_);
  nor (_08007_, _04932_, _07925_);
  or (_08008_, _07924_, _04953_);
  nor (_08009_, _08008_, _08007_);
  or (_08010_, _08009_, _02334_);
  nor (_08011_, _08010_, _08006_);
  nor (_08012_, _04940_, _07925_);
  nor (_08013_, _08012_, _07924_);
  nor (_08014_, _08013_, _04958_);
  or (_08015_, _08014_, _08011_);
  and (_08016_, _08015_, _02778_);
  nor (_08017_, _07936_, _02778_);
  or (_08018_, _08017_, _08016_);
  and (_08019_, _08018_, _01698_);
  nor (_08020_, _07953_, _01698_);
  or (_08021_, _08020_, _08019_);
  and (_08022_, _08021_, _02082_);
  and (_08023_, _04426_, _03844_);
  nor (_08024_, _08023_, _07924_);
  nor (_08025_, _08024_, _02082_);
  or (_08026_, _08025_, _08022_);
  or (_08027_, _08026_, _39633_);
  or (_08028_, _39632_, \oc8051_golden_model_1.IP [7]);
  and (_08029_, _08028_, _39026_);
  and (_38588_, _08029_, _08027_);
  nor (_08030_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_08031_, _08030_, _00001_);
  not (_08032_, _03885_);
  and (_08033_, _08032_, \oc8051_golden_model_1.P0 [7]);
  not (_08034_, _04162_);
  nor (_08035_, _08034_, _03796_);
  or (_08036_, _08035_, _08033_);
  or (_08037_, _08036_, _05444_);
  or (_08038_, _08036_, _02519_);
  and (_08039_, _04650_, _04162_);
  or (_08040_, _08039_, _08033_);
  or (_08041_, _08040_, _03006_);
  and (_08042_, _03885_, \oc8051_golden_model_1.ACC [7]);
  or (_08043_, _08042_, _08033_);
  and (_08044_, _08043_, _02062_);
  and (_08045_, _02063_, \oc8051_golden_model_1.P0 [7]);
  or (_08046_, _08045_, _02158_);
  or (_08047_, _08046_, _08044_);
  and (_08048_, _08047_, _02058_);
  and (_08049_, _08048_, _08041_);
  not (_08050_, _03825_);
  and (_08051_, _08050_, \oc8051_golden_model_1.P0 [7]);
  and (_08052_, _04521_, _03825_);
  or (_08053_, _08052_, _08051_);
  and (_08054_, _08053_, _02057_);
  or (_08055_, _08054_, _02155_);
  or (_08056_, _08055_, _08049_);
  and (_08057_, _08056_, _08038_);
  or (_08058_, _08057_, _02153_);
  or (_08059_, _08043_, _02549_);
  and (_08060_, _08059_, _02054_);
  and (_08061_, _08060_, _08058_);
  and (_08062_, _04517_, _03825_);
  or (_08063_, _08062_, _08051_);
  and (_08064_, _08063_, _02053_);
  or (_08065_, _08064_, _08061_);
  and (_08066_, _08065_, _02047_);
  and (_08067_, _04688_, _03825_);
  or (_08068_, _08067_, _08051_);
  and (_08069_, _08068_, _02046_);
  or (_08070_, _08069_, _08066_);
  and (_08071_, _08070_, _02043_);
  or (_08072_, _04517_, _04502_);
  and (_08073_, _08072_, _03825_);
  or (_08074_, _08073_, _08051_);
  and (_08075_, _08074_, _02042_);
  or (_08076_, _08075_, _06188_);
  or (_08077_, _08076_, _08071_);
  and (_08078_, _08077_, _08037_);
  or (_08079_, _08078_, _02031_);
  or (_08080_, _08033_, _02032_);
  and (_08081_, _04637_, _03885_);
  or (_08082_, _08081_, _08080_);
  and (_08083_, _08082_, _02037_);
  and (_08084_, _08083_, _08079_);
  and (_08085_, _04882_, \oc8051_golden_model_1.P1 [7]);
  and (_08086_, _04875_, \oc8051_golden_model_1.P0 [7]);
  and (_08087_, _04885_, \oc8051_golden_model_1.P2 [7]);
  and (_08088_, _04821_, _04817_);
  and (_08089_, _08088_, \oc8051_golden_model_1.P3 [7]);
  or (_08090_, _08089_, _08087_);
  or (_08091_, _08090_, _08086_);
  or (_08092_, _08091_, _08085_);
  nor (_08093_, _08092_, _04873_);
  and (_08094_, _08093_, _04905_);
  and (_08095_, _08094_, _04871_);
  nand (_08096_, _08095_, _04856_);
  or (_08097_, _08096_, _04717_);
  and (_08098_, _08097_, _04162_);
  or (_08099_, _08098_, _08033_);
  and (_08100_, _08099_, _01765_);
  or (_08101_, _08100_, _07629_);
  or (_08102_, _08101_, _08084_);
  and (_08103_, _04933_, _04162_);
  or (_08104_, _08033_, _03059_);
  or (_08105_, _08104_, _08103_);
  and (_08106_, _04716_, _03885_);
  or (_08107_, _08106_, _08033_);
  or (_08108_, _08107_, _01995_);
  and (_08109_, _08108_, _03061_);
  and (_08110_, _08109_, _08105_);
  and (_08111_, _08110_, _08102_);
  and (_08112_, _04942_, _04162_);
  or (_08113_, _08112_, _08033_);
  and (_08114_, _08113_, _02331_);
  or (_08115_, _08114_, _08111_);
  and (_08116_, _08115_, _02208_);
  or (_08117_, _08033_, _03903_);
  and (_08118_, _08107_, _02206_);
  and (_08119_, _08118_, _08117_);
  or (_08120_, _08119_, _08116_);
  and (_08121_, _08120_, _03065_);
  and (_08122_, _08043_, _02342_);
  and (_08123_, _08122_, _08117_);
  or (_08124_, _08123_, _02202_);
  or (_08125_, _08124_, _08121_);
  nor (_08126_, _04932_, _08034_);
  or (_08127_, _08033_, _04953_);
  or (_08128_, _08127_, _08126_);
  and (_08129_, _08128_, _04958_);
  and (_08130_, _08129_, _08125_);
  nor (_08131_, _04940_, _08034_);
  or (_08132_, _08131_, _08033_);
  and (_08133_, _08132_, _02334_);
  or (_08134_, _08133_, _02366_);
  or (_08135_, _08134_, _08130_);
  or (_08136_, _08040_, _02778_);
  and (_08137_, _08136_, _01698_);
  and (_08138_, _08137_, _08135_);
  and (_08139_, _08063_, _01697_);
  or (_08140_, _08139_, _02081_);
  or (_08141_, _08140_, _08138_);
  and (_08142_, _04426_, _04162_);
  or (_08143_, _08033_, _02082_);
  or (_08144_, _08143_, _08142_);
  and (_08145_, _08144_, _39632_);
  and (_08146_, _08145_, _08141_);
  or (_38589_, _08146_, _08031_);
  not (_08147_, \oc8051_golden_model_1.P1 [7]);
  nor (_08148_, _03859_, _08147_);
  not (_08149_, _03859_);
  nor (_08150_, _08149_, _03796_);
  or (_08151_, _08150_, _08148_);
  or (_08152_, _08151_, _05444_);
  or (_08153_, _08151_, _02519_);
  and (_08154_, _04650_, _03859_);
  or (_08155_, _08154_, _08148_);
  or (_08156_, _08155_, _03006_);
  and (_08157_, _03859_, \oc8051_golden_model_1.ACC [7]);
  or (_08158_, _08157_, _08148_);
  and (_08159_, _08158_, _02062_);
  nor (_08160_, _02062_, _08147_);
  or (_08161_, _08160_, _02158_);
  or (_08162_, _08161_, _08159_);
  and (_08163_, _08162_, _02058_);
  and (_08164_, _08163_, _08156_);
  nor (_08165_, _04489_, _08147_);
  and (_08166_, _04521_, _04489_);
  or (_08167_, _08166_, _08165_);
  and (_08168_, _08167_, _02057_);
  or (_08169_, _08168_, _02155_);
  or (_08170_, _08169_, _08164_);
  and (_08171_, _08170_, _08153_);
  or (_08172_, _08171_, _02153_);
  or (_08173_, _08158_, _02549_);
  and (_08174_, _08173_, _02054_);
  and (_08175_, _08174_, _08172_);
  and (_08176_, _04517_, _04489_);
  or (_08177_, _08176_, _08165_);
  and (_08178_, _08177_, _02053_);
  or (_08179_, _08178_, _08175_);
  and (_08180_, _08179_, _02047_);
  or (_08181_, _08165_, _04687_);
  and (_08182_, _08181_, _02046_);
  and (_08183_, _08182_, _08167_);
  or (_08184_, _08183_, _08180_);
  and (_08185_, _08184_, _02043_);
  and (_08186_, _08072_, _04489_);
  or (_08187_, _08186_, _08165_);
  and (_08188_, _08187_, _02042_);
  or (_08189_, _08188_, _06188_);
  or (_08190_, _08189_, _08185_);
  and (_08191_, _08190_, _08152_);
  or (_08192_, _08191_, _02031_);
  and (_08193_, _04637_, _03859_);
  or (_08194_, _08148_, _02032_);
  or (_08195_, _08194_, _08193_);
  and (_08196_, _08195_, _02037_);
  and (_08197_, _08196_, _08192_);
  and (_08198_, _08097_, _03859_);
  or (_08199_, _08198_, _08148_);
  and (_08200_, _08199_, _01765_);
  or (_08201_, _08200_, _07629_);
  or (_08202_, _08201_, _08197_);
  and (_08203_, _04933_, _03859_);
  or (_08204_, _08148_, _03059_);
  or (_08205_, _08204_, _08203_);
  and (_08206_, _04716_, _03859_);
  or (_08207_, _08206_, _08148_);
  or (_08208_, _08207_, _01995_);
  and (_08209_, _08208_, _03061_);
  and (_08211_, _08209_, _08205_);
  and (_08212_, _08211_, _08202_);
  and (_08213_, _04942_, _03859_);
  or (_08214_, _08213_, _08148_);
  and (_08215_, _08214_, _02331_);
  or (_08216_, _08215_, _08212_);
  and (_08217_, _08216_, _02208_);
  or (_08218_, _08148_, _03903_);
  and (_08219_, _08207_, _02206_);
  and (_08220_, _08219_, _08218_);
  or (_08221_, _08220_, _08217_);
  and (_08222_, _08221_, _03065_);
  and (_08223_, _08158_, _02342_);
  and (_08224_, _08223_, _08218_);
  or (_08225_, _08224_, _02202_);
  or (_08226_, _08225_, _08222_);
  nor (_08227_, _04932_, _08149_);
  or (_08228_, _08148_, _04953_);
  or (_08229_, _08228_, _08227_);
  and (_08230_, _08229_, _04958_);
  and (_08231_, _08230_, _08226_);
  nor (_08232_, _04940_, _08149_);
  or (_08233_, _08232_, _08148_);
  and (_08234_, _08233_, _02334_);
  or (_08235_, _08234_, _02366_);
  or (_08236_, _08235_, _08231_);
  or (_08237_, _08155_, _02778_);
  and (_08238_, _08237_, _01698_);
  and (_08239_, _08238_, _08236_);
  and (_08240_, _08177_, _01697_);
  or (_08241_, _08240_, _02081_);
  or (_08242_, _08241_, _08239_);
  and (_08243_, _04426_, _03859_);
  or (_08244_, _08148_, _02082_);
  or (_08245_, _08244_, _08243_);
  and (_08246_, _08245_, _39632_);
  and (_08247_, _08246_, _08242_);
  nor (_08248_, _39632_, _08147_);
  or (_08249_, _08248_, rst);
  or (_38590_, _08249_, _08247_);
  not (_08250_, _03830_);
  and (_08251_, _08250_, \oc8051_golden_model_1.P2 [7]);
  nor (_08252_, _08250_, _03796_);
  or (_08253_, _08252_, _08251_);
  or (_08254_, _08253_, _05444_);
  not (_08255_, \oc8051_golden_model_1.P2 [7]);
  nor (_08256_, _04492_, _08255_);
  and (_08257_, _04517_, _04492_);
  or (_08258_, _08257_, _08256_);
  and (_08259_, _08258_, _02053_);
  or (_08260_, _08253_, _02519_);
  and (_08261_, _04650_, _03830_);
  or (_08262_, _08261_, _08251_);
  or (_08263_, _08262_, _03006_);
  and (_08264_, _03830_, \oc8051_golden_model_1.ACC [7]);
  or (_08265_, _08264_, _08251_);
  and (_08266_, _08265_, _02062_);
  nor (_08267_, _02062_, _08255_);
  or (_08268_, _08267_, _02158_);
  or (_08269_, _08268_, _08266_);
  and (_08270_, _08269_, _02058_);
  and (_08271_, _08270_, _08263_);
  and (_08272_, _04521_, _04492_);
  or (_08273_, _08272_, _08256_);
  and (_08274_, _08273_, _02057_);
  or (_08275_, _08274_, _02155_);
  or (_08276_, _08275_, _08271_);
  and (_08277_, _08276_, _08260_);
  or (_08278_, _08277_, _02153_);
  or (_08279_, _08265_, _02549_);
  and (_08280_, _08279_, _02054_);
  and (_08281_, _08280_, _08278_);
  or (_08282_, _08281_, _08259_);
  and (_08283_, _08282_, _02047_);
  or (_08284_, _08256_, _04687_);
  and (_08285_, _08284_, _02046_);
  and (_08286_, _08285_, _08273_);
  or (_08287_, _08286_, _08283_);
  and (_08288_, _08287_, _02043_);
  and (_08289_, _08072_, _04492_);
  or (_08290_, _08289_, _08256_);
  and (_08291_, _08290_, _02042_);
  or (_08292_, _08291_, _06188_);
  or (_08293_, _08292_, _08288_);
  and (_08294_, _08293_, _08254_);
  or (_08295_, _08294_, _02031_);
  and (_08296_, _04637_, _03830_);
  or (_08297_, _08251_, _02032_);
  or (_08298_, _08297_, _08296_);
  and (_08299_, _08298_, _02037_);
  and (_08300_, _08299_, _08295_);
  and (_08301_, _08097_, _03830_);
  or (_08302_, _08301_, _08251_);
  and (_08303_, _08302_, _01765_);
  or (_08304_, _08303_, _07629_);
  or (_08305_, _08304_, _08300_);
  and (_08306_, _04933_, _03830_);
  or (_08308_, _08251_, _03059_);
  or (_08309_, _08308_, _08306_);
  and (_08311_, _04716_, _03830_);
  or (_08312_, _08311_, _08251_);
  or (_08314_, _08312_, _01995_);
  and (_08315_, _08314_, _03061_);
  and (_08317_, _08315_, _08309_);
  and (_08318_, _08317_, _08305_);
  and (_08319_, _04942_, _03830_);
  or (_08320_, _08319_, _08251_);
  and (_08321_, _08320_, _02331_);
  or (_08322_, _08321_, _08318_);
  and (_08323_, _08322_, _02208_);
  or (_08324_, _08251_, _03903_);
  and (_08325_, _08312_, _02206_);
  and (_08326_, _08325_, _08324_);
  or (_08327_, _08326_, _08323_);
  and (_08328_, _08327_, _03065_);
  and (_08329_, _08265_, _02342_);
  and (_08330_, _08329_, _08324_);
  or (_08331_, _08330_, _02202_);
  or (_08332_, _08331_, _08328_);
  nor (_08333_, _04932_, _08250_);
  or (_08334_, _08251_, _04953_);
  or (_08335_, _08334_, _08333_);
  and (_08336_, _08335_, _04958_);
  and (_08337_, _08336_, _08332_);
  nor (_08338_, _04940_, _08250_);
  or (_08339_, _08338_, _08251_);
  and (_08340_, _08339_, _02334_);
  or (_08341_, _08340_, _02366_);
  or (_08342_, _08341_, _08337_);
  or (_08343_, _08262_, _02778_);
  and (_08344_, _08343_, _01698_);
  and (_08345_, _08344_, _08342_);
  and (_08346_, _08258_, _01697_);
  or (_08347_, _08346_, _02081_);
  or (_08348_, _08347_, _08345_);
  and (_08349_, _04426_, _03830_);
  or (_08350_, _08251_, _02082_);
  or (_08351_, _08350_, _08349_);
  and (_08352_, _08351_, _39632_);
  and (_08353_, _08352_, _08348_);
  nor (_08354_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_08355_, _08354_, _00001_);
  or (_38592_, _08355_, _08353_);
  not (_08356_, \oc8051_golden_model_1.P3 [7]);
  nor (_08357_, _03820_, _08356_);
  not (_08358_, _03820_);
  nor (_08359_, _08358_, _03796_);
  or (_08360_, _08359_, _08357_);
  or (_08361_, _08360_, _05444_);
  nor (_08362_, _04467_, _08356_);
  and (_08363_, _04517_, _04467_);
  or (_08364_, _08363_, _08362_);
  and (_08365_, _08364_, _02053_);
  or (_08366_, _08360_, _02519_);
  and (_08367_, _04650_, _03820_);
  or (_08368_, _08367_, _08357_);
  or (_08369_, _08368_, _03006_);
  and (_08370_, _03820_, \oc8051_golden_model_1.ACC [7]);
  or (_08371_, _08370_, _08357_);
  and (_08372_, _08371_, _02062_);
  nor (_08373_, _02062_, _08356_);
  or (_08374_, _08373_, _02158_);
  or (_08375_, _08374_, _08372_);
  and (_08376_, _08375_, _02058_);
  and (_08377_, _08376_, _08369_);
  and (_08378_, _04521_, _04467_);
  or (_08379_, _08378_, _08362_);
  and (_08380_, _08379_, _02057_);
  or (_08381_, _08380_, _02155_);
  or (_08382_, _08381_, _08377_);
  and (_08383_, _08382_, _08366_);
  or (_08384_, _08383_, _02153_);
  or (_08385_, _08371_, _02549_);
  and (_08386_, _08385_, _02054_);
  and (_08387_, _08386_, _08384_);
  or (_08388_, _08387_, _08365_);
  and (_08389_, _08388_, _02047_);
  and (_08390_, _04688_, _04467_);
  or (_08391_, _08390_, _08362_);
  and (_08392_, _08391_, _02046_);
  or (_08393_, _08392_, _08389_);
  and (_08394_, _08393_, _02043_);
  and (_08395_, _08072_, _04467_);
  or (_08396_, _08395_, _08362_);
  and (_08397_, _08396_, _02042_);
  or (_08398_, _08397_, _06188_);
  or (_08399_, _08398_, _08394_);
  and (_08400_, _08399_, _08361_);
  or (_08401_, _08400_, _02031_);
  and (_08402_, _04637_, _03820_);
  or (_08403_, _08357_, _02032_);
  or (_08404_, _08403_, _08402_);
  and (_08405_, _08404_, _02037_);
  and (_08406_, _08405_, _08401_);
  and (_08407_, _08097_, _03820_);
  or (_08408_, _08407_, _08357_);
  and (_08409_, _08408_, _01765_);
  or (_08410_, _08409_, _07629_);
  or (_08411_, _08410_, _08406_);
  and (_08412_, _04933_, _03820_);
  or (_08413_, _08357_, _03059_);
  or (_08414_, _08413_, _08412_);
  and (_08415_, _04716_, _03820_);
  or (_08416_, _08415_, _08357_);
  or (_08417_, _08416_, _01995_);
  and (_08418_, _08417_, _03061_);
  and (_08419_, _08418_, _08414_);
  and (_08420_, _08419_, _08411_);
  and (_08421_, _04942_, _03820_);
  or (_08422_, _08421_, _08357_);
  and (_08423_, _08422_, _02331_);
  or (_08424_, _08423_, _08420_);
  and (_08425_, _08424_, _02208_);
  or (_08426_, _08357_, _03903_);
  and (_08427_, _08416_, _02206_);
  and (_08428_, _08427_, _08426_);
  or (_08429_, _08428_, _08425_);
  and (_08430_, _08429_, _03065_);
  and (_08431_, _08371_, _02342_);
  and (_08432_, _08431_, _08426_);
  or (_08433_, _08432_, _02202_);
  or (_08434_, _08433_, _08430_);
  nor (_08435_, _04932_, _08358_);
  or (_08436_, _08357_, _04953_);
  or (_08437_, _08436_, _08435_);
  and (_08438_, _08437_, _04958_);
  and (_08439_, _08438_, _08434_);
  nor (_08440_, _04940_, _08358_);
  or (_08441_, _08440_, _08357_);
  and (_08442_, _08441_, _02334_);
  or (_08443_, _08442_, _02366_);
  or (_08444_, _08443_, _08439_);
  or (_08445_, _08368_, _02778_);
  and (_08446_, _08445_, _01698_);
  and (_08447_, _08446_, _08444_);
  and (_08448_, _08364_, _01697_);
  or (_08449_, _08448_, _02081_);
  or (_08450_, _08449_, _08447_);
  and (_08451_, _04426_, _03820_);
  or (_08452_, _08357_, _02082_);
  or (_08453_, _08452_, _08451_);
  and (_08454_, _08453_, _39632_);
  and (_08455_, _08454_, _08450_);
  nor (_08456_, _39632_, _08356_);
  or (_08457_, _08456_, rst);
  or (_38593_, _08457_, _08455_);
  not (_08458_, _07487_);
  not (_08459_, _06616_);
  nor (_08460_, _06649_, _06615_);
  nor (_08461_, _08460_, _06614_);
  and (_08462_, _08461_, _08459_);
  nor (_08463_, _06945_, _04939_);
  nor (_08464_, _08463_, _07378_);
  and (_08465_, _06942_, _04637_);
  nor (_08466_, _08465_, _07356_);
  and (_08468_, _08466_, _08464_);
  and (_08470_, _06656_, _05350_);
  not (_08472_, _08470_);
  nor (_08474_, _06660_, _04939_);
  nor (_08476_, _08474_, _06724_);
  and (_08478_, _08476_, _08472_);
  nor (_08480_, _08478_, _06727_);
  nor (_08482_, _08480_, _06730_);
  nor (_08484_, _03838_, _06707_);
  not (_08485_, _08484_);
  nand (_08486_, _04942_, _03838_);
  and (_08487_, _08486_, _08485_);
  or (_08488_, _08487_, _03061_);
  not (_08489_, _03838_);
  or (_08490_, _04910_, _08489_);
  and (_08491_, _08490_, _08485_);
  or (_08492_, _08491_, _02037_);
  or (_08493_, _08489_, _03796_);
  and (_08494_, _08493_, _08485_);
  and (_08495_, _08494_, _06188_);
  and (_08496_, _06952_, _06948_);
  nor (_08497_, _08496_, _06946_);
  not (_08498_, _08497_);
  and (_08499_, _07358_, _06948_);
  not (_08500_, _08499_);
  nor (_08501_, _08500_, _07007_);
  nor (_08502_, _08501_, _08498_);
  or (_08503_, _08465_, _06941_);
  nor (_08504_, _08503_, _08502_);
  not (_08505_, _02182_);
  not (_08506_, _04179_);
  and (_08507_, _04476_, \oc8051_golden_model_1.PSW [2]);
  and (_08508_, _04478_, \oc8051_golden_model_1.B [2]);
  nor (_08509_, _08508_, _08507_);
  and (_08510_, _04481_, \oc8051_golden_model_1.IP [2]);
  and (_08511_, _04483_, \oc8051_golden_model_1.ACC [2]);
  nor (_08512_, _08511_, _08510_);
  and (_08513_, _08512_, _08509_);
  and (_08514_, _04489_, \oc8051_golden_model_1.P1INREG [2]);
  not (_08515_, _08514_);
  and (_08516_, _03825_, \oc8051_golden_model_1.P0INREG [2]);
  and (_08517_, _04492_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_08518_, _08517_, _08516_);
  and (_08519_, _08518_, _08515_);
  and (_08520_, _04471_, \oc8051_golden_model_1.SCON [2]);
  and (_08521_, _04473_, \oc8051_golden_model_1.IE [2]);
  nor (_08522_, _08521_, _08520_);
  and (_08523_, _04487_, \oc8051_golden_model_1.TCON [2]);
  and (_08524_, _04467_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_08525_, _08524_, _08523_);
  and (_08526_, _08525_, _08522_);
  and (_08527_, _08526_, _08519_);
  and (_08528_, _08527_, _08513_);
  and (_08529_, _08528_, _04259_);
  nor (_08530_, _08529_, _08506_);
  not (_08531_, _03803_);
  and (_08532_, _04471_, \oc8051_golden_model_1.SCON [1]);
  and (_08533_, _04473_, \oc8051_golden_model_1.IE [1]);
  nor (_08534_, _08533_, _08532_);
  and (_08535_, _04487_, \oc8051_golden_model_1.TCON [1]);
  and (_08536_, _04467_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_08537_, _08536_, _08535_);
  and (_08538_, _08537_, _08534_);
  and (_08539_, _04476_, \oc8051_golden_model_1.PSW [1]);
  and (_08540_, _04483_, \oc8051_golden_model_1.ACC [1]);
  nor (_08541_, _08540_, _08539_);
  and (_08542_, _04481_, \oc8051_golden_model_1.IP [1]);
  and (_08543_, _04478_, \oc8051_golden_model_1.B [1]);
  nor (_08544_, _08543_, _08542_);
  and (_08545_, _08544_, _08541_);
  and (_08546_, _04489_, \oc8051_golden_model_1.P1INREG [1]);
  and (_08547_, _04492_, \oc8051_golden_model_1.P2INREG [1]);
  and (_08548_, _03825_, \oc8051_golden_model_1.P0INREG [1]);
  or (_08549_, _08548_, _08547_);
  nor (_08550_, _08549_, _08546_);
  and (_08551_, _08550_, _08545_);
  and (_08552_, _08551_, _08538_);
  and (_08553_, _08552_, _04154_);
  nor (_08554_, _08553_, _08531_);
  nor (_08555_, _08554_, _08530_);
  and (_08556_, _03807_, _02453_);
  not (_08557_, _08556_);
  and (_08558_, _04487_, \oc8051_golden_model_1.TCON [4]);
  and (_08559_, _04483_, \oc8051_golden_model_1.ACC [4]);
  nor (_08560_, _08559_, _08558_);
  and (_08561_, _04481_, \oc8051_golden_model_1.IP [4]);
  not (_08562_, _08561_);
  and (_08563_, _04476_, \oc8051_golden_model_1.PSW [4]);
  and (_08564_, _04478_, \oc8051_golden_model_1.B [4]);
  nor (_08565_, _08564_, _08563_);
  and (_08566_, _08565_, _08562_);
  and (_08567_, _08566_, _08560_);
  and (_08568_, _04471_, \oc8051_golden_model_1.SCON [4]);
  and (_08569_, _04473_, \oc8051_golden_model_1.IE [4]);
  nor (_08570_, _08569_, _08568_);
  and (_08571_, _04489_, \oc8051_golden_model_1.P1INREG [4]);
  and (_08572_, _04467_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_08573_, _08572_, _08571_);
  and (_08574_, _03825_, \oc8051_golden_model_1.P0INREG [4]);
  and (_08575_, _04492_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_08576_, _08575_, _08574_);
  and (_08577_, _08576_, _08573_);
  and (_08578_, _08577_, _08570_);
  and (_08579_, _08578_, _08567_);
  and (_08580_, _08579_, _04373_);
  nor (_08581_, _08580_, _08557_);
  nor (_08582_, _04500_, _04520_);
  nor (_08583_, _08582_, _08581_);
  and (_08584_, _08583_, _08555_);
  not (_08585_, _03808_);
  and (_08586_, _04487_, \oc8051_golden_model_1.TCON [0]);
  and (_08587_, _04478_, \oc8051_golden_model_1.B [0]);
  nor (_08588_, _08587_, _08586_);
  and (_08589_, _04476_, \oc8051_golden_model_1.PSW [0]);
  not (_08590_, _08589_);
  and (_08591_, _04481_, \oc8051_golden_model_1.IP [0]);
  and (_08592_, _04483_, \oc8051_golden_model_1.ACC [0]);
  nor (_08593_, _08592_, _08591_);
  and (_08594_, _08593_, _08590_);
  and (_08595_, _08594_, _08588_);
  and (_08596_, _04471_, \oc8051_golden_model_1.SCON [0]);
  and (_08597_, _04473_, \oc8051_golden_model_1.IE [0]);
  nor (_08598_, _08597_, _08596_);
  and (_08599_, _03825_, \oc8051_golden_model_1.P0INREG [0]);
  and (_08600_, _04492_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_08601_, _08600_, _08599_);
  and (_08602_, _04489_, \oc8051_golden_model_1.P1INREG [0]);
  and (_08603_, _04467_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_08604_, _08603_, _08602_);
  and (_08605_, _08604_, _08601_);
  and (_08606_, _08605_, _08598_);
  and (_08607_, _08606_, _08595_);
  and (_08608_, _08607_, _04210_);
  nor (_08609_, _08608_, _08585_);
  and (_08610_, _03874_, _02453_);
  not (_08611_, _08610_);
  and (_08612_, _04487_, \oc8051_golden_model_1.TCON [6]);
  and (_08613_, _04483_, \oc8051_golden_model_1.ACC [6]);
  nor (_08614_, _08613_, _08612_);
  and (_08615_, _04476_, \oc8051_golden_model_1.PSW [6]);
  not (_08616_, _08615_);
  and (_08617_, _04481_, \oc8051_golden_model_1.IP [6]);
  and (_08618_, _04478_, \oc8051_golden_model_1.B [6]);
  nor (_08619_, _08618_, _08617_);
  and (_08620_, _08619_, _08616_);
  and (_08621_, _08620_, _08614_);
  and (_08622_, _04471_, \oc8051_golden_model_1.SCON [6]);
  and (_08623_, _04473_, \oc8051_golden_model_1.IE [6]);
  nor (_08624_, _08623_, _08622_);
  and (_08625_, _03825_, \oc8051_golden_model_1.P0INREG [6]);
  and (_08626_, _04492_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_08627_, _08626_, _08625_);
  and (_08628_, _04489_, \oc8051_golden_model_1.P1INREG [6]);
  and (_08629_, _04467_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_08630_, _08629_, _08628_);
  and (_08631_, _08630_, _08627_);
  and (_08632_, _08631_, _08624_);
  and (_08633_, _08632_, _08621_);
  and (_08634_, _08633_, _03965_);
  nor (_08635_, _08634_, _08611_);
  nor (_08636_, _08635_, _08609_);
  not (_08637_, _04201_);
  and (_08638_, _04487_, \oc8051_golden_model_1.TCON [3]);
  and (_08639_, _04483_, \oc8051_golden_model_1.ACC [3]);
  nor (_08640_, _08639_, _08638_);
  and (_08641_, _04481_, \oc8051_golden_model_1.IP [3]);
  not (_08642_, _08641_);
  and (_08643_, _04476_, \oc8051_golden_model_1.PSW [3]);
  and (_08644_, _04478_, \oc8051_golden_model_1.B [3]);
  nor (_08645_, _08644_, _08643_);
  and (_08646_, _08645_, _08642_);
  and (_08647_, _08646_, _08640_);
  and (_08648_, _04471_, \oc8051_golden_model_1.SCON [3]);
  and (_08649_, _04473_, \oc8051_golden_model_1.IE [3]);
  nor (_08650_, _08649_, _08648_);
  and (_08651_, _03825_, \oc8051_golden_model_1.P0INREG [3]);
  and (_08652_, _04492_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_08653_, _08652_, _08651_);
  and (_08654_, _04489_, \oc8051_golden_model_1.P1INREG [3]);
  and (_08655_, _04467_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08656_, _08655_, _08654_);
  and (_08657_, _08656_, _08653_);
  and (_08658_, _08657_, _08650_);
  and (_08659_, _08658_, _08647_);
  and (_08660_, _08659_, _04105_);
  nor (_08661_, _08660_, _08637_);
  and (_08662_, _03802_, _02453_);
  not (_08663_, _08662_);
  and (_08664_, _04487_, \oc8051_golden_model_1.TCON [5]);
  and (_08665_, _04478_, \oc8051_golden_model_1.B [5]);
  nor (_08666_, _08665_, _08664_);
  and (_08667_, _04476_, \oc8051_golden_model_1.PSW [5]);
  not (_08668_, _08667_);
  and (_08669_, _04481_, \oc8051_golden_model_1.IP [5]);
  and (_08670_, _04483_, \oc8051_golden_model_1.ACC [5]);
  nor (_08671_, _08670_, _08669_);
  and (_08672_, _08671_, _08668_);
  and (_08673_, _08672_, _08666_);
  and (_08674_, _04471_, \oc8051_golden_model_1.SCON [5]);
  and (_08675_, _04473_, \oc8051_golden_model_1.IE [5]);
  nor (_08676_, _08675_, _08674_);
  and (_08677_, _03825_, \oc8051_golden_model_1.P0INREG [5]);
  and (_08678_, _04492_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_08679_, _08678_, _08677_);
  and (_08680_, _04489_, \oc8051_golden_model_1.P1INREG [5]);
  and (_08681_, _04467_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_08682_, _08681_, _08680_);
  and (_08683_, _08682_, _08679_);
  and (_08684_, _08683_, _08676_);
  and (_08685_, _08684_, _08673_);
  and (_08686_, _08685_, _04058_);
  nor (_08687_, _08686_, _08663_);
  nor (_08688_, _08687_, _08661_);
  and (_08689_, _08688_, _08636_);
  and (_08690_, _08689_, _08584_);
  or (_08691_, _08690_, _08505_);
  nor (_08692_, _02246_, _02171_);
  nor (_08693_, _02141_, _01749_);
  not (_08694_, _08693_);
  and (_08695_, _08694_, _02229_);
  and (_08696_, _04650_, _03838_);
  nor (_08697_, _08696_, _08484_);
  and (_08698_, _08697_, _02158_);
  and (_08699_, _03838_, \oc8051_golden_model_1.ACC [7]);
  nor (_08700_, _08699_, _08484_);
  or (_08701_, _08700_, _02063_);
  or (_08702_, _02062_, _06707_);
  and (_08703_, _08702_, _03006_);
  and (_08704_, _08703_, _08701_);
  or (_08705_, _08704_, _06823_);
  or (_08706_, _08705_, _08698_);
  nor (_08707_, _01774_, _01744_);
  not (_08708_, _08707_);
  nor (_08709_, _06828_, \oc8051_golden_model_1.PSW [7]);
  not (_08710_, _08709_);
  nor (_08711_, _08710_, _06838_);
  not (_08712_, _08711_);
  nand (_08713_, _08712_, _06823_);
  and (_08714_, _08713_, _08708_);
  and (_08715_, _08714_, _02058_);
  and (_08716_, _08715_, _08706_);
  nor (_08717_, _04476_, _06707_);
  not (_08718_, _08717_);
  nand (_08719_, _04521_, _04476_);
  and (_08720_, _08719_, _08718_);
  and (_08721_, _08720_, _02057_);
  or (_08722_, _08721_, _08716_);
  or (_08723_, _08722_, _02155_);
  or (_08724_, _08494_, _02519_);
  and (_08725_, _08724_, _02549_);
  and (_08726_, _08725_, _08723_);
  and (_08727_, _08700_, _02153_);
  nor (_08728_, _01774_, _01756_);
  or (_08729_, _08728_, _02053_);
  or (_08730_, _08729_, _08727_);
  or (_08731_, _08730_, _08726_);
  and (_08732_, _04517_, _04476_);
  nor (_08733_, _08732_, _08717_);
  or (_08734_, _08733_, _02054_);
  nand (_08735_, _08734_, _08731_);
  nand (_08736_, _08735_, _08695_);
  and (_08737_, _03796_, _01952_);
  not (_08738_, _08737_);
  and (_08739_, _08738_, _03797_);
  and (_08740_, _03964_, _02118_);
  nor (_08741_, _03964_, _02118_);
  or (_08742_, _08741_, _08740_);
  and (_08743_, _08742_, _08739_);
  nor (_08744_, _04057_, _03810_);
  and (_08745_, _04057_, _03810_);
  nor (_08746_, _08745_, _08744_);
  and (_08747_, _04372_, _02825_);
  nor (_08748_, _04372_, _02825_);
  or (_08749_, _08748_, _08747_);
  and (_08750_, _08749_, _08746_);
  and (_08751_, _08750_, _08743_);
  and (_08752_, _03020_, _02028_);
  not (_08753_, _08752_);
  nor (_08754_, _03624_, _02453_);
  not (_08755_, _08754_);
  and (_08756_, _03624_, _02453_);
  not (_08757_, _08756_);
  and (_08758_, _03434_, _02120_);
  nor (_08759_, _03434_, _02120_);
  nor (_08760_, _08759_, _08758_);
  and (_08761_, _08760_, _08757_);
  and (_08762_, _08761_, _08755_);
  nor (_08763_, _03161_, _02860_);
  and (_08764_, _03002_, _02027_);
  and (_08765_, _03161_, _02860_);
  or (_08766_, _08765_, _08764_);
  nor (_08767_, _08766_, _08763_);
  and (_08768_, _08767_, _08762_);
  and (_08769_, _08768_, _08753_);
  and (_08770_, _08769_, _08751_);
  or (_08771_, _08767_, _08765_);
  nand (_08772_, _08771_, _08762_);
  nor (_08773_, _08757_, _08759_);
  nor (_08774_, _08773_, _08758_);
  nand (_08775_, _08774_, _08772_);
  nand (_08776_, _08775_, _08751_);
  and (_08777_, _04372_, _03799_);
  and (_08778_, _08746_, _08777_);
  or (_08779_, _08778_, _08745_);
  nand (_08780_, _08779_, _08743_);
  and (_08781_, _03964_, _03495_);
  nand (_08782_, _08739_, _08781_);
  and (_08783_, _08782_, _08738_);
  and (_08784_, _08783_, _08780_);
  and (_08785_, _08784_, _08776_);
  or (_08786_, _08785_, _08770_);
  or (_08787_, _08786_, _08695_);
  and (_08788_, _08787_, _02233_);
  and (_08789_, _08788_, _08736_);
  and (_08790_, _02030_, _02045_);
  and (_08791_, _08786_, _02232_);
  or (_08792_, _08791_, _08790_);
  or (_08793_, _08792_, _08789_);
  or (_08794_, _05166_, _01983_);
  or (_08795_, _05211_, _02452_);
  and (_08796_, _05166_, _01983_);
  or (_08797_, _08796_, _08795_);
  and (_08798_, _08797_, _08794_);
  or (_08799_, _05075_, _02859_);
  and (_08800_, _05120_, _02027_);
  or (_08801_, _05075_, _02860_);
  nand (_08802_, _05075_, _02860_);
  and (_08803_, _08802_, _08801_);
  or (_08804_, _08803_, _08800_);
  nand (_08805_, _08804_, _08799_);
  not (_08806_, _08796_);
  and (_08807_, _08806_, _08794_);
  nand (_08808_, _05211_, _02452_);
  and (_08809_, _08808_, _08807_);
  and (_08810_, _08809_, _08795_);
  nand (_08811_, _08810_, _08805_);
  nand (_08812_, _08811_, _08798_);
  or (_08813_, _05303_, _02825_);
  or (_08814_, _05258_, _02410_);
  nand (_08815_, _05258_, _02410_);
  and (_08816_, _08815_, _08814_);
  and (_08817_, _08816_, _08813_);
  nand (_08818_, _05303_, _02825_);
  nand (_08819_, _05029_, _02118_);
  or (_08820_, _05029_, _02118_);
  or (_08821_, _04637_, _03835_);
  and (_08822_, _08821_, _04699_);
  and (_08823_, _08822_, _08820_);
  and (_08824_, _08823_, _08819_);
  and (_08825_, _08824_, _08818_);
  and (_08826_, _08825_, _08817_);
  nand (_08827_, _08826_, _08812_);
  nand (_08828_, _08813_, _08814_);
  and (_08829_, _08824_, _08828_);
  nand (_08830_, _08829_, _08815_);
  not (_08831_, _04699_);
  or (_08832_, _08820_, _08831_);
  and (_08833_, _08832_, _08821_);
  and (_08834_, _08833_, _08830_);
  and (_08835_, _08834_, _08827_);
  not (_08836_, _08790_);
  or (_08837_, _05120_, _02028_);
  nand (_08838_, _05120_, _02028_);
  and (_08839_, _08838_, _08837_);
  nor (_08840_, _08803_, _08839_);
  and (_08841_, _08840_, _08810_);
  and (_08842_, _08841_, _08826_);
  or (_08843_, _08842_, _08836_);
  or (_08844_, _08843_, _08835_);
  nand (_08845_, _08844_, _08793_);
  nand (_08846_, _08845_, _08692_);
  nor (_08847_, _07056_, \oc8051_golden_model_1.ACC [3]);
  and (_08848_, _07056_, \oc8051_golden_model_1.ACC [3]);
  nor (_08849_, _08848_, _08847_);
  and (_08850_, _08849_, _07509_);
  not (_08851_, _07189_);
  and (_08852_, _07094_, \oc8051_golden_model_1.ACC [0]);
  nor (_08853_, _08852_, _08851_);
  or (_08854_, _08853_, _07187_);
  nand (_08855_, _08854_, _08850_);
  and (_08856_, _08849_, _07508_);
  nor (_08857_, _08856_, _08847_);
  nand (_08858_, _08857_, _08855_);
  and (_08859_, _07500_, _07504_);
  not (_08860_, _07492_);
  and (_08861_, _08860_, _07496_);
  and (_08862_, _08861_, _08859_);
  nand (_08863_, _08862_, _08858_);
  and (_08864_, _07500_, _07503_);
  or (_08865_, _08864_, _07498_);
  nand (_08866_, _08865_, _08861_);
  or (_08867_, _04682_, \oc8051_golden_model_1.ACC [7]);
  nand (_08868_, _08860_, _07495_);
  and (_08870_, _08868_, _08867_);
  and (_08871_, _08870_, _08866_);
  and (_08872_, _08871_, _08863_);
  nor (_08873_, _07094_, \oc8051_golden_model_1.ACC [0]);
  nor (_08874_, _08852_, _08873_);
  and (_08875_, _08874_, _07189_);
  and (_08876_, _08875_, _08850_);
  and (_08877_, _08862_, _08876_);
  or (_08878_, _08877_, _02547_);
  or (_08879_, _08878_, _08872_);
  nor (_08881_, _01774_, _01749_);
  not (_08882_, _08881_);
  nor (_08883_, _07544_, _07545_);
  nor (_08884_, _08883_, _07548_);
  or (_08885_, _02859_, \oc8051_golden_model_1.ACC [1]);
  and (_08886_, _02859_, \oc8051_golden_model_1.ACC [1]);
  and (_08887_, _02027_, \oc8051_golden_model_1.ACC [0]);
  or (_08888_, _08887_, _08886_);
  nand (_08889_, _08888_, _08885_);
  nand (_08890_, _08889_, _08884_);
  and (_08892_, _01983_, \oc8051_golden_model_1.ACC [3]);
  nor (_08893_, _01983_, \oc8051_golden_model_1.ACC [3]);
  nor (_08894_, _02452_, \oc8051_golden_model_1.ACC [2]);
  nor (_08895_, _08894_, _08893_);
  or (_08896_, _08895_, _08892_);
  nand (_08897_, _08896_, _08890_);
  not (_08898_, _07543_);
  and (_08899_, _07540_, _08898_);
  nor (_08900_, _07537_, _07280_);
  and (_08901_, _08900_, _08899_);
  nand (_08903_, _08901_, _08897_);
  and (_08904_, _02410_, \oc8051_golden_model_1.ACC [5]);
  nor (_08905_, _02410_, \oc8051_golden_model_1.ACC [5]);
  nor (_08906_, _02825_, \oc8051_golden_model_1.ACC [4]);
  nor (_08907_, _08906_, _08905_);
  nor (_08908_, _08907_, _08904_);
  nand (_08909_, _08900_, _08908_);
  nand (_08910_, _01952_, _04939_);
  or (_08911_, _02118_, \oc8051_golden_model_1.ACC [6]);
  or (_08912_, _08911_, _07280_);
  and (_08914_, _08912_, _08910_);
  and (_08915_, _08914_, _08909_);
  and (_08916_, _08915_, _08903_);
  not (_08917_, _02246_);
  and (_08918_, _02027_, _01887_);
  nor (_08919_, _08918_, _07553_);
  nor (_08920_, _08919_, _07552_);
  and (_08921_, _08920_, _08884_);
  and (_08922_, _08901_, _08921_);
  or (_08923_, _08922_, _08917_);
  or (_08925_, _08923_, _08916_);
  and (_08926_, _08925_, _08882_);
  and (_08927_, _08926_, _08879_);
  and (_08928_, _08927_, _08846_);
  and (_08929_, _08881_, \oc8051_golden_model_1.PSW [7]);
  or (_08930_, _08929_, _02046_);
  or (_08931_, _08930_, _08928_);
  and (_08932_, _08718_, _04686_);
  or (_08933_, _08720_, _02047_);
  or (_08934_, _08933_, _08932_);
  and (_08936_, _08934_, _08931_);
  or (_08937_, _08936_, _02147_);
  and (_08938_, _04467_, \oc8051_golden_model_1.P3 [2]);
  not (_08939_, _08938_);
  and (_08940_, _04492_, \oc8051_golden_model_1.P2 [2]);
  nor (_08941_, _08940_, _08523_);
  and (_08942_, _08941_, _08939_);
  and (_08943_, _03825_, \oc8051_golden_model_1.P0 [2]);
  and (_08944_, _04489_, \oc8051_golden_model_1.P1 [2]);
  nor (_08945_, _08944_, _08943_);
  and (_08946_, _08945_, _08522_);
  and (_08947_, _08946_, _08942_);
  and (_08948_, _08947_, _08513_);
  and (_08949_, _08948_, _04259_);
  nor (_08950_, _08949_, _08506_);
  and (_08951_, _03825_, \oc8051_golden_model_1.P0 [1]);
  and (_08952_, _04489_, \oc8051_golden_model_1.P1 [1]);
  nor (_08953_, _08952_, _08951_);
  and (_08954_, _04467_, \oc8051_golden_model_1.P3 [1]);
  and (_08955_, _04492_, \oc8051_golden_model_1.P2 [1]);
  or (_08956_, _08955_, _08954_);
  nor (_08957_, _08956_, _08535_);
  and (_08958_, _08957_, _08545_);
  and (_08959_, _08958_, _08534_);
  and (_08960_, _08959_, _08953_);
  and (_08961_, _08960_, _04154_);
  nor (_08962_, _08961_, _08531_);
  nor (_08963_, _08962_, _08950_);
  and (_08964_, _04492_, \oc8051_golden_model_1.P2 [4]);
  and (_08965_, _04467_, \oc8051_golden_model_1.P3 [4]);
  nor (_08966_, _08965_, _08964_);
  and (_08967_, _03825_, \oc8051_golden_model_1.P0 [4]);
  and (_08968_, _04489_, \oc8051_golden_model_1.P1 [4]);
  nor (_08969_, _08968_, _08967_);
  and (_08970_, _08969_, _08966_);
  and (_08971_, _08970_, _08570_);
  and (_08972_, _08971_, _08567_);
  and (_08973_, _08972_, _04373_);
  nor (_08974_, _08557_, _08973_);
  nor (_08975_, _08974_, _04686_);
  and (_08976_, _08975_, _08963_);
  and (_08977_, _04492_, \oc8051_golden_model_1.P2 [0]);
  and (_08978_, _04467_, \oc8051_golden_model_1.P3 [0]);
  nor (_08979_, _08978_, _08977_);
  and (_08980_, _03825_, \oc8051_golden_model_1.P0 [0]);
  and (_08981_, _04489_, \oc8051_golden_model_1.P1 [0]);
  nor (_08982_, _08981_, _08980_);
  and (_08983_, _08982_, _08979_);
  and (_08984_, _08983_, _08598_);
  and (_08985_, _08984_, _08595_);
  and (_08986_, _08985_, _04210_);
  nor (_08987_, _08986_, _08585_);
  and (_08988_, _04492_, \oc8051_golden_model_1.P2 [6]);
  and (_08989_, _04467_, \oc8051_golden_model_1.P3 [6]);
  nor (_08990_, _08989_, _08988_);
  and (_08991_, _03825_, \oc8051_golden_model_1.P0 [6]);
  and (_08992_, _04489_, \oc8051_golden_model_1.P1 [6]);
  nor (_08993_, _08992_, _08991_);
  and (_08994_, _08993_, _08990_);
  and (_08995_, _08994_, _08624_);
  and (_08996_, _08995_, _08621_);
  and (_08997_, _08996_, _03965_);
  nor (_08998_, _08611_, _08997_);
  nor (_08999_, _08998_, _08987_);
  and (_09000_, _04492_, \oc8051_golden_model_1.P2 [3]);
  and (_09001_, _04467_, \oc8051_golden_model_1.P3 [3]);
  nor (_09002_, _09001_, _09000_);
  and (_09003_, _03825_, \oc8051_golden_model_1.P0 [3]);
  and (_09004_, _04489_, \oc8051_golden_model_1.P1 [3]);
  nor (_09005_, _09004_, _09003_);
  and (_09006_, _09005_, _09002_);
  and (_09007_, _09006_, _08650_);
  and (_09008_, _09007_, _08647_);
  and (_09009_, _09008_, _04105_);
  nor (_09010_, _09009_, _08637_);
  and (_09011_, _04492_, \oc8051_golden_model_1.P2 [5]);
  and (_09012_, _04467_, \oc8051_golden_model_1.P3 [5]);
  nor (_09013_, _09012_, _09011_);
  and (_09014_, _03825_, \oc8051_golden_model_1.P0 [5]);
  and (_09015_, _04489_, \oc8051_golden_model_1.P1 [5]);
  nor (_09016_, _09015_, _09014_);
  and (_09017_, _09016_, _09013_);
  and (_09018_, _09017_, _08676_);
  and (_09019_, _09018_, _08673_);
  and (_09020_, _09019_, _04058_);
  nor (_09021_, _08663_, _09020_);
  nor (_09022_, _09021_, _09010_);
  and (_09023_, _09022_, _08999_);
  and (_09024_, _09023_, _08976_);
  and (_09025_, _02147_, \oc8051_golden_model_1.PSW [7]);
  nand (_09026_, _09025_, _09024_);
  and (_09027_, _09026_, _08937_);
  or (_09028_, _05474_, _02182_);
  or (_09029_, _09028_, _09027_);
  and (_09030_, _09029_, _08691_);
  or (_09031_, _09030_, _02181_);
  not (_09032_, _02181_);
  nor (_09033_, _09024_, \oc8051_golden_model_1.PSW [7]);
  or (_09034_, _09033_, _09032_);
  and (_09035_, _02133_, _01766_);
  not (_09036_, _09035_);
  and (_09037_, _02129_, _02235_);
  nor (_09038_, _09037_, _02137_);
  nor (_09039_, _09038_, _01777_);
  nor (_09040_, _09039_, _02628_);
  and (_09041_, _09040_, _09036_);
  and (_09042_, _09041_, _09034_);
  and (_09043_, _09042_, _09031_);
  and (_09044_, _06667_, _06663_);
  nor (_09045_, _09044_, _06661_);
  not (_09046_, _09045_);
  and (_09047_, _06669_, _06663_);
  not (_09048_, _09047_);
  nor (_09049_, _09048_, _06932_);
  nor (_09050_, _09049_, _09046_);
  nor (_09051_, _09050_, _08470_);
  or (_09052_, _09051_, _02625_);
  and (_09053_, _09052_, _06817_);
  or (_09054_, _09053_, _09043_);
  or (_09055_, _09051_, _02626_);
  and (_09056_, _09055_, _06941_);
  and (_09057_, _09056_, _09054_);
  or (_09058_, _09057_, _08504_);
  and (_09059_, _09058_, _02191_);
  and (_09060_, _07139_, _07135_);
  nor (_09061_, _09060_, _07133_);
  not (_09062_, _09061_);
  and (_09063_, _07388_, _07135_);
  not (_09064_, _09063_);
  nor (_09065_, _09064_, _07201_);
  nor (_09066_, _09065_, _09062_);
  not (_09067_, _04682_);
  and (_09068_, _07129_, _09067_);
  or (_09069_, _09068_, _02191_);
  nor (_09070_, _09069_, _09066_);
  or (_09071_, _09070_, _06740_);
  or (_09072_, _09071_, _09059_);
  and (_09073_, _06743_, _03846_);
  and (_09074_, _06757_, _06751_);
  and (_09075_, _09074_, _06805_);
  and (_09076_, _09074_, _06807_);
  not (_09077_, _09076_);
  and (_09078_, _06755_, _06751_);
  nor (_09079_, _09078_, _06749_);
  and (_09080_, _09079_, _09077_);
  not (_09081_, _09080_);
  nor (_09082_, _09081_, _09075_);
  nor (_09083_, _09082_, _09073_);
  or (_09084_, _09083_, _06741_);
  and (_09085_, _09084_, _05444_);
  and (_09086_, _09085_, _09072_);
  or (_09087_, _09086_, _08495_);
  and (_09088_, _09087_, _02032_);
  or (_09089_, _04698_, _08489_);
  nor (_09090_, _08484_, _02032_);
  and (_09091_, _09090_, _09089_);
  or (_09092_, _09091_, _01765_);
  or (_09093_, _09092_, _09088_);
  and (_09094_, _09093_, _08492_);
  or (_09095_, _06202_, _02124_);
  or (_09096_, _09095_, _09094_);
  nand (_09097_, _02124_, \oc8051_golden_model_1.PSW [7]);
  or (_09098_, _09097_, _09024_);
  and (_09099_, _09098_, _01995_);
  and (_09100_, _09099_, _09096_);
  and (_09101_, _04716_, _03838_);
  nor (_09102_, _09101_, _08484_);
  and (_09103_, _09102_, _01994_);
  or (_09104_, _09103_, _09100_);
  and (_09105_, _09104_, _02688_);
  and (_09106_, _09024_, _06707_);
  and (_09107_, _09106_, _02123_);
  or (_09108_, _09107_, _09105_);
  and (_09109_, _09108_, _03059_);
  nand (_09110_, _04933_, _03838_);
  nor (_09111_, _08484_, _03059_);
  and (_09112_, _09111_, _09110_);
  or (_09113_, _09112_, _02331_);
  or (_09114_, _09113_, _09109_);
  and (_09115_, _09114_, _08488_);
  or (_09116_, _09115_, _02206_);
  and (_09117_, _08485_, _03902_);
  or (_09118_, _09102_, _02208_);
  or (_09119_, _09118_, _09117_);
  and (_09120_, _09119_, _09116_);
  or (_09121_, _09120_, _02342_);
  or (_09122_, _08700_, _03065_);
  or (_09123_, _09122_, _09117_);
  and (_09124_, _09123_, _04953_);
  and (_09125_, _09124_, _09121_);
  or (_09126_, _04932_, _08489_);
  nor (_09127_, _08484_, _04953_);
  and (_09128_, _09127_, _09126_);
  or (_09129_, _09128_, _02334_);
  or (_09130_, _09129_, _09125_);
  or (_09131_, _04940_, _08489_);
  and (_09132_, _09131_, _08485_);
  or (_09133_, _09132_, _04958_);
  and (_09134_, _09133_, _06729_);
  and (_09135_, _09134_, _09130_);
  or (_09136_, _09135_, _08482_);
  or (_09137_, _08478_, _06728_);
  and (_09138_, _09137_, _07356_);
  and (_09139_, _09138_, _09136_);
  or (_09140_, _09139_, _08468_);
  nor (_09141_, _09140_, _02345_);
  nor (_09142_, _07132_, _04939_);
  or (_09143_, _09142_, _07409_);
  nor (_09144_, _09143_, _09068_);
  nor (_09145_, _09144_, _02346_);
  or (_09146_, _09145_, _09141_);
  nor (_09147_, _09146_, _07384_);
  nor (_09148_, _06748_, _04939_);
  nor (_09149_, _09148_, _07437_);
  nor (_09150_, _09073_, _07417_);
  and (_09151_, _09150_, _09149_);
  nor (_09152_, _09151_, _07415_);
  not (_09153_, _09152_);
  nor (_09154_, _09153_, _09147_);
  not (_09155_, _06614_);
  and (_09156_, _07415_, \oc8051_golden_model_1.ACC [7]);
  nor (_09157_, _09156_, _09155_);
  not (_09158_, _09157_);
  nor (_09159_, _09158_, _09154_);
  nor (_09160_, _09159_, _08462_);
  nor (_09161_, _09160_, _06609_);
  not (_09162_, _07270_);
  nor (_09163_, _07480_, _07269_);
  nor (_09164_, _09163_, _07448_);
  and (_09165_, _09164_, _09162_);
  nor (_09166_, _09165_, _02085_);
  not (_09167_, _09166_);
  nor (_09168_, _09167_, _09161_);
  not (_09169_, _07491_);
  and (_09170_, _07526_, _09169_);
  nor (_09171_, _09170_, _07490_);
  and (_09172_, _09171_, _02085_);
  or (_09173_, _09172_, _09168_);
  and (_09174_, _09173_, _08458_);
  not (_09175_, _07278_);
  not (_09176_, _07279_);
  nand (_09177_, _07565_, _09176_);
  and (_09178_, _09177_, _09175_);
  and (_09179_, _09178_, _07487_);
  or (_09180_, _09179_, _09174_);
  nor (_09181_, _09180_, _02366_);
  and (_09182_, _08697_, _02366_);
  nor (_09183_, _09182_, _07580_);
  not (_09184_, _09183_);
  nor (_09185_, _09184_, _09181_);
  and (_09186_, _07580_, \oc8051_golden_model_1.ACC [0]);
  or (_09187_, _09186_, _09185_);
  and (_09188_, _09187_, _01698_);
  nor (_09189_, _08733_, _01698_);
  or (_09190_, _09189_, _09188_);
  nor (_09191_, _09190_, _02081_);
  and (_09192_, _04426_, _03838_);
  nor (_09193_, _09192_, _08484_);
  and (_09194_, _09193_, _02081_);
  nor (_09195_, _09194_, _09191_);
  or (_09196_, _09195_, _39633_);
  or (_09197_, _39632_, \oc8051_golden_model_1.PSW [7]);
  and (_09198_, _09197_, _39026_);
  and (_38594_, _09198_, _09196_);
  not (_09199_, \oc8051_golden_model_1.PCON [7]);
  nor (_09200_, _03828_, _09199_);
  not (_09201_, _03828_);
  nor (_09202_, _04940_, _09201_);
  nor (_09203_, _09202_, _09200_);
  nor (_09204_, _09203_, _04958_);
  and (_09205_, _04942_, _03828_);
  nor (_09206_, _09205_, _09200_);
  nor (_09207_, _09206_, _03061_);
  and (_09208_, _04637_, _03828_);
  or (_09209_, _09208_, _09200_);
  and (_09210_, _09209_, _02031_);
  and (_09211_, _03828_, \oc8051_golden_model_1.ACC [7]);
  nor (_09212_, _09211_, _09200_);
  nor (_09213_, _09212_, _02063_);
  nor (_09214_, _02062_, _09199_);
  or (_09215_, _09214_, _09213_);
  and (_09216_, _09215_, _03006_);
  and (_09217_, _04650_, _03828_);
  nor (_09218_, _09217_, _09200_);
  nor (_09219_, _09218_, _03006_);
  or (_09220_, _09219_, _09216_);
  and (_09221_, _09220_, _02519_);
  nor (_09222_, _09201_, _03796_);
  nor (_09223_, _09222_, _09200_);
  nor (_09224_, _09223_, _02519_);
  nor (_09225_, _09224_, _09221_);
  nor (_09226_, _09225_, _02153_);
  nor (_09227_, _09212_, _02549_);
  nor (_09228_, _09227_, _06188_);
  not (_09229_, _09228_);
  nor (_09230_, _09229_, _09226_);
  and (_09231_, _09223_, _06188_);
  or (_09232_, _09231_, _02031_);
  nor (_09233_, _09232_, _09230_);
  or (_09234_, _09233_, _09210_);
  and (_09235_, _09234_, _02037_);
  nor (_09236_, _04910_, _09201_);
  nor (_09237_, _09236_, _09200_);
  nor (_09238_, _09237_, _02037_);
  or (_09239_, _09238_, _07629_);
  or (_09240_, _09239_, _09235_);
  and (_09241_, _04933_, _03828_);
  or (_09242_, _09200_, _03059_);
  or (_09243_, _09242_, _09241_);
  and (_09244_, _04716_, _03828_);
  nor (_09245_, _09244_, _09200_);
  and (_09246_, _09245_, _01994_);
  nor (_09247_, _09246_, _02331_);
  and (_09248_, _09247_, _09243_);
  and (_09249_, _09248_, _09240_);
  nor (_09250_, _09249_, _09207_);
  nor (_09251_, _09250_, _02206_);
  nor (_09252_, _09200_, _03903_);
  not (_09253_, _09252_);
  nor (_09254_, _09245_, _02208_);
  and (_09255_, _09254_, _09253_);
  nor (_09256_, _09255_, _09251_);
  nor (_09257_, _09256_, _02342_);
  or (_09258_, _09252_, _03065_);
  nor (_09259_, _09258_, _09212_);
  or (_09260_, _09259_, _02202_);
  nor (_09261_, _09260_, _09257_);
  nor (_09262_, _04932_, _09201_);
  or (_09263_, _09200_, _04953_);
  nor (_09264_, _09263_, _09262_);
  or (_09265_, _09264_, _02334_);
  nor (_09266_, _09265_, _09261_);
  nor (_09267_, _09266_, _09204_);
  nor (_09268_, _09267_, _02366_);
  nor (_09269_, _09218_, _02778_);
  or (_09270_, _09269_, _02081_);
  nor (_09271_, _09270_, _09268_);
  and (_09272_, _04426_, _03828_);
  nor (_09273_, _09272_, _09200_);
  and (_09274_, _09273_, _02081_);
  nor (_09275_, _09274_, _09271_);
  or (_09276_, _09275_, _39633_);
  or (_09277_, _39632_, \oc8051_golden_model_1.PCON [7]);
  and (_09278_, _09277_, _39026_);
  and (_38595_, _09278_, _09276_);
  not (_09279_, \oc8051_golden_model_1.SBUF [7]);
  nor (_09280_, _03805_, _09279_);
  not (_09281_, _03805_);
  nor (_09282_, _04940_, _09281_);
  nor (_09283_, _09282_, _09280_);
  nor (_09284_, _09283_, _04958_);
  and (_09285_, _04942_, _03805_);
  nor (_09286_, _09285_, _09280_);
  nor (_09287_, _09286_, _03061_);
  and (_09288_, _04637_, _03805_);
  or (_09289_, _09288_, _09280_);
  and (_09290_, _09289_, _02031_);
  and (_09291_, _03805_, \oc8051_golden_model_1.ACC [7]);
  nor (_09292_, _09291_, _09280_);
  nor (_09293_, _09292_, _02549_);
  nor (_09294_, _09292_, _02063_);
  nor (_09295_, _02062_, _09279_);
  or (_09296_, _09295_, _09294_);
  and (_09297_, _09296_, _03006_);
  and (_09298_, _04650_, _03805_);
  nor (_09299_, _09298_, _09280_);
  nor (_09300_, _09299_, _03006_);
  or (_09301_, _09300_, _09297_);
  and (_09302_, _09301_, _02519_);
  nor (_09303_, _09281_, _03796_);
  nor (_09304_, _09303_, _09280_);
  nor (_09305_, _09304_, _02519_);
  nor (_09306_, _09305_, _09302_);
  nor (_09307_, _09306_, _02153_);
  or (_09308_, _09307_, _06188_);
  nor (_09309_, _09308_, _09293_);
  and (_09310_, _09304_, _06188_);
  or (_09311_, _09310_, _02031_);
  nor (_09312_, _09311_, _09309_);
  or (_09313_, _09312_, _09290_);
  and (_09314_, _09313_, _02037_);
  nor (_09315_, _04910_, _09281_);
  nor (_09316_, _09315_, _09280_);
  nor (_09317_, _09316_, _02037_);
  or (_09318_, _09317_, _07629_);
  or (_09319_, _09318_, _09314_);
  and (_09320_, _04933_, _03805_);
  or (_09321_, _09280_, _03059_);
  or (_09322_, _09321_, _09320_);
  and (_09323_, _04716_, _03805_);
  nor (_09324_, _09323_, _09280_);
  and (_09325_, _09324_, _01994_);
  nor (_09326_, _09325_, _02331_);
  and (_09327_, _09326_, _09322_);
  and (_09328_, _09327_, _09319_);
  nor (_09329_, _09328_, _09287_);
  nor (_09330_, _09329_, _02206_);
  nor (_09331_, _09280_, _03903_);
  not (_09332_, _09331_);
  nor (_09333_, _09324_, _02208_);
  and (_09334_, _09333_, _09332_);
  nor (_09335_, _09334_, _09330_);
  nor (_09336_, _09335_, _02342_);
  or (_09337_, _09331_, _03065_);
  nor (_09338_, _09337_, _09292_);
  or (_09339_, _09338_, _02202_);
  nor (_09340_, _09339_, _09336_);
  nor (_09341_, _04932_, _09281_);
  or (_09342_, _09280_, _04953_);
  nor (_09343_, _09342_, _09341_);
  or (_09344_, _09343_, _02334_);
  nor (_09345_, _09344_, _09340_);
  nor (_09346_, _09345_, _09284_);
  nor (_09347_, _09346_, _02366_);
  nor (_09348_, _09299_, _02778_);
  or (_09349_, _09348_, _02081_);
  nor (_09350_, _09349_, _09347_);
  and (_09351_, _04426_, _03805_);
  nor (_09352_, _09351_, _09280_);
  and (_09353_, _09352_, _02081_);
  nor (_09354_, _09353_, _09350_);
  or (_09355_, _09354_, _39633_);
  or (_09356_, _39632_, \oc8051_golden_model_1.SBUF [7]);
  and (_09357_, _09356_, _39026_);
  and (_38596_, _09357_, _09355_);
  not (_09358_, \oc8051_golden_model_1.SCON [7]);
  nor (_09359_, _03868_, _09358_);
  not (_09360_, _03868_);
  nor (_09361_, _09360_, _03796_);
  nor (_09362_, _09361_, _09359_);
  and (_09363_, _09362_, _06188_);
  and (_09364_, _03868_, \oc8051_golden_model_1.ACC [7]);
  nor (_09365_, _09364_, _09359_);
  nor (_09366_, _09365_, _02063_);
  nor (_09367_, _02062_, _09358_);
  or (_09368_, _09367_, _09366_);
  and (_09369_, _09368_, _03006_);
  and (_09370_, _04650_, _03868_);
  nor (_09371_, _09370_, _09359_);
  nor (_09372_, _09371_, _03006_);
  or (_09373_, _09372_, _09369_);
  and (_09374_, _09373_, _02058_);
  nor (_09375_, _04471_, _09358_);
  and (_09376_, _04521_, _04471_);
  nor (_09377_, _09376_, _09375_);
  nor (_09378_, _09377_, _02058_);
  or (_09379_, _09378_, _09374_);
  and (_09380_, _09379_, _02519_);
  nor (_09381_, _09362_, _02519_);
  or (_09382_, _09381_, _09380_);
  and (_09383_, _09382_, _02549_);
  nor (_09384_, _09365_, _02549_);
  or (_09385_, _09384_, _09383_);
  and (_09386_, _09385_, _02054_);
  and (_09387_, _04517_, _04471_);
  nor (_09388_, _09387_, _09375_);
  nor (_09389_, _09388_, _02054_);
  nor (_09390_, _09389_, _09386_);
  nor (_09391_, _09390_, _02046_);
  and (_09392_, _04688_, _04471_);
  nor (_09393_, _09392_, _09375_);
  nor (_09394_, _09393_, _02047_);
  nor (_09395_, _09394_, _09391_);
  nor (_09396_, _09395_, _02042_);
  not (_09397_, _04471_);
  nor (_09398_, _04503_, _09397_);
  nor (_09399_, _09398_, _09375_);
  nor (_09400_, _09399_, _02043_);
  nor (_09401_, _09400_, _06188_);
  not (_09402_, _09401_);
  nor (_09403_, _09402_, _09396_);
  nor (_09404_, _09403_, _09363_);
  nor (_09405_, _09404_, _02031_);
  and (_09406_, _04637_, _03868_);
  nor (_09407_, _09359_, _02032_);
  not (_09408_, _09407_);
  nor (_09409_, _09408_, _09406_);
  nor (_09410_, _09409_, _01765_);
  not (_09411_, _09410_);
  nor (_09412_, _09411_, _09405_);
  nor (_09413_, _04910_, _09360_);
  nor (_09414_, _09413_, _09359_);
  nor (_09415_, _09414_, _02037_);
  or (_09416_, _09415_, _07629_);
  or (_09417_, _09416_, _09412_);
  and (_09418_, _04933_, _03868_);
  or (_09419_, _09359_, _03059_);
  or (_09420_, _09419_, _09418_);
  and (_09421_, _04716_, _03868_);
  nor (_09422_, _09421_, _09359_);
  and (_09423_, _09422_, _01994_);
  nor (_09424_, _09423_, _02331_);
  and (_09425_, _09424_, _09420_);
  and (_09426_, _09425_, _09417_);
  and (_09427_, _04942_, _03868_);
  nor (_09428_, _09427_, _09359_);
  nor (_09429_, _09428_, _03061_);
  nor (_09430_, _09429_, _09426_);
  nor (_09431_, _09430_, _02206_);
  nor (_09432_, _09359_, _03903_);
  not (_09433_, _09432_);
  nor (_09434_, _09422_, _02208_);
  and (_09435_, _09434_, _09433_);
  nor (_09436_, _09435_, _09431_);
  nor (_09437_, _09436_, _02342_);
  or (_09438_, _09432_, _03065_);
  nor (_09439_, _09438_, _09365_);
  or (_09440_, _09439_, _02202_);
  nor (_09441_, _09440_, _09437_);
  nor (_09442_, _04932_, _09360_);
  or (_09443_, _09359_, _04953_);
  nor (_09444_, _09443_, _09442_);
  or (_09445_, _09444_, _02334_);
  nor (_09446_, _09445_, _09441_);
  nor (_09447_, _04940_, _09360_);
  nor (_09448_, _09447_, _09359_);
  nor (_09449_, _09448_, _04958_);
  or (_09450_, _09449_, _09446_);
  and (_09451_, _09450_, _02778_);
  nor (_09452_, _09371_, _02778_);
  or (_09453_, _09452_, _09451_);
  and (_09454_, _09453_, _01698_);
  nor (_09455_, _09388_, _01698_);
  or (_09456_, _09455_, _09454_);
  and (_09457_, _09456_, _02082_);
  and (_09458_, _04426_, _03868_);
  nor (_09459_, _09458_, _09359_);
  nor (_09460_, _09459_, _02082_);
  or (_09461_, _09460_, _09457_);
  or (_09462_, _09461_, _39633_);
  or (_09463_, _39632_, \oc8051_golden_model_1.SCON [7]);
  and (_09464_, _09463_, _39026_);
  and (_38597_, _09464_, _09462_);
  and (_09465_, _03441_, \oc8051_golden_model_1.SP [4]);
  and (_09466_, _09465_, \oc8051_golden_model_1.SP [5]);
  and (_09467_, _09466_, \oc8051_golden_model_1.SP [6]);
  nor (_09468_, _09467_, \oc8051_golden_model_1.SP [7]);
  and (_09469_, _09467_, \oc8051_golden_model_1.SP [7]);
  nor (_09470_, _09469_, _09468_);
  nor (_09471_, _09470_, _01990_);
  not (_09472_, _02350_);
  not (_09473_, \oc8051_golden_model_1.SP [7]);
  nor (_09474_, _04182_, _09473_);
  and (_09475_, _04942_, _04182_);
  nor (_09476_, _09475_, _09474_);
  nor (_09477_, _09476_, _03061_);
  not (_09478_, _03893_);
  nor (_09479_, _09478_, _03796_);
  nor (_09480_, _09479_, _09474_);
  nor (_09481_, _09480_, _05444_);
  or (_09482_, _09481_, _02031_);
  and (_09483_, _09467_, \oc8051_golden_model_1.SP [0]);
  nor (_09484_, _09483_, \oc8051_golden_model_1.SP [7]);
  and (_09485_, _09483_, \oc8051_golden_model_1.SP [7]);
  nor (_09486_, _09485_, _09484_);
  and (_09487_, _09486_, _02052_);
  not (_09488_, _03311_);
  and (_09489_, _04650_, _04182_);
  nor (_09490_, _09489_, _09474_);
  and (_09491_, _09490_, _02158_);
  and (_09492_, _03893_, \oc8051_golden_model_1.ACC [7]);
  nor (_09493_, _09492_, _09474_);
  or (_09494_, _09493_, _02063_);
  nor (_09495_, _02062_, _02060_);
  nand (_09496_, _09495_, \oc8051_golden_model_1.SP [7]);
  not (_09497_, _09470_);
  nor (_09498_, _09497_, _01747_);
  nor (_09499_, _09498_, _02158_);
  and (_09500_, _09499_, _09496_);
  and (_09501_, _09500_, _09494_);
  nor (_09502_, _09501_, _03446_);
  not (_09503_, _09502_);
  nor (_09504_, _09503_, _09491_);
  nor (_09505_, _09497_, _01745_);
  or (_09506_, _09505_, _02155_);
  nor (_09507_, _09506_, _09504_);
  not (_09508_, \oc8051_golden_model_1.SP [6]);
  not (_09509_, \oc8051_golden_model_1.SP [5]);
  not (_09510_, \oc8051_golden_model_1.SP [4]);
  and (_09511_, _04555_, _09510_);
  and (_09512_, _09511_, _09509_);
  and (_09513_, _09512_, _09508_);
  and (_09514_, _09513_, _01986_);
  nor (_09515_, _09514_, _09473_);
  and (_09516_, _09514_, _09473_);
  nor (_09517_, _09516_, _09515_);
  and (_09518_, _09517_, _02155_);
  nor (_09519_, _09518_, _09507_);
  and (_09520_, _09519_, _02549_);
  nor (_09521_, _09493_, _02549_);
  or (_09522_, _09521_, _09520_);
  and (_09523_, _09522_, _03114_);
  or (_09524_, _09523_, _09488_);
  nor (_09525_, _09524_, _09487_);
  nor (_09526_, _09470_, _03311_);
  or (_09527_, _09526_, _06188_);
  nor (_09528_, _09527_, _09525_);
  nor (_09529_, _09528_, _09482_);
  nor (_09530_, _09474_, _02032_);
  not (_09531_, _04182_);
  or (_09532_, _04698_, _09531_);
  and (_09533_, _09532_, _09530_);
  or (_09534_, _09533_, _01765_);
  nor (_09535_, _09534_, _09529_);
  nor (_09536_, _04910_, _09478_);
  nor (_09537_, _09536_, _09474_);
  nor (_09538_, _09537_, _02037_);
  or (_09539_, _09538_, _01994_);
  or (_09540_, _09539_, _09535_);
  and (_09541_, _04716_, _03893_);
  nor (_09542_, _09541_, _09474_);
  nand (_09543_, _09542_, _01994_);
  and (_09544_, _09543_, _09540_);
  nor (_09545_, _09544_, _01718_);
  and (_09546_, _09497_, _01718_);
  nor (_09547_, _09546_, _09545_);
  and (_09548_, _09547_, _03059_);
  and (_09549_, _04933_, _03893_);
  nor (_09550_, _09549_, _09474_);
  nor (_09551_, _09550_, _03059_);
  or (_09552_, _09551_, _09548_);
  and (_09553_, _09552_, _03061_);
  nor (_09554_, _09553_, _09477_);
  nor (_09555_, _09554_, _02206_);
  nor (_09556_, _09474_, _03903_);
  not (_09557_, _09556_);
  nor (_09558_, _09542_, _02208_);
  and (_09559_, _09558_, _09557_);
  nor (_09560_, _09559_, _09555_);
  nor (_09561_, _02342_, _01728_);
  not (_09562_, _09561_);
  nor (_09563_, _09562_, _09560_);
  and (_09564_, _09470_, _01728_);
  or (_09565_, _09556_, _03065_);
  nor (_09566_, _09565_, _09493_);
  or (_09567_, _09566_, _09564_);
  or (_09568_, _09567_, _02202_);
  nor (_09569_, _09568_, _09563_);
  nor (_09570_, _04932_, _09478_);
  nor (_09571_, _09570_, _09474_);
  and (_09572_, _09571_, _02202_);
  nor (_09573_, _09572_, _09569_);
  and (_09574_, _09573_, _04958_);
  nor (_09575_, _04940_, _09478_);
  nor (_09576_, _09575_, _09474_);
  nor (_09577_, _09576_, _04958_);
  or (_09578_, _09577_, _09574_);
  and (_09579_, _09578_, _09472_);
  nor (_09580_, _09513_, \oc8051_golden_model_1.SP [7]);
  and (_09581_, _09513_, \oc8051_golden_model_1.SP [7]);
  nor (_09582_, _09581_, _09580_);
  and (_09583_, _09582_, _02350_);
  or (_09584_, _09583_, _01726_);
  nor (_09585_, _09584_, _09579_);
  and (_09586_, _09497_, _01726_);
  nor (_09587_, _09586_, _09585_);
  and (_09588_, _09587_, _02084_);
  and (_09589_, _09582_, _02083_);
  or (_09590_, _09589_, _09588_);
  and (_09591_, _09590_, _02778_);
  nor (_09592_, _09490_, _02778_);
  nor (_09593_, _09592_, _03537_);
  not (_09594_, _09593_);
  nor (_09595_, _09594_, _09591_);
  nor (_09596_, _09595_, _09471_);
  nor (_09597_, _09596_, _02081_);
  and (_09598_, _04426_, _03893_);
  nor (_09599_, _09598_, _09474_);
  and (_09600_, _09599_, _02081_);
  nor (_09601_, _09600_, _09597_);
  or (_09602_, _09601_, _39633_);
  or (_09603_, _39632_, \oc8051_golden_model_1.SP [7]);
  and (_09604_, _09603_, _39026_);
  and (_38598_, _09604_, _09602_);
  not (_09605_, \oc8051_golden_model_1.TCON [7]);
  nor (_09606_, _03856_, _09605_);
  not (_09607_, _03856_);
  nor (_09608_, _09607_, _03796_);
  nor (_09609_, _09608_, _09606_);
  and (_09610_, _09609_, _06188_);
  and (_09611_, _03856_, \oc8051_golden_model_1.ACC [7]);
  nor (_09612_, _09611_, _09606_);
  nor (_09613_, _09612_, _02063_);
  nor (_09614_, _02062_, _09605_);
  or (_09615_, _09614_, _09613_);
  and (_09616_, _09615_, _03006_);
  and (_09617_, _04650_, _03856_);
  nor (_09618_, _09617_, _09606_);
  nor (_09619_, _09618_, _03006_);
  or (_09620_, _09619_, _09616_);
  and (_09621_, _09620_, _02058_);
  nor (_09622_, _04487_, _09605_);
  and (_09623_, _04521_, _04487_);
  nor (_09624_, _09623_, _09622_);
  nor (_09625_, _09624_, _02058_);
  or (_09626_, _09625_, _09621_);
  and (_09627_, _09626_, _02519_);
  nor (_09628_, _09609_, _02519_);
  or (_09629_, _09628_, _09627_);
  and (_09630_, _09629_, _02549_);
  nor (_09631_, _09612_, _02549_);
  or (_09632_, _09631_, _09630_);
  and (_09633_, _09632_, _02054_);
  and (_09634_, _04517_, _04487_);
  nor (_09635_, _09634_, _09622_);
  nor (_09636_, _09635_, _02054_);
  nor (_09637_, _09636_, _09633_);
  nor (_09638_, _09637_, _02046_);
  nor (_09639_, _09622_, _04687_);
  or (_09640_, _09624_, _02047_);
  nor (_09641_, _09640_, _09639_);
  nor (_09642_, _09641_, _09638_);
  nor (_09643_, _09642_, _02042_);
  not (_09644_, _04487_);
  nor (_09645_, _04503_, _09644_);
  nor (_09646_, _09645_, _09622_);
  nor (_09647_, _09646_, _02043_);
  nor (_09648_, _09647_, _06188_);
  not (_09649_, _09648_);
  nor (_09650_, _09649_, _09643_);
  nor (_09651_, _09650_, _09610_);
  nor (_09652_, _09651_, _02031_);
  and (_09653_, _04637_, _03856_);
  nor (_09654_, _09606_, _02032_);
  not (_09655_, _09654_);
  nor (_09656_, _09655_, _09653_);
  nor (_09657_, _09656_, _01765_);
  not (_09658_, _09657_);
  nor (_09659_, _09658_, _09652_);
  nor (_09660_, _04910_, _09607_);
  nor (_09661_, _09660_, _09606_);
  nor (_09662_, _09661_, _02037_);
  or (_09663_, _09662_, _07629_);
  or (_09664_, _09663_, _09659_);
  and (_09665_, _04933_, _03856_);
  or (_09666_, _09606_, _03059_);
  or (_09667_, _09666_, _09665_);
  and (_09668_, _04716_, _03856_);
  nor (_09669_, _09668_, _09606_);
  and (_09670_, _09669_, _01994_);
  nor (_09671_, _09670_, _02331_);
  and (_09672_, _09671_, _09667_);
  and (_09673_, _09672_, _09664_);
  and (_09674_, _04942_, _03856_);
  nor (_09675_, _09674_, _09606_);
  nor (_09676_, _09675_, _03061_);
  nor (_09677_, _09676_, _09673_);
  nor (_09678_, _09677_, _02206_);
  nor (_09679_, _09606_, _03903_);
  not (_09680_, _09679_);
  nor (_09681_, _09669_, _02208_);
  and (_09682_, _09681_, _09680_);
  nor (_09683_, _09682_, _09678_);
  nor (_09684_, _09683_, _02342_);
  or (_09685_, _09679_, _03065_);
  nor (_09686_, _09685_, _09612_);
  or (_09687_, _09686_, _02202_);
  nor (_09688_, _09687_, _09684_);
  nor (_09689_, _04932_, _09607_);
  or (_09690_, _09606_, _04953_);
  nor (_09691_, _09690_, _09689_);
  or (_09692_, _09691_, _02334_);
  nor (_09693_, _09692_, _09688_);
  nor (_09694_, _04940_, _09607_);
  nor (_09695_, _09694_, _09606_);
  nor (_09696_, _09695_, _04958_);
  or (_09697_, _09696_, _09693_);
  and (_09698_, _09697_, _02778_);
  nor (_09699_, _09618_, _02778_);
  or (_09700_, _09699_, _09698_);
  and (_09701_, _09700_, _01698_);
  nor (_09702_, _09635_, _01698_);
  or (_09703_, _09702_, _09701_);
  and (_09704_, _09703_, _02082_);
  and (_09705_, _04426_, _03856_);
  nor (_09706_, _09705_, _09606_);
  nor (_09707_, _09706_, _02082_);
  or (_09708_, _09707_, _09704_);
  or (_09709_, _09708_, _39633_);
  or (_09710_, _39632_, \oc8051_golden_model_1.TCON [7]);
  and (_09711_, _09710_, _39026_);
  and (_38599_, _09711_, _09709_);
  not (_09712_, \oc8051_golden_model_1.TH0 [7]);
  nor (_09713_, _03854_, _09712_);
  not (_09714_, _03854_);
  nor (_09715_, _04940_, _09714_);
  nor (_09716_, _09715_, _09713_);
  nor (_09717_, _09716_, _04958_);
  and (_09718_, _04942_, _03854_);
  nor (_09719_, _09718_, _09713_);
  nor (_09720_, _09719_, _03061_);
  and (_09721_, _04637_, _03854_);
  or (_09722_, _09721_, _09713_);
  and (_09723_, _09722_, _02031_);
  and (_09724_, _03854_, \oc8051_golden_model_1.ACC [7]);
  nor (_09725_, _09724_, _09713_);
  nor (_09726_, _09725_, _02549_);
  nor (_09727_, _09725_, _02063_);
  nor (_09728_, _02062_, _09712_);
  or (_09729_, _09728_, _09727_);
  and (_09730_, _09729_, _03006_);
  and (_09731_, _04650_, _03854_);
  nor (_09732_, _09731_, _09713_);
  nor (_09733_, _09732_, _03006_);
  or (_09734_, _09733_, _09730_);
  and (_09735_, _09734_, _02519_);
  nor (_09736_, _09714_, _03796_);
  nor (_09737_, _09736_, _09713_);
  nor (_09738_, _09737_, _02519_);
  nor (_09739_, _09738_, _09735_);
  nor (_09740_, _09739_, _02153_);
  or (_09741_, _09740_, _06188_);
  nor (_09742_, _09741_, _09726_);
  and (_09743_, _09737_, _06188_);
  or (_09744_, _09743_, _02031_);
  nor (_09745_, _09744_, _09742_);
  or (_09746_, _09745_, _09723_);
  and (_09747_, _09746_, _02037_);
  nor (_09748_, _04910_, _09714_);
  nor (_09749_, _09748_, _09713_);
  nor (_09750_, _09749_, _02037_);
  or (_09751_, _09750_, _07629_);
  or (_09752_, _09751_, _09747_);
  and (_09753_, _04933_, _03854_);
  or (_09754_, _09713_, _03059_);
  or (_09755_, _09754_, _09753_);
  and (_09756_, _04716_, _03854_);
  nor (_09757_, _09756_, _09713_);
  and (_09758_, _09757_, _01994_);
  nor (_09759_, _09758_, _02331_);
  and (_09760_, _09759_, _09755_);
  and (_09761_, _09760_, _09752_);
  nor (_09762_, _09761_, _09720_);
  nor (_09763_, _09762_, _02206_);
  nor (_09764_, _09713_, _03903_);
  not (_09765_, _09764_);
  nor (_09766_, _09757_, _02208_);
  and (_09767_, _09766_, _09765_);
  nor (_09768_, _09767_, _09763_);
  nor (_09769_, _09768_, _02342_);
  or (_09770_, _09764_, _03065_);
  nor (_09771_, _09770_, _09725_);
  or (_09772_, _09771_, _02202_);
  nor (_09773_, _09772_, _09769_);
  nor (_09774_, _04932_, _09714_);
  or (_09775_, _09713_, _04953_);
  nor (_09776_, _09775_, _09774_);
  or (_09777_, _09776_, _02334_);
  nor (_09778_, _09777_, _09773_);
  nor (_09779_, _09778_, _09717_);
  nor (_09780_, _09779_, _02366_);
  nor (_09781_, _09732_, _02778_);
  or (_09782_, _09781_, _02081_);
  nor (_09783_, _09782_, _09780_);
  and (_09784_, _04426_, _03854_);
  nor (_09785_, _09784_, _09713_);
  and (_09786_, _09785_, _02081_);
  nor (_09787_, _09786_, _09783_);
  or (_09788_, _09787_, _39633_);
  or (_09789_, _39632_, \oc8051_golden_model_1.TH0 [7]);
  and (_09790_, _09789_, _39026_);
  and (_38600_, _09790_, _09788_);
  not (_09791_, \oc8051_golden_model_1.TH1 [7]);
  nor (_09792_, _03871_, _09791_);
  not (_09793_, _03871_);
  nor (_09794_, _04940_, _09793_);
  nor (_09795_, _09794_, _09792_);
  nor (_09796_, _09795_, _04958_);
  nor (_09797_, _09792_, _03903_);
  not (_09798_, _09797_);
  and (_09799_, _04716_, _03871_);
  nor (_09800_, _09799_, _09792_);
  nor (_09801_, _09800_, _02208_);
  and (_09802_, _09801_, _09798_);
  and (_09803_, _04942_, _03871_);
  nor (_09804_, _09803_, _09792_);
  nor (_09805_, _09804_, _03061_);
  and (_09806_, _04637_, _03871_);
  or (_09807_, _09806_, _09792_);
  and (_09808_, _09807_, _02031_);
  and (_09809_, _03871_, \oc8051_golden_model_1.ACC [7]);
  nor (_09810_, _09809_, _09792_);
  nor (_09811_, _09810_, _02549_);
  nor (_09812_, _09810_, _02063_);
  nor (_09813_, _02062_, _09791_);
  or (_09814_, _09813_, _09812_);
  and (_09815_, _09814_, _03006_);
  and (_09816_, _04650_, _03871_);
  nor (_09817_, _09816_, _09792_);
  nor (_09818_, _09817_, _03006_);
  or (_09819_, _09818_, _09815_);
  and (_09820_, _09819_, _02519_);
  nor (_09821_, _09793_, _03796_);
  nor (_09822_, _09821_, _09792_);
  nor (_09823_, _09822_, _02519_);
  nor (_09824_, _09823_, _09820_);
  nor (_09825_, _09824_, _02153_);
  or (_09826_, _09825_, _06188_);
  nor (_09827_, _09826_, _09811_);
  and (_09828_, _09822_, _06188_);
  or (_09829_, _09828_, _02031_);
  nor (_09830_, _09829_, _09827_);
  or (_09831_, _09830_, _09808_);
  and (_09832_, _09831_, _02037_);
  nor (_09833_, _04910_, _09793_);
  nor (_09834_, _09833_, _09792_);
  nor (_09835_, _09834_, _02037_);
  or (_09836_, _09835_, _07629_);
  or (_09837_, _09836_, _09832_);
  and (_09838_, _04933_, _03871_);
  or (_09839_, _09792_, _03059_);
  or (_09840_, _09839_, _09838_);
  and (_09841_, _09800_, _01994_);
  nor (_09842_, _09841_, _02331_);
  and (_09843_, _09842_, _09840_);
  and (_09844_, _09843_, _09837_);
  nor (_09845_, _09844_, _09805_);
  nor (_09846_, _09845_, _02206_);
  nor (_09847_, _09846_, _09802_);
  nor (_09848_, _09847_, _02342_);
  or (_09849_, _09797_, _03065_);
  nor (_09850_, _09849_, _09810_);
  or (_09851_, _09850_, _02202_);
  nor (_09852_, _09851_, _09848_);
  nor (_09853_, _04932_, _09793_);
  or (_09854_, _09792_, _04953_);
  nor (_09855_, _09854_, _09853_);
  or (_09856_, _09855_, _02334_);
  nor (_09857_, _09856_, _09852_);
  nor (_09858_, _09857_, _09796_);
  nor (_09859_, _09858_, _02366_);
  nor (_09860_, _09817_, _02778_);
  or (_09861_, _09860_, _02081_);
  nor (_09862_, _09861_, _09859_);
  and (_09863_, _04426_, _03871_);
  nor (_09864_, _09863_, _09792_);
  and (_09865_, _09864_, _02081_);
  nor (_09866_, _09865_, _09862_);
  or (_09867_, _09866_, _39633_);
  or (_09868_, _39632_, \oc8051_golden_model_1.TH1 [7]);
  and (_09869_, _09868_, _39026_);
  and (_38601_, _09869_, _09867_);
  not (_09870_, \oc8051_golden_model_1.TL0 [7]);
  nor (_09871_, _03876_, _09870_);
  not (_09872_, _03876_);
  nor (_09873_, _04940_, _09872_);
  nor (_09874_, _09873_, _09871_);
  nor (_09875_, _09874_, _04958_);
  and (_09876_, _04942_, _03876_);
  nor (_09877_, _09876_, _09871_);
  nor (_09878_, _09877_, _03061_);
  and (_09879_, _04637_, _03876_);
  or (_09880_, _09879_, _09871_);
  and (_09881_, _09880_, _02031_);
  and (_09882_, _03876_, \oc8051_golden_model_1.ACC [7]);
  nor (_09883_, _09882_, _09871_);
  nor (_09884_, _09883_, _02549_);
  nor (_09885_, _09883_, _02063_);
  nor (_09886_, _02062_, _09870_);
  or (_09887_, _09886_, _09885_);
  and (_09888_, _09887_, _03006_);
  and (_09889_, _04650_, _03876_);
  nor (_09890_, _09889_, _09871_);
  nor (_09891_, _09890_, _03006_);
  or (_09892_, _09891_, _09888_);
  and (_09893_, _09892_, _02519_);
  nor (_09894_, _09872_, _03796_);
  nor (_09895_, _09894_, _09871_);
  nor (_09896_, _09895_, _02519_);
  nor (_09897_, _09896_, _09893_);
  nor (_09898_, _09897_, _02153_);
  or (_09899_, _09898_, _06188_);
  nor (_09900_, _09899_, _09884_);
  and (_09901_, _09895_, _06188_);
  or (_09902_, _09901_, _02031_);
  nor (_09903_, _09902_, _09900_);
  or (_09904_, _09903_, _09881_);
  and (_09905_, _09904_, _02037_);
  nor (_09906_, _04910_, _09872_);
  nor (_09907_, _09906_, _09871_);
  nor (_09908_, _09907_, _02037_);
  or (_09909_, _09908_, _07629_);
  or (_09910_, _09909_, _09905_);
  and (_09911_, _04933_, _03876_);
  or (_09912_, _09871_, _03059_);
  or (_09913_, _09912_, _09911_);
  and (_09914_, _04716_, _03876_);
  nor (_09915_, _09914_, _09871_);
  and (_09916_, _09915_, _01994_);
  nor (_09917_, _09916_, _02331_);
  and (_09918_, _09917_, _09913_);
  and (_09919_, _09918_, _09910_);
  nor (_09920_, _09919_, _09878_);
  nor (_09921_, _09920_, _02206_);
  nor (_09922_, _09871_, _03903_);
  not (_09923_, _09922_);
  nor (_09924_, _09915_, _02208_);
  and (_09925_, _09924_, _09923_);
  nor (_09926_, _09925_, _09921_);
  nor (_09927_, _09926_, _02342_);
  or (_09928_, _09922_, _03065_);
  nor (_09929_, _09928_, _09883_);
  or (_09930_, _09929_, _02202_);
  nor (_09931_, _09930_, _09927_);
  nor (_09932_, _04932_, _09872_);
  or (_09933_, _09871_, _04953_);
  nor (_09934_, _09933_, _09932_);
  or (_09935_, _09934_, _02334_);
  nor (_09936_, _09935_, _09931_);
  nor (_09937_, _09936_, _09875_);
  nor (_09938_, _09937_, _02366_);
  nor (_09939_, _09890_, _02778_);
  or (_09940_, _09939_, _02081_);
  nor (_09941_, _09940_, _09938_);
  and (_09942_, _04426_, _03876_);
  nor (_09943_, _09942_, _09871_);
  and (_09944_, _09943_, _02081_);
  nor (_09945_, _09944_, _09941_);
  or (_09946_, _09945_, _39633_);
  or (_09947_, _39632_, \oc8051_golden_model_1.TL0 [7]);
  and (_09948_, _09947_, _39026_);
  and (_38603_, _09948_, _09946_);
  not (_09949_, \oc8051_golden_model_1.TL1 [7]);
  nor (_09950_, _03864_, _09949_);
  not (_09951_, _04197_);
  nor (_09952_, _04940_, _09951_);
  nor (_09953_, _09952_, _09950_);
  nor (_09954_, _09953_, _04958_);
  nor (_09955_, _09950_, _03903_);
  not (_09956_, _09955_);
  and (_09957_, _04716_, _03864_);
  nor (_09958_, _09957_, _09950_);
  nor (_09959_, _09958_, _02208_);
  and (_09960_, _09959_, _09956_);
  and (_09961_, _04942_, _04197_);
  nor (_09962_, _09961_, _09950_);
  nor (_09963_, _09962_, _03061_);
  and (_09964_, _04637_, _03864_);
  or (_09965_, _09964_, _09950_);
  and (_09966_, _09965_, _02031_);
  and (_09967_, _03864_, \oc8051_golden_model_1.ACC [7]);
  nor (_09968_, _09967_, _09950_);
  nor (_09969_, _09968_, _02549_);
  nor (_09970_, _09968_, _02063_);
  nor (_09971_, _02062_, _09949_);
  or (_09972_, _09971_, _09970_);
  and (_09973_, _09972_, _03006_);
  and (_09974_, _04650_, _04197_);
  nor (_09975_, _09974_, _09950_);
  nor (_09976_, _09975_, _03006_);
  or (_09977_, _09976_, _09973_);
  and (_09978_, _09977_, _02519_);
  nor (_09979_, _09951_, _03796_);
  nor (_09980_, _09979_, _09950_);
  nor (_09981_, _09980_, _02519_);
  nor (_09982_, _09981_, _09978_);
  nor (_09983_, _09982_, _02153_);
  or (_09984_, _09983_, _06188_);
  nor (_09985_, _09984_, _09969_);
  and (_09986_, _09980_, _06188_);
  or (_09987_, _09986_, _02031_);
  nor (_09988_, _09987_, _09985_);
  or (_09989_, _09988_, _09966_);
  and (_09990_, _09989_, _02037_);
  nor (_09991_, _04910_, _09951_);
  nor (_09992_, _09991_, _09950_);
  nor (_09993_, _09992_, _02037_);
  or (_09994_, _09993_, _07629_);
  or (_09995_, _09994_, _09990_);
  and (_09996_, _04933_, _04197_);
  or (_09997_, _09950_, _03059_);
  or (_09998_, _09997_, _09996_);
  and (_09999_, _09958_, _01994_);
  nor (_10000_, _09999_, _02331_);
  and (_10001_, _10000_, _09998_);
  and (_10002_, _10001_, _09995_);
  nor (_10003_, _10002_, _09963_);
  nor (_10004_, _10003_, _02206_);
  nor (_10005_, _10004_, _09960_);
  nor (_10006_, _10005_, _02342_);
  or (_10007_, _09955_, _03065_);
  nor (_10008_, _10007_, _09968_);
  or (_10009_, _10008_, _02202_);
  nor (_10010_, _10009_, _10006_);
  or (_10011_, _04932_, _09951_);
  nor (_10012_, _09950_, _04953_);
  and (_10013_, _10012_, _10011_);
  or (_10014_, _10013_, _02334_);
  nor (_10015_, _10014_, _10010_);
  nor (_10016_, _10015_, _09954_);
  nor (_10017_, _10016_, _02366_);
  nor (_10018_, _09975_, _02778_);
  or (_10019_, _10018_, _02081_);
  nor (_10020_, _10019_, _10017_);
  and (_10021_, _04426_, _03864_);
  nor (_10022_, _10021_, _09950_);
  and (_10023_, _10022_, _02081_);
  nor (_10024_, _10023_, _10020_);
  or (_10025_, _10024_, _39633_);
  or (_10026_, _39632_, \oc8051_golden_model_1.TL1 [7]);
  and (_10027_, _10026_, _39026_);
  and (_38604_, _10027_, _10025_);
  not (_10028_, \oc8051_golden_model_1.TMOD [7]);
  nor (_10029_, _03878_, _10028_);
  not (_10030_, _03878_);
  nor (_10031_, _04940_, _10030_);
  nor (_10032_, _10031_, _10029_);
  nor (_10033_, _10032_, _04958_);
  and (_10034_, _04942_, _03878_);
  nor (_10035_, _10034_, _10029_);
  nor (_10036_, _10035_, _03061_);
  and (_10037_, _04637_, _03878_);
  or (_10038_, _10037_, _10029_);
  and (_10039_, _10038_, _02031_);
  and (_10040_, _03878_, \oc8051_golden_model_1.ACC [7]);
  nor (_10041_, _10040_, _10029_);
  nor (_10042_, _10041_, _02549_);
  nor (_10043_, _10041_, _02063_);
  nor (_10044_, _02062_, _10028_);
  or (_10045_, _10044_, _10043_);
  and (_10046_, _10045_, _03006_);
  and (_10047_, _04650_, _03878_);
  nor (_10048_, _10047_, _10029_);
  nor (_10049_, _10048_, _03006_);
  or (_10050_, _10049_, _10046_);
  and (_10051_, _10050_, _02519_);
  nor (_10052_, _10030_, _03796_);
  nor (_10053_, _10052_, _10029_);
  nor (_10054_, _10053_, _02519_);
  nor (_10055_, _10054_, _10051_);
  nor (_10056_, _10055_, _02153_);
  or (_10057_, _10056_, _06188_);
  nor (_10058_, _10057_, _10042_);
  and (_10059_, _10053_, _06188_);
  or (_10060_, _10059_, _02031_);
  nor (_10061_, _10060_, _10058_);
  or (_10062_, _10061_, _10039_);
  and (_10063_, _10062_, _02037_);
  nor (_10064_, _04910_, _10030_);
  nor (_10065_, _10064_, _10029_);
  nor (_10066_, _10065_, _02037_);
  or (_10067_, _10066_, _07629_);
  or (_10068_, _10067_, _10063_);
  and (_10069_, _04933_, _03878_);
  or (_10070_, _10029_, _03059_);
  or (_10071_, _10070_, _10069_);
  and (_10072_, _04716_, _03878_);
  nor (_10073_, _10072_, _10029_);
  and (_10074_, _10073_, _01994_);
  nor (_10075_, _10074_, _02331_);
  and (_10076_, _10075_, _10071_);
  and (_10077_, _10076_, _10068_);
  nor (_10078_, _10077_, _10036_);
  nor (_10079_, _10078_, _02206_);
  nor (_10080_, _10029_, _03903_);
  not (_10081_, _10080_);
  nor (_10082_, _10073_, _02208_);
  and (_10083_, _10082_, _10081_);
  nor (_10084_, _10083_, _10079_);
  nor (_10085_, _10084_, _02342_);
  or (_10086_, _10080_, _03065_);
  nor (_10087_, _10086_, _10041_);
  or (_10088_, _10087_, _02202_);
  nor (_10089_, _10088_, _10085_);
  nor (_10090_, _04932_, _10030_);
  or (_10091_, _10029_, _04953_);
  nor (_10092_, _10091_, _10090_);
  or (_10093_, _10092_, _02334_);
  nor (_10094_, _10093_, _10089_);
  nor (_10095_, _10094_, _10033_);
  nor (_10096_, _10095_, _02366_);
  nor (_10097_, _10048_, _02778_);
  or (_10098_, _10097_, _02081_);
  nor (_10099_, _10098_, _10096_);
  and (_10100_, _04426_, _03878_);
  nor (_10101_, _10100_, _10029_);
  and (_10102_, _10101_, _02081_);
  nor (_10103_, _10102_, _10099_);
  or (_10104_, _10103_, _39633_);
  or (_10105_, _39632_, \oc8051_golden_model_1.TMOD [7]);
  and (_10106_, _10105_, _39026_);
  and (_38605_, _10106_, _10104_);
  not (_10107_, _01426_);
  and (_10108_, _04539_, _10107_);
  and (_10109_, _10108_, \oc8051_golden_model_1.PC [7]);
  and (_10110_, _10109_, _05397_);
  and (_10111_, _10110_, \oc8051_golden_model_1.PC [11]);
  and (_10112_, _10111_, \oc8051_golden_model_1.PC [12]);
  and (_10113_, _10112_, \oc8051_golden_model_1.PC [13]);
  and (_10114_, _10113_, \oc8051_golden_model_1.PC [14]);
  nor (_10115_, _10114_, \oc8051_golden_model_1.PC [15]);
  and (_10116_, _10114_, \oc8051_golden_model_1.PC [15]);
  nor (_10117_, _10116_, _10115_);
  and (_10118_, _06614_, _07448_);
  or (_10119_, _10118_, _10117_);
  and (_10120_, _06729_, _02731_);
  or (_10121_, _10120_, _10117_);
  and (_10122_, _01735_, _01696_);
  not (_10123_, _10122_);
  nor (_10124_, _02334_, _01736_);
  or (_10125_, _10124_, _05428_);
  and (_10126_, _10125_, _10123_);
  not (_10127_, _07331_);
  and (_10128_, _07325_, _01773_);
  nor (_10129_, _10128_, _02719_);
  not (_10130_, _01735_);
  or (_10131_, _09038_, _10130_);
  and (_10132_, _10131_, _10129_);
  and (_10133_, _10132_, _10127_);
  or (_10134_, _10133_, _10117_);
  nor (_10135_, _07312_, _02340_);
  not (_10136_, _10135_);
  nor (_10137_, _02702_, _07304_);
  nor (_10138_, _07298_, _07292_);
  and (_10139_, _10138_, _10137_);
  or (_10140_, _10139_, _10117_);
  and (_10141_, _09037_, _01721_);
  or (_10142_, _10141_, _02693_);
  not (_10143_, _10142_);
  nor (_10144_, _07258_, _02691_);
  and (_10145_, _10144_, _07251_);
  and (_10146_, _10145_, _10143_);
  and (_10147_, _10146_, _07264_);
  or (_10148_, _10147_, _10117_);
  and (_10149_, _02201_, _01717_);
  not (_10150_, _10149_);
  or (_10151_, _05428_, _04919_);
  and (_10152_, _05412_, _01765_);
  nor (_10153_, _06817_, _06815_);
  or (_10154_, _10153_, _10117_);
  and (_10155_, _01764_, _02128_);
  not (_10156_, _10155_);
  nor (_10157_, _07648_, _05474_);
  and (_10158_, _10157_, _10156_);
  not (_10159_, _10158_);
  and (_10160_, _10159_, _10117_);
  nor (_10161_, _05401_, \oc8051_golden_model_1.PC [14]);
  nor (_10162_, _10161_, _05402_);
  not (_10163_, _10162_);
  nor (_10164_, _10163_, _04458_);
  and (_10165_, _10163_, _04458_);
  nor (_10166_, _10165_, _10164_);
  not (_10167_, _10166_);
  nor (_10168_, _05400_, \oc8051_golden_model_1.PC [13]);
  nor (_10169_, _10168_, _05401_);
  and (_10170_, _10169_, _04716_);
  nor (_10171_, _10169_, _04716_);
  nor (_10172_, _05399_, \oc8051_golden_model_1.PC [12]);
  nor (_10173_, _10172_, _05400_);
  not (_10174_, _10173_);
  nor (_10175_, _10174_, _04458_);
  not (_10176_, \oc8051_golden_model_1.PC [11]);
  nor (_10177_, _05398_, _10176_);
  and (_10178_, _05398_, _10176_);
  or (_10179_, _10178_, _10177_);
  not (_10180_, _10179_);
  nor (_10181_, _10180_, _04458_);
  and (_10182_, _10180_, _04458_);
  nor (_10183_, _10182_, _10181_);
  nor (_10184_, _05405_, \oc8051_golden_model_1.PC [10]);
  nor (_10185_, _10184_, _05398_);
  not (_10186_, _10185_);
  nor (_10187_, _10186_, _04458_);
  and (_10188_, _10186_, _04458_);
  nor (_10189_, _10188_, _10187_);
  and (_10190_, _10189_, _10183_);
  nor (_10191_, _05404_, \oc8051_golden_model_1.PC [9]);
  nor (_10192_, _10191_, _05405_);
  not (_10193_, _10192_);
  nor (_10194_, _10193_, _04458_);
  and (_10195_, _10193_, _04458_);
  nor (_10196_, _10195_, _10194_);
  nor (_10197_, _05323_, _04458_);
  and (_10198_, _05323_, _04458_);
  and (_10199_, _05317_, _04538_);
  nor (_10200_, _10199_, \oc8051_golden_model_1.PC [6]);
  nor (_10201_, _10200_, _05318_);
  not (_10202_, _10201_);
  nor (_10203_, _10202_, _04752_);
  and (_10204_, _10202_, _04752_);
  nor (_10205_, _10204_, _10203_);
  not (_10206_, _10205_);
  and (_10207_, _05317_, \oc8051_golden_model_1.PC [4]);
  nor (_10208_, _10207_, \oc8051_golden_model_1.PC [5]);
  nor (_10209_, _10208_, _10199_);
  not (_10210_, _10209_);
  nor (_10211_, _10210_, _04815_);
  and (_10212_, _10210_, _04815_);
  nor (_10213_, _05317_, \oc8051_golden_model_1.PC [4]);
  nor (_10214_, _10213_, _10207_);
  not (_10215_, _10214_);
  nor (_10216_, _10215_, _04784_);
  nor (_10217_, _05316_, \oc8051_golden_model_1.PC [3]);
  nor (_10218_, _10217_, _05317_);
  not (_10219_, _10218_);
  nor (_10220_, _10219_, _02324_);
  and (_10221_, _10219_, _02324_);
  nor (_10222_, _01443_, \oc8051_golden_model_1.PC [2]);
  nor (_10223_, _10222_, _05316_);
  not (_10224_, _10223_);
  nor (_10225_, _10224_, _02494_);
  not (_10226_, _01805_);
  nor (_10227_, _02893_, _10226_);
  nor (_10228_, _02679_, \oc8051_golden_model_1.PC [0]);
  and (_10229_, _02893_, _10226_);
  nor (_10230_, _10229_, _10227_);
  and (_10231_, _10230_, _10228_);
  nor (_10232_, _10231_, _10227_);
  and (_10233_, _10224_, _02494_);
  nor (_10234_, _10233_, _10225_);
  not (_10235_, _10234_);
  nor (_10236_, _10235_, _10232_);
  nor (_10237_, _10236_, _10225_);
  nor (_10238_, _10237_, _10221_);
  nor (_10239_, _10238_, _10220_);
  and (_10240_, _10215_, _04784_);
  nor (_10241_, _10240_, _10216_);
  not (_10242_, _10241_);
  nor (_10243_, _10242_, _10239_);
  nor (_10244_, _10243_, _10216_);
  nor (_10245_, _10244_, _10212_);
  nor (_10246_, _10245_, _10211_);
  nor (_10247_, _10246_, _10206_);
  nor (_10248_, _10247_, _10203_);
  nor (_10249_, _10248_, _10198_);
  or (_10250_, _10249_, _10197_);
  nor (_10251_, _05321_, \oc8051_golden_model_1.PC [8]);
  nor (_10252_, _10251_, _05404_);
  not (_10253_, _10252_);
  nor (_10254_, _10253_, _04458_);
  and (_10255_, _10253_, _04458_);
  nor (_10256_, _10255_, _10254_);
  and (_10257_, _10256_, _10250_);
  and (_10258_, _10257_, _10196_);
  and (_10259_, _10258_, _10190_);
  nor (_10260_, _10254_, _10194_);
  not (_10261_, _10260_);
  and (_10262_, _10261_, _10190_);
  or (_10263_, _10262_, _10187_);
  or (_10264_, _10263_, _10259_);
  nor (_10265_, _10264_, _10181_);
  and (_10266_, _10174_, _04458_);
  nor (_10267_, _10266_, _10175_);
  not (_10268_, _10267_);
  nor (_10269_, _10268_, _10265_);
  nor (_10270_, _10269_, _10175_);
  nor (_10271_, _10270_, _10171_);
  nor (_10272_, _10271_, _10170_);
  nor (_10273_, _10272_, _10167_);
  nor (_10274_, _10273_, _10164_);
  not (_10275_, _05412_);
  and (_10276_, _10275_, _04458_);
  nor (_10277_, _10275_, _04458_);
  nor (_10278_, _10277_, _10276_);
  and (_10279_, _10278_, _10274_);
  nor (_10280_, _10278_, _10274_);
  or (_10281_, _10280_, _10279_);
  or (_10282_, _10281_, _08922_);
  nand (_10283_, _08922_, _10275_);
  and (_10284_, _10283_, _02246_);
  and (_10285_, _10284_, _10282_);
  and (_10286_, _05428_, _02153_);
  nor (_10287_, _08707_, _06823_);
  not (_10288_, _10287_);
  and (_10289_, _04257_, _04208_);
  and (_10290_, _04644_, _10289_);
  and (_10291_, _04010_, _03902_);
  and (_10292_, _10291_, _04641_);
  and (_10293_, _10292_, _10290_);
  or (_10294_, _10293_, _10281_);
  nand (_10295_, _10292_, _10290_);
  or (_10296_, _10295_, _05412_);
  and (_10297_, _10296_, _10294_);
  or (_10298_, _10297_, _03006_);
  not (_10299_, _06845_);
  nor (_10300_, _02030_, _01693_);
  nor (_10301_, _10300_, _01746_);
  not (_10302_, _10301_);
  and (_10303_, _10302_, \oc8051_golden_model_1.PC [15]);
  nor (_10304_, _10303_, _02062_);
  nor (_10305_, _10304_, _06855_);
  or (_10306_, _10305_, _02060_);
  and (_10307_, _10306_, _06859_);
  or (_10308_, _10307_, _02160_);
  and (_10309_, _10308_, _10299_);
  or (_10310_, _10309_, _10117_);
  and (_10311_, _06859_, _01747_);
  nor (_10312_, _10301_, _06855_);
  nand (_10313_, _10312_, _06847_);
  nor (_10314_, _10313_, _10305_);
  nand (_10315_, _10314_, _10311_);
  not (_10316_, _05428_);
  nand (_10317_, _09495_, _06847_);
  nand (_10318_, _10317_, _10316_);
  and (_10319_, _10318_, _10315_);
  or (_10320_, _10319_, _06845_);
  and (_10321_, _10320_, _01752_);
  and (_10322_, _10321_, _10310_);
  not (_10323_, _01752_);
  nand (_10324_, _05428_, _10323_);
  nand (_10325_, _10324_, _04534_);
  or (_10326_, _10325_, _10322_);
  nor (_10327_, _05417_, \oc8051_golden_model_1.PC [14]);
  nor (_10328_, _10327_, _05418_);
  and (_10329_, _10328_, _01952_);
  nor (_10330_, _10328_, _01952_);
  nor (_10331_, _10330_, _10329_);
  not (_10332_, _10331_);
  nor (_10333_, _05416_, \oc8051_golden_model_1.PC [13]);
  nor (_10334_, _10333_, _05417_);
  and (_10335_, _10334_, _01952_);
  nor (_10336_, _10334_, _01952_);
  nor (_10337_, _05415_, \oc8051_golden_model_1.PC [12]);
  nor (_10338_, _10337_, _05416_);
  and (_10339_, _10338_, _01952_);
  nor (_10340_, _05422_, \oc8051_golden_model_1.PC [11]);
  nor (_10341_, _10340_, _05423_);
  and (_10342_, _10341_, _01952_);
  nor (_10343_, _10341_, _01952_);
  nor (_10344_, _10343_, _10342_);
  nor (_10345_, _05421_, \oc8051_golden_model_1.PC [10]);
  nor (_10346_, _10345_, _05414_);
  and (_10347_, _10346_, _01952_);
  nor (_10348_, _10346_, _01952_);
  nor (_10349_, _10348_, _10347_);
  and (_10350_, _10349_, _10344_);
  nor (_10351_, _05420_, \oc8051_golden_model_1.PC [9]);
  nor (_10352_, _10351_, _05421_);
  and (_10353_, _10352_, _01952_);
  nor (_10354_, _10352_, _01952_);
  nor (_10355_, _10354_, _10353_);
  and (_10356_, _04543_, _01952_);
  nor (_10357_, _04543_, _01952_);
  and (_10358_, _04538_, _01824_);
  nor (_10359_, _10358_, \oc8051_golden_model_1.PC [6]);
  nor (_10360_, _10359_, _04540_);
  not (_10361_, _10360_);
  nor (_10362_, _10361_, _02118_);
  and (_10363_, _10361_, _02118_);
  nor (_10364_, _10363_, _10362_);
  not (_10365_, _10364_);
  and (_10366_, _01824_, \oc8051_golden_model_1.PC [4]);
  nor (_10367_, _10366_, \oc8051_golden_model_1.PC [5]);
  nor (_10368_, _10367_, _10358_);
  not (_10369_, _10368_);
  nor (_10370_, _10369_, _02410_);
  and (_10371_, _10369_, _02410_);
  nor (_10372_, _01824_, \oc8051_golden_model_1.PC [4]);
  nor (_10373_, _10372_, _10366_);
  not (_10374_, _10373_);
  nor (_10375_, _10374_, _02825_);
  nor (_10376_, _01983_, _02264_);
  and (_10377_, _01983_, _02264_);
  nor (_10378_, _02452_, _01702_);
  nor (_10379_, _02859_, \oc8051_golden_model_1.PC [1]);
  nor (_10380_, _02027_, _01439_);
  and (_10381_, _02859_, \oc8051_golden_model_1.PC [1]);
  nor (_10382_, _10381_, _10379_);
  and (_10383_, _10382_, _10380_);
  nor (_10384_, _10383_, _10379_);
  and (_10385_, _02452_, _01702_);
  nor (_10386_, _10385_, _10378_);
  not (_10387_, _10386_);
  nor (_10388_, _10387_, _10384_);
  nor (_10389_, _10388_, _10378_);
  nor (_10390_, _10389_, _10377_);
  nor (_10391_, _10390_, _10376_);
  and (_10392_, _10374_, _02825_);
  nor (_10393_, _10392_, _10375_);
  not (_10394_, _10393_);
  nor (_10395_, _10394_, _10391_);
  nor (_10396_, _10395_, _10375_);
  nor (_10397_, _10396_, _10371_);
  nor (_10398_, _10397_, _10370_);
  nor (_10399_, _10398_, _10365_);
  nor (_10400_, _10399_, _10362_);
  nor (_10401_, _10400_, _10357_);
  or (_10402_, _10401_, _10356_);
  nor (_10403_, _04542_, \oc8051_golden_model_1.PC [8]);
  nor (_10404_, _10403_, _05420_);
  and (_10405_, _10404_, _01952_);
  nor (_10406_, _10404_, _01952_);
  nor (_10407_, _10406_, _10405_);
  and (_10408_, _10407_, _10402_);
  and (_10409_, _10408_, _10355_);
  and (_10410_, _10409_, _10350_);
  nor (_10411_, _10405_, _10353_);
  not (_10412_, _10411_);
  and (_10413_, _10412_, _10350_);
  or (_10414_, _10413_, _10347_);
  or (_10415_, _10414_, _10410_);
  nor (_10416_, _10415_, _10342_);
  nor (_10417_, _10338_, _01952_);
  nor (_10418_, _10417_, _10339_);
  not (_10419_, _10418_);
  nor (_10420_, _10419_, _10416_);
  nor (_10421_, _10420_, _10339_);
  nor (_10422_, _10421_, _10336_);
  nor (_10423_, _10422_, _10335_);
  nor (_10424_, _10423_, _10332_);
  nor (_10425_, _10424_, _10329_);
  nor (_10426_, _05428_, _01952_);
  and (_10427_, _05428_, _01952_);
  nor (_10428_, _10427_, _10426_);
  and (_10429_, _10428_, _10425_);
  nor (_10430_, _10428_, _10425_);
  or (_10431_, _10430_, _10429_);
  and (_10432_, _04526_, _04524_);
  and (_10433_, _03161_, _03002_);
  and (_10434_, _05349_, _10433_);
  and (_10435_, _10434_, _10432_);
  or (_10436_, _10435_, _10431_);
  nand (_10437_, _10434_, _10432_);
  or (_10438_, _10437_, _05428_);
  and (_10439_, _10438_, _10436_);
  or (_10440_, _10439_, _04534_);
  nand (_10441_, _10440_, _10326_);
  nor (_10442_, _02158_, _02079_);
  nand (_10443_, _10442_, _10441_);
  and (_10444_, _10443_, _10298_);
  or (_10445_, _10444_, _10288_);
  nor (_10446_, _02155_, _03446_);
  and (_10447_, _10446_, _02058_);
  and (_10448_, _10287_, _04550_);
  or (_10449_, _10448_, _10117_);
  and (_10450_, _10449_, _10447_);
  and (_10451_, _10450_, _10445_);
  and (_10452_, _06820_, _06884_);
  or (_10453_, _10447_, _10316_);
  nand (_10454_, _10453_, _10452_);
  or (_10455_, _10454_, _10451_);
  or (_10456_, _10452_, _10117_);
  and (_10457_, _10456_, _02549_);
  and (_10458_, _10457_, _10455_);
  or (_10459_, _10458_, _10286_);
  nor (_10460_, _08728_, _06888_);
  and (_10461_, _10460_, _10459_);
  not (_10462_, _10460_);
  nand (_10463_, _10462_, _10117_);
  not (_10464_, _01757_);
  nor (_10465_, _02052_, _10464_);
  and (_10466_, _10465_, _02054_);
  nand (_10467_, _10466_, _10463_);
  or (_10468_, _10467_, _10461_);
  or (_10469_, _10466_, _05428_);
  nor (_10470_, _05442_, _01749_);
  nor (_10471_, _10470_, _02230_);
  and (_10472_, _10471_, _10469_);
  and (_10473_, _10472_, _10468_);
  nand (_10474_, _08770_, _10275_);
  not (_10475_, _10471_);
  or (_10476_, _10281_, _08770_);
  and (_10477_, _10476_, _10475_);
  and (_10478_, _10477_, _10474_);
  or (_10479_, _10478_, _08790_);
  or (_10480_, _10479_, _10473_);
  and (_10481_, _08842_, _05412_);
  nand (_10482_, _08841_, _08826_);
  and (_10483_, _10281_, _10482_);
  or (_10484_, _10483_, _10481_);
  or (_10485_, _10484_, _08836_);
  and (_10486_, _10485_, _10480_);
  or (_10487_, _10486_, _02171_);
  and (_10488_, _08877_, _05412_);
  not (_10489_, _08877_);
  and (_10490_, _10281_, _10489_);
  or (_10491_, _10490_, _02547_);
  or (_10492_, _10491_, _10488_);
  and (_10493_, _10492_, _08917_);
  and (_10494_, _10493_, _10487_);
  or (_10495_, _10494_, _10285_);
  and (_10496_, _10495_, _08882_);
  nand (_10497_, _10117_, _08881_);
  nor (_10498_, _04916_, _01754_);
  or (_10499_, _10498_, _02046_);
  nor (_10500_, _10499_, _02131_);
  nor (_10501_, _02147_, _03310_);
  and (_10502_, _02133_, _02128_);
  nor (_10503_, _02614_, _10502_);
  and (_10504_, _10503_, _10501_);
  and (_10505_, _10504_, _02143_);
  and (_10506_, _10505_, _10500_);
  nand (_10507_, _10506_, _10497_);
  or (_10508_, _10507_, _10496_);
  or (_10509_, _10506_, _05428_);
  and (_10510_, _10509_, _10158_);
  and (_10511_, _10510_, _10508_);
  or (_10512_, _10511_, _10160_);
  not (_10513_, _01755_);
  nor (_10514_, _02181_, _10513_);
  and (_10515_, _10514_, _08505_);
  and (_10516_, _10515_, _10512_);
  not (_10517_, _10153_);
  nor (_10518_, _10515_, _10316_);
  or (_10519_, _10518_, _10517_);
  or (_10520_, _10519_, _10516_);
  and (_10521_, _10520_, _10154_);
  or (_10522_, _10521_, _07017_);
  or (_10523_, _07016_, _05428_);
  and (_10524_, _10523_, _01778_);
  and (_10525_, _10524_, _10522_);
  and (_10526_, _10117_, _01876_);
  nor (_10527_, _02042_, _01767_);
  not (_10528_, _10527_);
  or (_10529_, _10528_, _10526_);
  or (_10530_, _10529_, _10525_);
  or (_10531_, _10527_, _05428_);
  and (_10532_, _10531_, _07633_);
  and (_10533_, _10532_, _10530_);
  and (_10534_, _05444_, _02032_);
  nand (_10535_, _05412_, _02218_);
  nand (_10536_, _10535_, _10534_);
  or (_10537_, _10536_, _10533_);
  or (_10538_, _10534_, _05428_);
  and (_10539_, _10538_, _02037_);
  and (_10540_, _10539_, _10537_);
  or (_10541_, _10540_, _10152_);
  nor (_10542_, _06202_, _01775_);
  and (_10543_, _10542_, _10541_);
  nor (_10544_, _02124_, _01711_);
  not (_10545_, _10544_);
  not (_10546_, _10542_);
  and (_10547_, _10546_, _10117_);
  or (_10548_, _10547_, _10545_);
  or (_10549_, _10548_, _10543_);
  and (_10550_, _01710_, _01696_);
  not (_10551_, _10550_);
  or (_10552_, _10544_, _05428_);
  and (_10553_, _10552_, _10551_);
  and (_10554_, _10553_, _10549_);
  and (_10555_, _10550_, _10431_);
  or (_10556_, _10555_, _04920_);
  or (_10557_, _10556_, _10554_);
  and (_10558_, _10557_, _10151_);
  or (_10559_, _10558_, _01994_);
  or (_10560_, _05412_, _01995_);
  and (_10561_, _10560_, _07240_);
  and (_10562_, _10561_, _10559_);
  and (_10563_, _07239_, _05428_);
  or (_10564_, _10563_, _10562_);
  and (_10565_, _10564_, _10150_);
  and (_10566_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_10567_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_10568_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_10569_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_10570_, _10569_, _10568_);
  not (_10571_, _10570_);
  and (_10572_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_10573_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_10574_, _10573_, _10572_);
  not (_10575_, _10574_);
  and (_10576_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10577_, _01843_, _01839_);
  nor (_10578_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_10579_, _10578_, _10576_);
  not (_10580_, _10579_);
  nor (_10581_, _10580_, _10577_);
  nor (_10582_, _10581_, _10576_);
  nor (_10583_, _10582_, _10575_);
  nor (_10584_, _10583_, _10572_);
  nor (_10585_, _10584_, _10571_);
  nor (_10586_, _10585_, _10568_);
  nor (_10587_, _10586_, _10567_);
  or (_10588_, _10587_, _10566_);
  and (_10589_, _10588_, \oc8051_golden_model_1.DPH [0]);
  and (_10590_, _10589_, \oc8051_golden_model_1.DPH [1]);
  and (_10591_, _10590_, \oc8051_golden_model_1.DPH [2]);
  and (_10592_, _10591_, \oc8051_golden_model_1.DPH [3]);
  and (_10593_, _10592_, \oc8051_golden_model_1.DPH [4]);
  and (_10594_, _10593_, \oc8051_golden_model_1.DPH [5]);
  and (_10595_, _10594_, \oc8051_golden_model_1.DPH [6]);
  nand (_10596_, _10595_, \oc8051_golden_model_1.DPH [7]);
  or (_10597_, _10595_, \oc8051_golden_model_1.DPH [7]);
  and (_10598_, _10597_, _10149_);
  and (_10599_, _10598_, _10596_);
  nor (_10600_, _02123_, _01718_);
  not (_10601_, _10600_);
  or (_10602_, _10601_, _10599_);
  or (_10603_, _10602_, _10565_);
  and (_10604_, _01717_, _01696_);
  not (_10605_, _10604_);
  or (_10606_, _10600_, _05428_);
  and (_10607_, _10606_, _10605_);
  and (_10608_, _10607_, _10603_);
  not (_10609_, _10147_);
  or (_10610_, _10431_, _07587_);
  not (_10611_, _07587_);
  or (_10612_, _10611_, _05428_);
  and (_10613_, _10612_, _10604_);
  and (_10614_, _10613_, _10610_);
  or (_10615_, _10614_, _10609_);
  or (_10616_, _10615_, _10608_);
  and (_10617_, _10616_, _10148_);
  nor (_10618_, _06734_, _02329_);
  not (_10619_, _10618_);
  or (_10620_, _10619_, _10617_);
  or (_10621_, _10618_, _05428_);
  and (_10622_, _10621_, _03059_);
  and (_10623_, _10622_, _10620_);
  and (_10624_, _05412_, _02210_);
  nor (_10625_, _02331_, _01722_);
  not (_10626_, _10625_);
  or (_10627_, _10626_, _10624_);
  or (_10628_, _10627_, _10623_);
  and (_10629_, _01721_, _01696_);
  not (_10630_, _10629_);
  or (_10631_, _10625_, _05428_);
  and (_10632_, _10631_, _10630_);
  and (_10633_, _10632_, _10628_);
  not (_10634_, _10139_);
  or (_10635_, _10431_, _10611_);
  or (_10636_, _07587_, _05428_);
  and (_10637_, _10636_, _10629_);
  and (_10638_, _10637_, _10635_);
  or (_10639_, _10638_, _10634_);
  or (_10640_, _10639_, _10633_);
  and (_10641_, _10640_, _10140_);
  or (_10642_, _10641_, _10136_);
  or (_10643_, _10135_, _05428_);
  and (_10644_, _10643_, _02208_);
  and (_10645_, _10644_, _10642_);
  and (_10646_, _05412_, _02206_);
  or (_10647_, _10646_, _09562_);
  or (_10648_, _10647_, _10645_);
  and (_10649_, _01727_, _01696_);
  not (_10650_, _10649_);
  or (_10651_, _09561_, _05428_);
  and (_10652_, _10651_, _10650_);
  and (_10653_, _10652_, _10648_);
  not (_10654_, _10133_);
  or (_10655_, _10431_, \oc8051_golden_model_1.PSW [7]);
  or (_10656_, _05428_, _06707_);
  and (_10657_, _10656_, _10649_);
  and (_10658_, _10657_, _10655_);
  or (_10659_, _10658_, _10654_);
  or (_10660_, _10659_, _10653_);
  and (_10661_, _10660_, _10134_);
  or (_10662_, _10661_, _07340_);
  or (_10663_, _07339_, _05428_);
  and (_10664_, _10663_, _04953_);
  and (_10665_, _10664_, _10662_);
  not (_10666_, _10124_);
  and (_10667_, _05412_, _02202_);
  or (_10668_, _10667_, _10666_);
  or (_10669_, _10668_, _10665_);
  and (_10670_, _10669_, _10126_);
  not (_10671_, _10120_);
  or (_10672_, _10431_, _06707_);
  or (_10673_, _05428_, \oc8051_golden_model_1.PSW [7]);
  and (_10674_, _10673_, _10122_);
  and (_10675_, _10674_, _10672_);
  or (_10676_, _10675_, _10671_);
  or (_10677_, _10676_, _10670_);
  and (_10678_, _10677_, _10121_);
  or (_10679_, _10678_, _07386_);
  or (_10680_, _07385_, _05428_);
  and (_10681_, _10680_, _07416_);
  and (_10682_, _10681_, _10679_);
  and (_10683_, _10117_, _07415_);
  or (_10684_, _10683_, _02350_);
  or (_10685_, _10684_, _10682_);
  nand (_10686_, _03796_, _02350_);
  and (_10687_, _10686_, _10685_);
  or (_10688_, _10687_, _01726_);
  not (_10689_, _02200_);
  or (_10690_, _05428_, _04964_);
  and (_10691_, _10690_, _10689_);
  and (_10692_, _10691_, _10688_);
  not (_10693_, _10118_);
  not (_10694_, _08690_);
  or (_10695_, _10281_, _10694_);
  or (_10696_, _08690_, _05412_);
  and (_10697_, _10696_, _02200_);
  and (_10698_, _10697_, _10695_);
  or (_10699_, _10698_, _10693_);
  or (_10700_, _10699_, _10692_);
  and (_10701_, _10700_, _10119_);
  or (_10702_, _10701_, _07489_);
  or (_10703_, _07488_, _05428_);
  and (_10704_, _10703_, _07534_);
  and (_10705_, _10704_, _10702_);
  and (_10706_, _10117_, _07533_);
  or (_10707_, _10706_, _02083_);
  or (_10708_, _10707_, _10705_);
  nand (_10709_, _03796_, _02083_);
  and (_10710_, _10709_, _10708_);
  or (_10711_, _10710_, _01738_);
  not (_10712_, _01738_);
  or (_10713_, _05428_, _10712_);
  and (_10714_, _10713_, _02367_);
  and (_10715_, _10714_, _10711_);
  or (_10716_, _10281_, _08690_);
  nand (_10717_, _08690_, _10275_);
  and (_10718_, _10717_, _10716_);
  and (_10719_, _10718_, _02243_);
  nor (_10720_, _05442_, _04969_);
  nor (_10721_, _10720_, _03273_);
  and (_10722_, _10721_, _04984_);
  not (_10723_, _10722_);
  or (_10724_, _10723_, _10719_);
  or (_10725_, _10724_, _10715_);
  or (_10726_, _10722_, _10117_);
  and (_10727_, _10726_, _02778_);
  and (_10728_, _10727_, _10725_);
  nand (_10729_, _05428_, _02366_);
  nand (_10730_, _10729_, _07581_);
  or (_10731_, _10730_, _10728_);
  or (_10732_, _10117_, _07581_);
  and (_10733_, _10732_, _05395_);
  and (_10734_, _10733_, _10731_);
  and (_10735_, _01989_, _01952_);
  or (_10736_, _10735_, _01733_);
  or (_10737_, _10736_, _10734_);
  not (_10738_, _01733_);
  or (_10739_, _05428_, _10738_);
  and (_10740_, _10739_, _01698_);
  and (_10741_, _10740_, _10737_);
  and (_10742_, _10718_, _01697_);
  not (_10743_, _01731_);
  nor (_10744_, _10300_, _10743_);
  or (_10745_, _10744_, _10742_);
  or (_10746_, _10745_, _10741_);
  not (_10747_, _10744_);
  or (_10748_, _10747_, _10117_);
  and (_10749_, _10748_, _02082_);
  and (_10750_, _10749_, _10746_);
  nor (_10751_, _07606_, _07599_);
  nand (_10752_, _05428_, _02081_);
  nand (_10753_, _10752_, _10751_);
  or (_10754_, _10753_, _10750_);
  not (_10755_, _02198_);
  or (_10756_, _10117_, _10751_);
  and (_10757_, _10756_, _10755_);
  and (_10758_, _10757_, _10754_);
  and (_10759_, _02198_, _01952_);
  or (_10760_, _10759_, _01732_);
  or (_10761_, _10760_, _10758_);
  and (_10762_, _01731_, _01696_);
  not (_10763_, _10762_);
  not (_10764_, _01732_);
  or (_10765_, _05428_, _10764_);
  and (_10766_, _10765_, _10763_);
  and (_10767_, _10766_, _10761_);
  and (_10768_, _10762_, _10117_);
  or (_10769_, _10768_, _10767_);
  or (_10770_, _10769_, _39633_);
  or (_10771_, _39632_, \oc8051_golden_model_1.PC [15]);
  and (_10772_, _10771_, _39026_);
  and (_38606_, _10772_, _10770_);
  and (_10773_, _39633_, \oc8051_golden_model_1.P0INREG [7]);
  or (_10774_, _10773_, _40036_);
  and (_38607_, _10774_, _39026_);
  and (_10775_, _39633_, \oc8051_golden_model_1.P1INREG [7]);
  or (_10776_, _10775_, _39694_);
  and (_38609_, _10776_, _39026_);
  and (_10777_, _39633_, \oc8051_golden_model_1.P2INREG [7]);
  or (_10778_, _10777_, _39818_);
  and (_38610_, _10778_, _39026_);
  and (_10779_, _39633_, \oc8051_golden_model_1.P3INREG [7]);
  or (_10780_, _10779_, _39750_);
  and (_38611_, _10780_, _39026_);
  and (_10781_, _03384_, _03101_);
  nor (_10782_, _10781_, _03386_);
  nor (_10783_, _03555_, _03385_);
  nor (_10784_, _10783_, _03743_);
  and (_10785_, _10784_, _10782_);
  and (_10786_, _10785_, _03384_);
  not (_10787_, _10786_);
  nand (_10788_, _01733_, _01439_);
  nor (_10789_, _04257_, \oc8051_golden_model_1.ACC [0]);
  nand (_10790_, _10789_, _04959_);
  and (_10791_, _04257_, \oc8051_golden_model_1.ACC [0]);
  nor (_10792_, _10791_, _10789_);
  and (_10793_, _10792_, _03062_);
  not (_10794_, _02035_);
  or (_10795_, _10794_, _03002_);
  nor (_10796_, _08608_, _03808_);
  and (_10797_, _03808_, \oc8051_golden_model_1.PSW [7]);
  nor (_10798_, _10797_, _10796_);
  nor (_10799_, _10798_, _04461_);
  nand (_10800_, _05120_, _03835_);
  nand (_10801_, _10800_, _07093_);
  and (_10802_, _10801_, _03041_);
  and (_10803_, _03015_, _03002_);
  nor (_10804_, _01747_, _01439_);
  and (_10805_, _01747_, \oc8051_golden_model_1.ACC [0]);
  or (_10806_, _10805_, _10804_);
  and (_10807_, _10806_, _04534_);
  and (_10808_, _04535_, _03020_);
  or (_10809_, _10808_, _10807_);
  and (_10810_, _10809_, _03165_);
  nor (_10811_, _04257_, _03165_);
  or (_10812_, _10811_, _10810_);
  and (_10813_, _10812_, _04519_);
  nand (_10814_, _08986_, _08585_);
  and (_10815_, _10814_, _03005_);
  or (_10816_, _10815_, _03446_);
  or (_10817_, _10816_, _10813_);
  nor (_10818_, _01745_, \oc8051_golden_model_1.PC [0]);
  nor (_10819_, _10818_, _03015_);
  and (_10820_, _10819_, _10817_);
  or (_10821_, _10820_, _10803_);
  and (_10822_, _10821_, _04505_);
  nor (_10823_, _08986_, _03808_);
  and (_10824_, _10823_, _03024_);
  or (_10825_, _10824_, _02052_);
  or (_10826_, _10825_, _10822_);
  nand (_10827_, _07094_, _02052_);
  and (_10828_, _10827_, _02050_);
  and (_10829_, _10828_, _10826_);
  nor (_10830_, _08987_, _02050_);
  and (_10831_, _10830_, _10814_);
  or (_10832_, _10831_, _10829_);
  and (_10833_, _10832_, _01750_);
  or (_10834_, _01750_, _01439_);
  nand (_10835_, _02144_, _10834_);
  or (_10836_, _10835_, _10833_);
  nand (_10837_, _07094_, _02145_);
  and (_10838_, _10837_, _04559_);
  and (_10839_, _10838_, _10836_);
  or (_10840_, _10839_, _10802_);
  and (_10841_, _10840_, _04461_);
  or (_10842_, _10841_, _10799_);
  and (_10843_, _10842_, _04460_);
  and (_10844_, _01767_, \oc8051_golden_model_1.PC [0]);
  or (_10845_, _02035_, _10844_);
  or (_10846_, _10845_, _10843_);
  and (_10847_, _10846_, _10795_);
  or (_10848_, _10847_, _02033_);
  or (_10849_, _05120_, _04712_);
  and (_10850_, _10849_, _02039_);
  and (_10851_, _10850_, _10848_);
  and (_10852_, _04458_, _03002_);
  and (_10853_, _04818_, \oc8051_golden_model_1.IP [0]);
  and (_10854_, _04833_, \oc8051_golden_model_1.PSW [0]);
  nor (_10855_, _10854_, _10853_);
  and (_10856_, _04829_, \oc8051_golden_model_1.ACC [0]);
  and (_10857_, _04824_, \oc8051_golden_model_1.B [0]);
  nor (_10858_, _10857_, _10856_);
  and (_10859_, _10858_, _10855_);
  and (_10860_, _04843_, \oc8051_golden_model_1.TH1 [0]);
  not (_10861_, _10860_);
  and (_10862_, _04849_, \oc8051_golden_model_1.TL0 [0]);
  and (_10863_, _04852_, \oc8051_golden_model_1.SP [0]);
  nor (_10864_, _10863_, _10862_);
  and (_10865_, _10864_, _10861_);
  and (_10866_, _10865_, _10859_);
  and (_10867_, _04864_, \oc8051_golden_model_1.TCON [0]);
  and (_10868_, _04857_, \oc8051_golden_model_1.TH0 [0]);
  nor (_10869_, _10868_, _10867_);
  and (_10870_, _04868_, \oc8051_golden_model_1.PCON [0]);
  and (_10871_, _04861_, \oc8051_golden_model_1.TL1 [0]);
  nor (_10872_, _10871_, _10870_);
  and (_10873_, _10872_, _10869_);
  and (_10874_, _04872_, \oc8051_golden_model_1.DPL [0]);
  not (_10875_, _10874_);
  and (_10876_, _04875_, \oc8051_golden_model_1.P0INREG [0]);
  not (_10877_, _10876_);
  nand (_10878_, _04879_, \oc8051_golden_model_1.P3INREG [0]);
  and (_10879_, _04882_, \oc8051_golden_model_1.P1INREG [0]);
  and (_10880_, _04885_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_10881_, _10880_, _10879_);
  and (_10882_, _10881_, _10878_);
  and (_10883_, _10882_, _10877_);
  and (_10884_, _10883_, _10875_);
  and (_10885_, _04891_, \oc8051_golden_model_1.IE [0]);
  and (_10886_, _04894_, \oc8051_golden_model_1.SBUF [0]);
  and (_10887_, _04896_, \oc8051_golden_model_1.SCON [0]);
  or (_10888_, _10887_, _10886_);
  nor (_10889_, _10888_, _10885_);
  and (_10890_, _04900_, \oc8051_golden_model_1.TMOD [0]);
  and (_10891_, _04902_, \oc8051_golden_model_1.DPH [0]);
  nor (_10892_, _10891_, _10890_);
  and (_10893_, _10892_, _10889_);
  and (_10894_, _10893_, _10884_);
  and (_10895_, _10894_, _10873_);
  and (_10896_, _10895_, _10866_);
  not (_10897_, _10896_);
  nor (_10898_, _10897_, _10852_);
  nor (_10899_, _10898_, _02039_);
  or (_10900_, _10899_, _04920_);
  or (_10901_, _10900_, _10851_);
  and (_10902_, _04920_, _02027_);
  nor (_10903_, _10902_, _01996_);
  and (_10904_, _10903_, _10901_);
  and (_10905_, _04837_, _01996_);
  or (_10906_, _10905_, _01718_);
  or (_10907_, _10906_, _10904_);
  nand (_10908_, _01718_, _01439_);
  and (_10909_, _10908_, _10907_);
  or (_10910_, _10909_, _03060_);
  not (_10911_, _03060_);
  and (_10912_, _04257_, _04837_);
  nor (_10913_, _04257_, _04837_);
  nor (_10914_, _10913_, _10912_);
  or (_10915_, _10914_, _10911_);
  and (_10916_, _10915_, _04938_);
  and (_10917_, _10916_, _10910_);
  or (_10918_, _10917_, _10793_);
  and (_10919_, _10918_, _04937_);
  and (_10920_, _10912_, _03064_);
  or (_10921_, _10920_, _03066_);
  or (_10922_, _10921_, _10919_);
  or (_10923_, _10791_, _04949_);
  and (_10924_, _10923_, _10922_);
  or (_10925_, _10924_, _01728_);
  and (_10926_, _01728_, _01439_);
  nor (_10927_, _10926_, _04954_);
  and (_10928_, _10927_, _10925_);
  nor (_10929_, _10913_, _04960_);
  or (_10930_, _10929_, _04959_);
  or (_10931_, _10930_, _10928_);
  and (_10932_, _10931_, _10790_);
  or (_10933_, _10932_, _01726_);
  nand (_10934_, _01726_, _01439_);
  and (_10935_, _10934_, _10721_);
  and (_10936_, _10935_, _10933_);
  nor (_10937_, _10721_, _03002_);
  or (_10938_, _10937_, _10936_);
  and (_10939_, _10938_, _04984_);
  nor (_10940_, _05120_, _04984_);
  or (_10941_, _10940_, _03083_);
  or (_10942_, _10941_, _10939_);
  nand (_10943_, _04257_, _03083_);
  and (_10944_, _10943_, _05395_);
  and (_10945_, _10944_, _10942_);
  and (_10946_, _01989_, _01439_);
  or (_10947_, _10946_, _01733_);
  or (_10948_, _10947_, _10945_);
  and (_10949_, _10948_, _10788_);
  or (_10950_, _10949_, _01992_);
  nand (_10951_, _01731_, _01693_);
  or (_10952_, _10796_, _03377_);
  and (_10953_, _10952_, _10951_);
  and (_10954_, _10953_, _10950_);
  nor (_10955_, _10951_, _03002_);
  or (_10956_, _10955_, _02785_);
  or (_10957_, _10956_, _10954_);
  nand (_10958_, _05120_, _02785_);
  and (_10959_, _10958_, _10957_);
  or (_10960_, _10959_, _03098_);
  nand (_10961_, _04257_, _03098_);
  and (_10962_, _10961_, _03384_);
  and (_10963_, _10962_, _10960_);
  or (_10964_, _10963_, _10787_);
  or (_10965_, _10786_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_10966_, _05390_, _05386_);
  nor (_10967_, _10966_, _05391_);
  and (_10968_, _10967_, _03106_);
  and (_10969_, _10968_, _05390_);
  not (_10970_, _10969_);
  and (_10971_, _10970_, _10965_);
  and (_10972_, _10971_, _10964_);
  and (_10973_, _05390_, _03106_);
  and (_10974_, _10973_, _10967_);
  nand (_10975_, _10253_, _01989_);
  or (_10976_, _10404_, _01989_);
  and (_10977_, _10976_, _10975_);
  and (_10978_, _10977_, _05390_);
  and (_10979_, _10978_, _10974_);
  or (_38643_, _10979_, _10972_);
  not (_10980_, _10951_);
  nor (_10981_, _05344_, _04525_);
  and (_10982_, _10981_, _10980_);
  nor (_10983_, _05364_, _05121_);
  nor (_10984_, _10983_, _04984_);
  not (_10985_, _03350_);
  and (_10986_, _01726_, _01412_);
  and (_10987_, _04208_, _02893_);
  nor (_10988_, _04208_, _02893_);
  nor (_10989_, _10988_, _10987_);
  and (_10990_, _10989_, _03060_);
  nand (_10991_, _03161_, _02035_);
  nor (_10992_, _08961_, _03803_);
  or (_10993_, _10992_, _04505_);
  nand (_10994_, _10981_, _04535_);
  and (_10995_, _01747_, \oc8051_golden_model_1.ACC [1]);
  or (_10996_, _01747_, \oc8051_golden_model_1.PC [1]);
  nand (_10997_, _04534_, _10996_);
  or (_10998_, _10997_, _10995_);
  and (_10999_, _10998_, _10994_);
  and (_11000_, _10999_, _03165_);
  nor (_11001_, _04643_, _04258_);
  nor (_11002_, _11001_, _03165_);
  or (_11003_, _11002_, _11000_);
  or (_11004_, _11003_, _03005_);
  nand (_11005_, _08961_, _08531_);
  or (_11006_, _11005_, _04519_);
  and (_11007_, _11006_, _11004_);
  or (_11008_, _11007_, _03446_);
  nor (_11009_, _01745_, _01412_);
  nor (_11010_, _11009_, _03015_);
  and (_11011_, _11010_, _11008_);
  and (_11012_, _03163_, _03015_);
  or (_11013_, _11012_, _03024_);
  or (_11014_, _11013_, _11011_);
  and (_11015_, _11014_, _10993_);
  or (_11016_, _11015_, _02052_);
  nand (_11017_, _07082_, _02052_);
  and (_11018_, _11017_, _02050_);
  and (_11019_, _11018_, _11016_);
  not (_11020_, _08962_);
  and (_11021_, _11005_, _11020_);
  and (_11022_, _11021_, _02049_);
  or (_11023_, _11022_, _11019_);
  and (_11024_, _11023_, _01750_);
  or (_11025_, _01750_, \oc8051_golden_model_1.PC [1]);
  nand (_11026_, _02144_, _11025_);
  or (_11027_, _11026_, _11024_);
  nand (_11028_, _07082_, _02145_);
  and (_11029_, _11028_, _04559_);
  and (_11030_, _11029_, _11027_);
  nand (_11031_, _05075_, _03835_);
  nand (_11032_, _11031_, _07081_);
  and (_11033_, _11032_, _03041_);
  or (_11034_, _11033_, _03040_);
  or (_11035_, _11034_, _11030_);
  nor (_11036_, _08553_, _03803_);
  and (_11037_, _03803_, \oc8051_golden_model_1.PSW [7]);
  nor (_11038_, _11037_, _11036_);
  nand (_11039_, _11038_, _03040_);
  and (_11040_, _11039_, _04460_);
  and (_11041_, _11040_, _11035_);
  and (_11042_, _01767_, _01412_);
  or (_11043_, _02035_, _11042_);
  or (_11044_, _11043_, _11041_);
  and (_11045_, _11044_, _10991_);
  or (_11046_, _11045_, _02033_);
  or (_11047_, _05075_, _04712_);
  and (_11048_, _11047_, _02039_);
  and (_11049_, _11048_, _11046_);
  nor (_11050_, _04716_, _03161_);
  and (_11051_, _04818_, \oc8051_golden_model_1.IP [1]);
  and (_11052_, _04824_, \oc8051_golden_model_1.B [1]);
  nor (_11053_, _11052_, _11051_);
  and (_11054_, _04829_, \oc8051_golden_model_1.ACC [1]);
  and (_11055_, _04833_, \oc8051_golden_model_1.PSW [1]);
  nor (_11056_, _11055_, _11054_);
  and (_11057_, _11056_, _11053_);
  and (_11058_, _04843_, \oc8051_golden_model_1.TH1 [1]);
  not (_11059_, _11058_);
  and (_11060_, _04849_, \oc8051_golden_model_1.TL0 [1]);
  and (_11061_, _04852_, \oc8051_golden_model_1.SP [1]);
  nor (_11062_, _11061_, _11060_);
  and (_11063_, _11062_, _11059_);
  and (_11064_, _11063_, _11057_);
  and (_11065_, _04864_, \oc8051_golden_model_1.TCON [1]);
  and (_11066_, _04857_, \oc8051_golden_model_1.TH0 [1]);
  nor (_11067_, _11066_, _11065_);
  and (_11068_, _04868_, \oc8051_golden_model_1.PCON [1]);
  and (_11069_, _04861_, \oc8051_golden_model_1.TL1 [1]);
  nor (_11070_, _11069_, _11068_);
  and (_11071_, _11070_, _11067_);
  and (_11072_, _04872_, \oc8051_golden_model_1.DPL [1]);
  not (_11073_, _11072_);
  and (_11074_, _04875_, \oc8051_golden_model_1.P0INREG [1]);
  not (_11075_, _11074_);
  nand (_11076_, _04879_, \oc8051_golden_model_1.P3INREG [1]);
  and (_11077_, _04882_, \oc8051_golden_model_1.P1INREG [1]);
  and (_11078_, _04885_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_11079_, _11078_, _11077_);
  and (_11080_, _11079_, _11076_);
  and (_11081_, _11080_, _11075_);
  and (_11082_, _11081_, _11073_);
  and (_11083_, _04891_, \oc8051_golden_model_1.IE [1]);
  and (_11084_, _04894_, \oc8051_golden_model_1.SBUF [1]);
  and (_11085_, _04896_, \oc8051_golden_model_1.SCON [1]);
  or (_11086_, _11085_, _11084_);
  nor (_11087_, _11086_, _11083_);
  and (_11088_, _04900_, \oc8051_golden_model_1.TMOD [1]);
  and (_11089_, _04902_, \oc8051_golden_model_1.DPH [1]);
  nor (_11090_, _11089_, _11088_);
  and (_11091_, _11090_, _11087_);
  and (_11092_, _11091_, _11082_);
  and (_11093_, _11092_, _11071_);
  and (_11094_, _11093_, _11064_);
  not (_11095_, _11094_);
  nor (_11096_, _11095_, _11050_);
  nor (_11097_, _11096_, _02039_);
  or (_11098_, _11097_, _04920_);
  or (_11099_, _11098_, _11049_);
  and (_11100_, _04920_, _02859_);
  nor (_11101_, _11100_, _01996_);
  and (_11102_, _11101_, _11099_);
  and (_11103_, _04846_, _01996_);
  or (_11104_, _11103_, _01718_);
  or (_11105_, _11104_, _11102_);
  and (_11106_, _01718_, \oc8051_golden_model_1.PC [1]);
  nor (_11107_, _11106_, _03060_);
  and (_11108_, _11107_, _11105_);
  or (_11109_, _11108_, _10990_);
  and (_11110_, _11109_, _04938_);
  nor (_11111_, _04208_, _01804_);
  and (_11112_, _04208_, _01804_);
  nor (_11113_, _11112_, _11111_);
  and (_11114_, _11113_, _03062_);
  or (_11115_, _11114_, _11110_);
  and (_11116_, _11115_, _04937_);
  and (_11117_, _10988_, _03064_);
  or (_11118_, _11117_, _11116_);
  and (_11119_, _11118_, _04949_);
  and (_11120_, _11111_, _03066_);
  or (_11121_, _11120_, _01728_);
  or (_11122_, _11121_, _11119_);
  and (_11123_, _01728_, \oc8051_golden_model_1.PC [1]);
  nor (_11124_, _11123_, _04954_);
  and (_11125_, _11124_, _11122_);
  nor (_11126_, _10987_, _04960_);
  or (_11127_, _11126_, _04959_);
  or (_11128_, _11127_, _11125_);
  nand (_11129_, _11112_, _04959_);
  and (_11130_, _11129_, _04964_);
  and (_11131_, _11130_, _11128_);
  or (_11132_, _11131_, _10986_);
  and (_11133_, _11132_, _10985_);
  nor (_11134_, _10981_, _10985_);
  or (_11135_, _11134_, _03276_);
  or (_11136_, _11135_, _11133_);
  nand (_11137_, _10981_, _03276_);
  and (_11138_, _11137_, _03723_);
  and (_11139_, _11138_, _11136_);
  nor (_11140_, _10981_, _03723_);
  or (_11141_, _11140_, _04979_);
  or (_11142_, _11141_, _11139_);
  nand (_11143_, _10981_, _04979_);
  and (_11144_, _11143_, _04984_);
  and (_11145_, _11144_, _11142_);
  or (_11146_, _11145_, _10984_);
  and (_11147_, _11146_, _04983_);
  nor (_11148_, _11001_, _04983_);
  or (_11149_, _11148_, _01989_);
  or (_11150_, _11149_, _11147_);
  nand (_11151_, _01989_, _10226_);
  and (_11152_, _11151_, _10738_);
  and (_11153_, _11152_, _11150_);
  and (_11154_, _01733_, _01412_);
  or (_11155_, _01992_, _11154_);
  or (_11156_, _11155_, _11153_);
  or (_11157_, _11036_, _03377_);
  and (_11158_, _11157_, _10951_);
  and (_11159_, _11158_, _11156_);
  or (_11160_, _11159_, _10982_);
  and (_11161_, _11160_, _05363_);
  and (_11162_, _10983_, _02785_);
  or (_11163_, _11162_, _03098_);
  or (_11164_, _11163_, _11161_);
  not (_11165_, _03098_);
  or (_11166_, _11001_, _11165_);
  and (_11167_, _11166_, _03384_);
  and (_11168_, _11167_, _11164_);
  or (_11169_, _11168_, _10787_);
  or (_11170_, _10786_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_11171_, _11170_, _10970_);
  and (_11172_, _11171_, _11169_);
  nand (_11173_, _10193_, _01989_);
  or (_11174_, _10352_, _01989_);
  and (_11175_, _11174_, _11173_);
  and (_11176_, _11175_, _05390_);
  and (_11177_, _11176_, _10974_);
  or (_38644_, _11177_, _11172_);
  not (_11178_, _05211_);
  and (_11179_, _05121_, _11178_);
  nor (_11180_, _05121_, _11178_);
  or (_11181_, _11180_, _11179_);
  and (_11182_, _11181_, _03084_);
  and (_11183_, _04525_, _03624_);
  nor (_11184_, _04525_, _03624_);
  or (_11185_, _11184_, _11183_);
  or (_11186_, _11185_, _04973_);
  and (_11187_, _04308_, _02494_);
  nor (_11188_, _04308_, _02494_);
  nor (_11189_, _11188_, _11187_);
  and (_11190_, _11189_, _03060_);
  nand (_11191_, _03624_, _02035_);
  nor (_11192_, _08949_, _04179_);
  or (_11193_, _11192_, _04505_);
  nand (_11194_, _08949_, _08506_);
  or (_11195_, _11194_, _04519_);
  and (_11196_, _04308_, _04208_);
  and (_11197_, _11196_, _04642_);
  nor (_11198_, _04643_, _04308_);
  nor (_11199_, _11198_, _11197_);
  nor (_11200_, _11199_, _03165_);
  or (_11201_, _11185_, _04534_);
  nor (_11202_, _01747_, _01702_);
  and (_11203_, _01747_, \oc8051_golden_model_1.ACC [2]);
  nor (_11204_, _11203_, _11202_);
  and (_11205_, _11204_, _04534_);
  nor (_11206_, _11205_, _03007_);
  and (_11207_, _11206_, _11201_);
  or (_11208_, _11207_, _03005_);
  or (_11209_, _11208_, _11200_);
  and (_11210_, _11209_, _11195_);
  or (_11211_, _11210_, _03446_);
  nor (_11212_, _01745_, _01701_);
  nor (_11213_, _11212_, _03015_);
  and (_11214_, _11213_, _11211_);
  and (_11215_, _03625_, _03015_);
  or (_11216_, _11215_, _03024_);
  or (_11217_, _11216_, _11214_);
  and (_11218_, _11217_, _11193_);
  or (_11219_, _11218_, _02052_);
  nand (_11220_, _07068_, _02052_);
  and (_11221_, _11220_, _02050_);
  and (_11222_, _11221_, _11219_);
  not (_11223_, _08950_);
  and (_11224_, _11194_, _11223_);
  and (_11225_, _11224_, _02049_);
  or (_11226_, _11225_, _11222_);
  and (_11227_, _11226_, _01750_);
  or (_11228_, _01750_, _01702_);
  nand (_11229_, _02144_, _11228_);
  or (_11230_, _11229_, _11227_);
  nand (_11231_, _07068_, _02145_);
  and (_11232_, _11231_, _11230_);
  or (_11233_, _11232_, _03041_);
  and (_11234_, _05211_, _03835_);
  nand (_11235_, _07067_, _03041_);
  or (_11236_, _11235_, _11234_);
  and (_11237_, _11236_, _11233_);
  or (_11238_, _11237_, _03040_);
  nor (_11239_, _08529_, _04179_);
  and (_11240_, _04179_, \oc8051_golden_model_1.PSW [7]);
  nor (_11241_, _11240_, _11239_);
  nand (_11242_, _11241_, _03040_);
  and (_11243_, _11242_, _04460_);
  and (_11244_, _11243_, _11238_);
  and (_11245_, _01767_, _01701_);
  or (_11246_, _02035_, _11245_);
  or (_11247_, _11246_, _11244_);
  and (_11248_, _11247_, _11191_);
  or (_11249_, _11248_, _02033_);
  or (_11250_, _05211_, _04712_);
  and (_11251_, _11250_, _02039_);
  and (_11252_, _11251_, _11249_);
  nor (_11253_, _04716_, _03624_);
  and (_11254_, _04882_, \oc8051_golden_model_1.P1INREG [2]);
  not (_11255_, _11254_);
  and (_11256_, _04875_, \oc8051_golden_model_1.P0INREG [2]);
  not (_11257_, _11256_);
  and (_11258_, _04885_, \oc8051_golden_model_1.P2INREG [2]);
  and (_11259_, _08088_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_11260_, _11259_, _11258_);
  and (_11261_, _11260_, _11257_);
  and (_11262_, _11261_, _11255_);
  and (_11263_, _04849_, \oc8051_golden_model_1.TL0 [2]);
  and (_11264_, _04852_, \oc8051_golden_model_1.SP [2]);
  nor (_11265_, _11264_, _11263_);
  and (_11266_, _11265_, _11262_);
  and (_11267_, _04818_, \oc8051_golden_model_1.IP [2]);
  and (_11268_, _04824_, \oc8051_golden_model_1.B [2]);
  nor (_11269_, _11268_, _11267_);
  and (_11270_, _04829_, \oc8051_golden_model_1.ACC [2]);
  and (_11271_, _04833_, \oc8051_golden_model_1.PSW [2]);
  nor (_11272_, _11271_, _11270_);
  and (_11273_, _11272_, _11269_);
  and (_11274_, _04891_, \oc8051_golden_model_1.IE [2]);
  and (_11275_, _04894_, \oc8051_golden_model_1.SBUF [2]);
  and (_11276_, _04896_, \oc8051_golden_model_1.SCON [2]);
  or (_11277_, _11276_, _11275_);
  nor (_11278_, _11277_, _11274_);
  and (_11279_, _11278_, _11273_);
  and (_11280_, _11279_, _11266_);
  and (_11281_, _04857_, \oc8051_golden_model_1.TH0 [2]);
  and (_11282_, _04861_, \oc8051_golden_model_1.TL1 [2]);
  nor (_11283_, _11282_, _11281_);
  and (_11284_, _04864_, \oc8051_golden_model_1.TCON [2]);
  and (_11285_, _04868_, \oc8051_golden_model_1.PCON [2]);
  nor (_11286_, _11285_, _11284_);
  and (_11287_, _11286_, _11283_);
  and (_11288_, _04902_, \oc8051_golden_model_1.DPH [2]);
  and (_11289_, _04900_, \oc8051_golden_model_1.TMOD [2]);
  nor (_11290_, _11289_, _11288_);
  and (_11291_, _04872_, \oc8051_golden_model_1.DPL [2]);
  and (_11292_, _04843_, \oc8051_golden_model_1.TH1 [2]);
  nor (_11293_, _11292_, _11291_);
  and (_11294_, _11293_, _11290_);
  and (_11295_, _11294_, _11287_);
  and (_11296_, _11295_, _11280_);
  not (_11297_, _11296_);
  nor (_11298_, _11297_, _11253_);
  nor (_11299_, _11298_, _02039_);
  or (_11300_, _11299_, _04920_);
  or (_11301_, _11300_, _11252_);
  and (_11302_, _04920_, _02452_);
  nor (_11303_, _11302_, _01996_);
  and (_11304_, _11303_, _11301_);
  and (_11305_, _04866_, _01996_);
  or (_11306_, _11305_, _01718_);
  or (_11307_, _11306_, _11304_);
  and (_11308_, _01718_, _01702_);
  nor (_11309_, _11308_, _03060_);
  and (_11310_, _11309_, _11307_);
  or (_11311_, _11310_, _11190_);
  and (_11312_, _11311_, _04938_);
  nor (_11313_, _04308_, _06383_);
  and (_11314_, _04308_, _06383_);
  nor (_11315_, _11314_, _11313_);
  and (_11316_, _11315_, _03062_);
  or (_11317_, _11316_, _11312_);
  and (_11318_, _11317_, _04937_);
  and (_11319_, _11188_, _03064_);
  or (_11320_, _11319_, _11318_);
  and (_11321_, _11320_, _04949_);
  and (_11322_, _11313_, _03066_);
  or (_11323_, _11322_, _01728_);
  or (_11324_, _11323_, _11321_);
  and (_11325_, _01728_, _01702_);
  nor (_11326_, _11325_, _04954_);
  and (_11327_, _11326_, _11324_);
  nor (_11328_, _11187_, _04960_);
  or (_11329_, _11328_, _04959_);
  or (_11330_, _11329_, _11327_);
  nand (_11331_, _11314_, _04959_);
  and (_11332_, _11331_, _04964_);
  and (_11333_, _11332_, _11330_);
  nand (_11334_, _01726_, _01701_);
  nand (_11335_, _04973_, _11334_);
  or (_11336_, _11335_, _11333_);
  and (_11337_, _11336_, _11186_);
  or (_11338_, _11337_, _04979_);
  or (_11339_, _11185_, _03275_);
  and (_11340_, _11339_, _04984_);
  and (_11341_, _11340_, _11338_);
  or (_11342_, _11341_, _11182_);
  and (_11343_, _11342_, _04983_);
  nor (_11344_, _11199_, _04983_);
  or (_11345_, _11344_, _01989_);
  or (_11346_, _11345_, _11343_);
  nand (_11347_, _10224_, _01989_);
  and (_11348_, _11347_, _10738_);
  and (_11349_, _11348_, _11346_);
  and (_11350_, _01733_, _01701_);
  or (_11351_, _01992_, _11350_);
  or (_11352_, _11351_, _11349_);
  or (_11353_, _11239_, _03377_);
  and (_11354_, _11353_, _10951_);
  and (_11355_, _11354_, _11352_);
  or (_11356_, _05344_, _03625_);
  nor (_11357_, _10951_, _06686_);
  and (_11358_, _11357_, _11356_);
  or (_11359_, _11358_, _02785_);
  or (_11360_, _11359_, _11355_);
  nor (_11361_, _05364_, _05211_);
  nor (_11362_, _11361_, _06972_);
  or (_11363_, _11362_, _05363_);
  and (_11364_, _11363_, _11360_);
  or (_11365_, _11364_, _03098_);
  nor (_11366_, _04309_, _04258_);
  nor (_11367_, _11366_, _04310_);
  or (_11368_, _11367_, _11165_);
  and (_11369_, _11368_, _03384_);
  and (_11370_, _11369_, _11365_);
  or (_11371_, _11370_, _10787_);
  or (_11372_, _10786_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_11373_, _11372_, _10970_);
  and (_11374_, _11373_, _11371_);
  nand (_11375_, _10186_, _01989_);
  or (_11376_, _10346_, _01989_);
  and (_11377_, _11376_, _11375_);
  and (_11378_, _11377_, _05390_);
  and (_11379_, _11378_, _10974_);
  or (_38646_, _11379_, _11374_);
  or (_11380_, _06686_, _06685_);
  nor (_11381_, _10951_, _05346_);
  and (_11382_, _11381_, _11380_);
  nand (_11383_, _03434_, _02035_);
  nor (_11384_, _11183_, _03434_);
  or (_11385_, _11384_, _04527_);
  or (_11386_, _11385_, _04534_);
  nor (_11387_, _02264_, _01747_);
  nand (_11388_, _01747_, \oc8051_golden_model_1.ACC [3]);
  nand (_11389_, _11388_, _04534_);
  or (_11390_, _11389_, _11387_);
  and (_11391_, _11390_, _11386_);
  and (_11392_, _11391_, _03165_);
  nor (_11393_, _11197_, _04152_);
  nor (_11394_, _11393_, _04645_);
  nor (_11395_, _11394_, _03165_);
  or (_11396_, _11395_, _11392_);
  or (_11397_, _11396_, _03005_);
  nand (_11398_, _09009_, _08637_);
  or (_11399_, _11398_, _04519_);
  and (_11400_, _11399_, _11397_);
  or (_11401_, _11400_, _03446_);
  nor (_11402_, _01825_, _01745_);
  nor (_11403_, _11402_, _03015_);
  and (_11404_, _11403_, _11401_);
  and (_11405_, _06685_, _03015_);
  or (_11406_, _11405_, _03024_);
  or (_11407_, _11406_, _11404_);
  nor (_11408_, _09009_, _04201_);
  or (_11409_, _11408_, _04505_);
  and (_11410_, _11409_, _11407_);
  or (_11411_, _11410_, _02052_);
  nand (_11412_, _07056_, _02052_);
  and (_11413_, _11412_, _02050_);
  and (_11414_, _11413_, _11411_);
  not (_11415_, _09010_);
  and (_11416_, _11398_, _11415_);
  and (_11417_, _11416_, _02049_);
  or (_11418_, _11417_, _11414_);
  and (_11419_, _11418_, _01750_);
  or (_11420_, _02264_, _01750_);
  nand (_11421_, _02144_, _11420_);
  or (_11422_, _11421_, _11419_);
  nand (_11423_, _07056_, _02145_);
  and (_11424_, _11423_, _11422_);
  or (_11425_, _11424_, _03041_);
  and (_11426_, _05166_, _03835_);
  nand (_11427_, _07055_, _03041_);
  or (_11428_, _11427_, _11426_);
  and (_11429_, _11428_, _11425_);
  or (_11430_, _11429_, _03040_);
  and (_11431_, _04201_, \oc8051_golden_model_1.PSW [7]);
  nor (_11432_, _08660_, _04201_);
  nor (_11433_, _11432_, _11431_);
  nand (_11434_, _11433_, _03040_);
  and (_11435_, _11434_, _04460_);
  and (_11436_, _11435_, _11430_);
  and (_11437_, _01825_, _01767_);
  or (_11438_, _02035_, _11437_);
  or (_11439_, _11438_, _11436_);
  and (_11440_, _11439_, _11383_);
  or (_11441_, _11440_, _02033_);
  or (_11442_, _05166_, _04712_);
  and (_11443_, _11442_, _02039_);
  and (_11444_, _11443_, _11441_);
  nor (_11445_, _04716_, _03434_);
  and (_11446_, _04882_, \oc8051_golden_model_1.P1INREG [3]);
  not (_11447_, _11446_);
  and (_11448_, _04875_, \oc8051_golden_model_1.P0INREG [3]);
  not (_11449_, _11448_);
  and (_11450_, _04885_, \oc8051_golden_model_1.P2INREG [3]);
  and (_11451_, _08088_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_11452_, _11451_, _11450_);
  and (_11453_, _11452_, _11449_);
  and (_11454_, _11453_, _11447_);
  and (_11455_, _04849_, \oc8051_golden_model_1.TL0 [3]);
  and (_11456_, _04852_, \oc8051_golden_model_1.SP [3]);
  nor (_11457_, _11456_, _11455_);
  and (_11458_, _11457_, _11454_);
  and (_11459_, _04818_, \oc8051_golden_model_1.IP [3]);
  and (_11460_, _04824_, \oc8051_golden_model_1.B [3]);
  nor (_11461_, _11460_, _11459_);
  and (_11462_, _04829_, \oc8051_golden_model_1.ACC [3]);
  and (_11463_, _04833_, \oc8051_golden_model_1.PSW [3]);
  nor (_11464_, _11463_, _11462_);
  and (_11465_, _11464_, _11461_);
  and (_11466_, _04891_, \oc8051_golden_model_1.IE [3]);
  and (_11467_, _04894_, \oc8051_golden_model_1.SBUF [3]);
  and (_11468_, _04896_, \oc8051_golden_model_1.SCON [3]);
  or (_11469_, _11468_, _11467_);
  nor (_11470_, _11469_, _11466_);
  and (_11471_, _11470_, _11465_);
  and (_11472_, _11471_, _11458_);
  and (_11473_, _04857_, \oc8051_golden_model_1.TH0 [3]);
  and (_11474_, _04861_, \oc8051_golden_model_1.TL1 [3]);
  nor (_11475_, _11474_, _11473_);
  and (_11476_, _04864_, \oc8051_golden_model_1.TCON [3]);
  and (_11477_, _04868_, \oc8051_golden_model_1.PCON [3]);
  nor (_11478_, _11477_, _11476_);
  and (_11479_, _11478_, _11475_);
  and (_11480_, _04902_, \oc8051_golden_model_1.DPH [3]);
  and (_11481_, _04900_, \oc8051_golden_model_1.TMOD [3]);
  nor (_11482_, _11481_, _11480_);
  and (_11483_, _04872_, \oc8051_golden_model_1.DPL [3]);
  and (_11484_, _04843_, \oc8051_golden_model_1.TH1 [3]);
  nor (_11485_, _11484_, _11483_);
  and (_11486_, _11485_, _11482_);
  and (_11487_, _11486_, _11479_);
  and (_11488_, _11487_, _11472_);
  not (_11489_, _11488_);
  nor (_11490_, _11489_, _11445_);
  nor (_11491_, _11490_, _02039_);
  or (_11492_, _11491_, _04920_);
  or (_11493_, _11492_, _11444_);
  and (_11494_, _04920_, _01983_);
  nor (_11495_, _11494_, _01996_);
  and (_11496_, _11495_, _11493_);
  and (_11497_, _04719_, _01996_);
  or (_11498_, _11497_, _01718_);
  or (_11499_, _11498_, _11496_);
  and (_11500_, _02264_, _01718_);
  nor (_11501_, _11500_, _03060_);
  and (_11502_, _11501_, _11499_);
  and (_11503_, _04152_, _02324_);
  nor (_11504_, _04152_, _02324_);
  nor (_11505_, _11504_, _11503_);
  and (_11506_, _11505_, _03060_);
  or (_11507_, _11506_, _11502_);
  and (_11508_, _11507_, _04938_);
  nor (_11509_, _04152_, _06377_);
  and (_11510_, _04152_, _06377_);
  nor (_11511_, _11510_, _11509_);
  and (_11512_, _11511_, _03062_);
  or (_11513_, _11512_, _11508_);
  and (_11514_, _11513_, _04937_);
  and (_11515_, _11504_, _03064_);
  or (_11516_, _11515_, _11514_);
  and (_11517_, _11516_, _04949_);
  and (_11518_, _11509_, _03066_);
  or (_11519_, _11518_, _01728_);
  or (_11520_, _11519_, _11517_);
  and (_11521_, _02264_, _01728_);
  nor (_11522_, _11521_, _04954_);
  and (_11523_, _11522_, _11520_);
  nor (_11524_, _11503_, _04960_);
  or (_11525_, _11524_, _04959_);
  or (_11526_, _11525_, _11523_);
  nand (_11527_, _11510_, _04959_);
  and (_11528_, _11527_, _04964_);
  and (_11529_, _11528_, _11526_);
  and (_11530_, _01825_, _01726_);
  or (_11531_, _10720_, _11530_);
  or (_11532_, _11531_, _11529_);
  not (_11533_, _03273_);
  and (_11534_, _11385_, _11533_);
  or (_11535_, _11534_, _10721_);
  and (_11536_, _11535_, _11532_);
  and (_11537_, _02765_, _01630_);
  and (_11538_, _11385_, _11537_);
  or (_11539_, _11538_, _03084_);
  or (_11540_, _11539_, _11536_);
  not (_11541_, _05166_);
  nor (_11542_, _11179_, _11541_);
  or (_11543_, _05213_, _04984_);
  or (_11544_, _11543_, _11542_);
  and (_11545_, _11544_, _04983_);
  and (_11546_, _11545_, _11540_);
  nor (_11547_, _11394_, _04983_);
  or (_11548_, _11547_, _01989_);
  or (_11549_, _11548_, _11546_);
  nand (_11550_, _10219_, _01989_);
  and (_11551_, _11550_, _10738_);
  and (_11552_, _11551_, _11549_);
  and (_11553_, _01825_, _01733_);
  or (_11554_, _01992_, _11553_);
  or (_11555_, _11554_, _11552_);
  or (_11556_, _11432_, _03377_);
  and (_11557_, _11556_, _10951_);
  and (_11558_, _11557_, _11555_);
  or (_11559_, _11558_, _11382_);
  and (_11560_, _11559_, _05363_);
  or (_11561_, _06972_, _05166_);
  nor (_11562_, _05366_, _05363_);
  and (_11563_, _11562_, _11561_);
  or (_11564_, _11563_, _03098_);
  or (_11565_, _11564_, _11560_);
  nor (_11566_, _04310_, _04153_);
  nor (_11567_, _11566_, _04311_);
  or (_11568_, _11567_, _11165_);
  and (_11569_, _11568_, _03384_);
  and (_11570_, _11569_, _11565_);
  and (_11571_, _11570_, _10785_);
  nor (_11572_, _10786_, _03388_);
  or (_11573_, _11572_, _10969_);
  or (_11574_, _11573_, _11571_);
  nand (_11575_, _10180_, _01989_);
  or (_11576_, _10341_, _01989_);
  and (_11577_, _11576_, _11575_);
  or (_11578_, _11577_, _10970_);
  and (_38647_, _11578_, _11574_);
  or (_11579_, _05346_, _05343_);
  nor (_11580_, _10951_, _05347_);
  and (_11581_, _11580_, _11579_);
  nor (_11582_, _04527_, _04372_);
  and (_11583_, _04527_, _04372_);
  or (_11584_, _11583_, _11582_);
  or (_11585_, _11584_, _04973_);
  nor (_11586_, _04419_, _06283_);
  and (_11587_, _04419_, _06283_);
  nor (_11588_, _11587_, _11586_);
  and (_11589_, _11588_, _03062_);
  and (_11590_, _04784_, _04419_);
  nor (_11591_, _04784_, _04419_);
  nor (_11592_, _11591_, _11590_);
  and (_11593_, _11592_, _03060_);
  and (_11594_, _10373_, _01767_);
  nor (_11595_, _08556_, _08973_);
  or (_11596_, _11595_, _04505_);
  nand (_11597_, _08557_, _08973_);
  or (_11598_, _11597_, _04519_);
  and (_11599_, _11584_, _04535_);
  and (_11600_, _01747_, \oc8051_golden_model_1.ACC [4]);
  nor (_11601_, _10374_, _01747_);
  or (_11602_, _11601_, _11600_);
  and (_11603_, _11602_, _04534_);
  or (_11604_, _11603_, _02079_);
  or (_11605_, _11604_, _11599_);
  or (_11606_, _05303_, _04550_);
  and (_11607_, _11606_, _11605_);
  or (_11608_, _11607_, _03007_);
  and (_11609_, _04645_, _04419_);
  nor (_11610_, _04645_, _04419_);
  nor (_11611_, _11610_, _11609_);
  nand (_11612_, _11611_, _03007_);
  and (_11613_, _11612_, _11608_);
  or (_11614_, _11613_, _03005_);
  and (_11615_, _11614_, _11598_);
  or (_11616_, _11615_, _03446_);
  nor (_11617_, _10373_, _01745_);
  nor (_11618_, _11617_, _03015_);
  and (_11619_, _11618_, _11616_);
  and (_11620_, _05343_, _03015_);
  or (_11621_, _11620_, _03024_);
  or (_11622_, _11621_, _11619_);
  and (_11623_, _11622_, _11596_);
  or (_11624_, _11623_, _02052_);
  nand (_11625_, _07126_, _02052_);
  and (_11626_, _11625_, _02050_);
  and (_11627_, _11626_, _11624_);
  not (_11628_, _08974_);
  and (_11629_, _11597_, _11628_);
  and (_11630_, _11629_, _02049_);
  or (_11631_, _11630_, _11627_);
  and (_11632_, _11631_, _01750_);
  or (_11633_, _10374_, _01750_);
  nand (_11634_, _11633_, _02144_);
  or (_11635_, _11634_, _11632_);
  nand (_11636_, _07126_, _02145_);
  and (_11637_, _11636_, _11635_);
  or (_11638_, _11637_, _03041_);
  and (_11639_, _05303_, _03835_);
  nand (_11640_, _07125_, _03041_);
  or (_11641_, _11640_, _11639_);
  and (_11642_, _11641_, _11638_);
  or (_11643_, _11642_, _03040_);
  nor (_11644_, _08580_, _08556_);
  and (_11645_, _08556_, \oc8051_golden_model_1.PSW [7]);
  nor (_11646_, _11645_, _11644_);
  nand (_11647_, _11646_, _03040_);
  and (_11648_, _11647_, _04460_);
  and (_11649_, _11648_, _11643_);
  or (_11650_, _11649_, _11594_);
  and (_11651_, _11650_, _10794_);
  nor (_11652_, _04372_, _10794_);
  or (_11653_, _11652_, _02033_);
  or (_11654_, _11653_, _11651_);
  or (_11655_, _05303_, _04712_);
  and (_11656_, _11655_, _02039_);
  and (_11657_, _11656_, _11654_);
  nor (_11658_, _04716_, _04372_);
  and (_11659_, _04818_, \oc8051_golden_model_1.IP [4]);
  and (_11660_, _04824_, \oc8051_golden_model_1.B [4]);
  nor (_11661_, _11660_, _11659_);
  and (_11662_, _04829_, \oc8051_golden_model_1.ACC [4]);
  and (_11663_, _04833_, \oc8051_golden_model_1.PSW [4]);
  nor (_11664_, _11663_, _11662_);
  and (_11665_, _11664_, _11661_);
  and (_11666_, _04843_, \oc8051_golden_model_1.TH1 [4]);
  not (_11667_, _11666_);
  and (_11668_, _04849_, \oc8051_golden_model_1.TL0 [4]);
  and (_11669_, _04852_, \oc8051_golden_model_1.SP [4]);
  nor (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _11667_);
  and (_11672_, _11671_, _11665_);
  and (_11673_, _04857_, \oc8051_golden_model_1.TH0 [4]);
  and (_11674_, _04861_, \oc8051_golden_model_1.TL1 [4]);
  nor (_11675_, _11674_, _11673_);
  and (_11676_, _04864_, \oc8051_golden_model_1.TCON [4]);
  and (_11677_, _04868_, \oc8051_golden_model_1.PCON [4]);
  nor (_11678_, _11677_, _11676_);
  and (_11679_, _11678_, _11675_);
  and (_11680_, _04872_, \oc8051_golden_model_1.DPL [4]);
  not (_11681_, _11680_);
  and (_11682_, _04875_, \oc8051_golden_model_1.P0INREG [4]);
  not (_11683_, _11682_);
  nand (_11684_, _04879_, \oc8051_golden_model_1.P3INREG [4]);
  and (_11685_, _04882_, \oc8051_golden_model_1.P1INREG [4]);
  and (_11686_, _04885_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_11687_, _11686_, _11685_);
  and (_11688_, _11687_, _11684_);
  and (_11689_, _11688_, _11683_);
  and (_11690_, _11689_, _11681_);
  and (_11691_, _04891_, \oc8051_golden_model_1.IE [4]);
  and (_11692_, _04894_, \oc8051_golden_model_1.SBUF [4]);
  and (_11693_, _04896_, \oc8051_golden_model_1.SCON [4]);
  or (_11694_, _11693_, _11692_);
  nor (_11695_, _11694_, _11691_);
  and (_11696_, _04900_, \oc8051_golden_model_1.TMOD [4]);
  and (_11697_, _04902_, \oc8051_golden_model_1.DPH [4]);
  nor (_11698_, _11697_, _11696_);
  and (_11699_, _11698_, _11695_);
  and (_11700_, _11699_, _11690_);
  and (_11701_, _11700_, _11679_);
  and (_11702_, _11701_, _11672_);
  not (_11703_, _11702_);
  nor (_11704_, _11703_, _11658_);
  nor (_11705_, _11704_, _02039_);
  or (_11706_, _11705_, _04920_);
  or (_11707_, _11706_, _11657_);
  and (_11708_, _04920_, _02825_);
  nor (_11709_, _11708_, _01996_);
  and (_11710_, _11709_, _11707_);
  and (_11711_, _04831_, _01996_);
  or (_11712_, _11711_, _01718_);
  or (_11713_, _11712_, _11710_);
  and (_11714_, _10374_, _01718_);
  nor (_11715_, _11714_, _03060_);
  and (_11716_, _11715_, _11713_);
  or (_11717_, _11716_, _11593_);
  and (_11718_, _11717_, _04938_);
  or (_11719_, _11718_, _11589_);
  and (_11720_, _11719_, _04937_);
  and (_11721_, _11591_, _03064_);
  or (_11722_, _11721_, _11720_);
  and (_11723_, _11722_, _04949_);
  and (_11724_, _11586_, _03066_);
  or (_11725_, _11724_, _01728_);
  or (_11726_, _11725_, _11723_);
  and (_11727_, _10374_, _01728_);
  nor (_11728_, _11727_, _04954_);
  and (_11729_, _11728_, _11726_);
  nor (_11730_, _11590_, _04960_);
  or (_11731_, _11730_, _04959_);
  or (_11732_, _11731_, _11729_);
  nand (_11733_, _11587_, _04959_);
  and (_11734_, _11733_, _04964_);
  and (_11735_, _11734_, _11732_);
  nand (_11736_, _10373_, _01726_);
  nand (_11737_, _11736_, _04973_);
  or (_11738_, _11737_, _11735_);
  and (_11739_, _11738_, _11585_);
  or (_11740_, _11739_, _04979_);
  or (_11741_, _11584_, _03275_);
  and (_11742_, _11741_, _04984_);
  and (_11743_, _11742_, _11740_);
  not (_11744_, _05303_);
  and (_11745_, _05213_, _11744_);
  nor (_11746_, _05213_, _11744_);
  or (_11747_, _11746_, _11745_);
  and (_11748_, _11747_, _03084_);
  or (_11749_, _11748_, _11743_);
  and (_11750_, _11749_, _04983_);
  nor (_11751_, _11611_, _04983_);
  or (_11752_, _11751_, _01989_);
  or (_11753_, _11752_, _11750_);
  nand (_11754_, _10215_, _01989_);
  and (_11755_, _11754_, _10738_);
  and (_11756_, _11755_, _11753_);
  and (_11757_, _10373_, _01733_);
  or (_11758_, _11757_, _01992_);
  or (_11759_, _11758_, _11756_);
  or (_11760_, _11644_, _03377_);
  and (_11761_, _11760_, _10951_);
  and (_11762_, _11761_, _11759_);
  or (_11763_, _11762_, _11581_);
  and (_11764_, _11763_, _05363_);
  or (_11765_, _05366_, _05303_);
  nor (_11766_, _06954_, _05363_);
  and (_11767_, _11766_, _11765_);
  or (_11768_, _11767_, _03098_);
  or (_11769_, _11768_, _11764_);
  nor (_11770_, _04420_, _04311_);
  nor (_11771_, _11770_, _04421_);
  or (_11772_, _11771_, _11165_);
  and (_11773_, _11772_, _03384_);
  and (_11774_, _11773_, _11769_);
  or (_11775_, _11774_, _10787_);
  or (_11776_, _10786_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_11777_, _11776_, _10970_);
  and (_11778_, _11777_, _11775_);
  nand (_11779_, _10174_, _01989_);
  or (_11780_, _10338_, _01989_);
  and (_11781_, _11780_, _11779_);
  and (_11782_, _11781_, _05390_);
  and (_11783_, _11782_, _10974_);
  or (_38649_, _11783_, _11778_);
  nor (_11784_, _04103_, _06277_);
  and (_11785_, _04103_, _06277_);
  nor (_11786_, _11785_, _11784_);
  and (_11787_, _11786_, _03062_);
  nand (_11788_, _04057_, _02035_);
  nand (_11789_, _08663_, _09020_);
  or (_11790_, _11789_, _04519_);
  or (_11791_, _05258_, _04550_);
  nor (_11792_, _11583_, _04057_);
  or (_11793_, _11792_, _04528_);
  and (_11794_, _11793_, _04535_);
  and (_11795_, _01747_, \oc8051_golden_model_1.ACC [5]);
  nor (_11796_, _10369_, _01747_);
  or (_11797_, _11796_, _11795_);
  and (_11798_, _11797_, _04534_);
  or (_11799_, _11798_, _02079_);
  or (_11800_, _11799_, _11794_);
  and (_11801_, _11800_, _11791_);
  or (_11802_, _11801_, _03007_);
  nor (_11803_, _11609_, _04103_);
  nor (_11804_, _11803_, _04646_);
  nand (_11805_, _11804_, _03007_);
  and (_11806_, _11805_, _11802_);
  or (_11807_, _11806_, _03005_);
  and (_11808_, _11807_, _11790_);
  or (_11809_, _11808_, _03446_);
  nor (_11810_, _10368_, _01745_);
  nor (_11811_, _11810_, _03015_);
  and (_11812_, _11811_, _11809_);
  and (_11813_, _05342_, _03015_);
  or (_11814_, _11813_, _03024_);
  or (_11815_, _11814_, _11812_);
  nor (_11816_, _08662_, _09020_);
  or (_11817_, _11816_, _04505_);
  and (_11818_, _11817_, _11815_);
  or (_11819_, _11818_, _02052_);
  nand (_11820_, _07115_, _02052_);
  and (_11821_, _11820_, _02050_);
  and (_11822_, _11821_, _11819_);
  not (_11823_, _09021_);
  and (_11824_, _11789_, _11823_);
  and (_11825_, _11824_, _02049_);
  or (_11826_, _11825_, _11822_);
  and (_11827_, _11826_, _01750_);
  or (_11828_, _10369_, _01750_);
  nand (_11829_, _11828_, _02144_);
  or (_11830_, _11829_, _11827_);
  nand (_11831_, _07115_, _02145_);
  and (_11832_, _11831_, _11830_);
  or (_11833_, _11832_, _03041_);
  and (_11834_, _05258_, _03835_);
  nand (_11835_, _07114_, _03041_);
  or (_11836_, _11835_, _11834_);
  and (_11837_, _11836_, _11833_);
  or (_11838_, _11837_, _03040_);
  nor (_11839_, _08686_, _08662_);
  and (_11840_, _08662_, \oc8051_golden_model_1.PSW [7]);
  nor (_11841_, _11840_, _11839_);
  nand (_11842_, _11841_, _03040_);
  and (_11843_, _11842_, _04460_);
  and (_11844_, _11843_, _11838_);
  and (_11845_, _10368_, _01767_);
  or (_11846_, _11845_, _02035_);
  or (_11847_, _11846_, _11844_);
  and (_11848_, _11847_, _11788_);
  or (_11849_, _11848_, _02033_);
  or (_11850_, _05258_, _04712_);
  and (_11851_, _11850_, _02039_);
  and (_11852_, _11851_, _11849_);
  nor (_11853_, _04716_, _04057_);
  and (_11854_, _04818_, \oc8051_golden_model_1.IP [5]);
  and (_11855_, _04824_, \oc8051_golden_model_1.B [5]);
  nor (_11856_, _11855_, _11854_);
  and (_11857_, _04829_, \oc8051_golden_model_1.ACC [5]);
  and (_11858_, _04833_, \oc8051_golden_model_1.PSW [5]);
  nor (_11859_, _11858_, _11857_);
  and (_11860_, _11859_, _11856_);
  and (_11861_, _04852_, \oc8051_golden_model_1.SP [5]);
  not (_11862_, _11861_);
  and (_11863_, _04872_, \oc8051_golden_model_1.DPL [5]);
  and (_11864_, _04851_, _04718_);
  and (_11865_, _11864_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_11866_, _11865_, _11863_);
  and (_11867_, _11866_, _11862_);
  and (_11868_, _11867_, _11860_);
  and (_11869_, _04879_, \oc8051_golden_model_1.P3INREG [5]);
  not (_11870_, _11869_);
  and (_11871_, _04882_, \oc8051_golden_model_1.P1INREG [5]);
  and (_11872_, _04885_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_11873_, _11872_, _11871_);
  and (_11874_, _11873_, _11870_);
  and (_11875_, _04891_, \oc8051_golden_model_1.IE [5]);
  not (_11876_, _11875_);
  and (_11877_, _04896_, \oc8051_golden_model_1.SCON [5]);
  and (_11878_, _04894_, \oc8051_golden_model_1.SBUF [5]);
  nor (_11879_, _11878_, _11877_);
  and (_11880_, _11879_, _11876_);
  and (_11881_, _11880_, _11874_);
  and (_11882_, _04902_, \oc8051_golden_model_1.DPH [5]);
  and (_11883_, _04900_, \oc8051_golden_model_1.TMOD [5]);
  nor (_11884_, _11883_, _11882_);
  and (_11885_, _04843_, \oc8051_golden_model_1.TH1 [5]);
  and (_11886_, _04849_, \oc8051_golden_model_1.TL0 [5]);
  nor (_11887_, _11886_, _11885_);
  and (_11888_, _11887_, _11884_);
  and (_11889_, _04857_, \oc8051_golden_model_1.TH0 [5]);
  and (_11890_, _04861_, \oc8051_golden_model_1.TL1 [5]);
  nor (_11891_, _11890_, _11889_);
  and (_11892_, _04864_, \oc8051_golden_model_1.TCON [5]);
  and (_11893_, _04868_, \oc8051_golden_model_1.PCON [5]);
  nor (_11894_, _11893_, _11892_);
  and (_11895_, _11894_, _11891_);
  and (_11896_, _11895_, _11888_);
  and (_11897_, _11896_, _11881_);
  and (_11898_, _11897_, _11868_);
  not (_11899_, _11898_);
  nor (_11900_, _11899_, _11853_);
  nor (_11901_, _11900_, _02039_);
  or (_11902_, _11901_, _04920_);
  or (_11903_, _11902_, _11852_);
  and (_11904_, _04920_, _02410_);
  nor (_11905_, _11904_, _01996_);
  and (_11906_, _11905_, _11903_);
  and (_11907_, _04827_, _01996_);
  or (_11908_, _11907_, _01718_);
  or (_11909_, _11908_, _11906_);
  and (_11910_, _10369_, _01718_);
  nor (_11911_, _11910_, _03060_);
  and (_11912_, _11911_, _11909_);
  and (_11913_, _04815_, _04103_);
  nor (_11914_, _04815_, _04103_);
  nor (_11915_, _11914_, _11913_);
  and (_11916_, _11915_, _03060_);
  or (_11917_, _11916_, _11912_);
  and (_11918_, _11917_, _04938_);
  or (_11919_, _11918_, _11787_);
  and (_11920_, _11919_, _04937_);
  and (_11921_, _11914_, _03064_);
  or (_11922_, _11921_, _03066_);
  or (_11923_, _11922_, _11920_);
  or (_11924_, _11784_, _04949_);
  and (_11925_, _11924_, _11923_);
  or (_11926_, _11925_, _01728_);
  and (_11927_, _10369_, _01728_);
  nor (_11928_, _11927_, _04954_);
  and (_11929_, _11928_, _11926_);
  nor (_11930_, _11913_, _04960_);
  or (_11931_, _11930_, _04959_);
  or (_11932_, _11931_, _11929_);
  nand (_11933_, _11785_, _04959_);
  and (_11934_, _11933_, _04964_);
  and (_11935_, _11934_, _11932_);
  and (_11936_, _10368_, _01726_);
  or (_11937_, _11936_, _10720_);
  or (_11938_, _11937_, _11935_);
  and (_11939_, _11793_, _11533_);
  or (_11940_, _11939_, _10721_);
  and (_11941_, _11940_, _11938_);
  and (_11942_, _11793_, _11537_);
  or (_11943_, _11942_, _03084_);
  or (_11944_, _11943_, _11941_);
  not (_11945_, _05258_);
  nor (_11946_, _11745_, _11945_);
  or (_11947_, _05305_, _04984_);
  or (_11948_, _11947_, _11946_);
  and (_11949_, _11948_, _04983_);
  and (_11950_, _11949_, _11944_);
  nor (_11951_, _11804_, _04983_);
  or (_11952_, _11951_, _01989_);
  or (_11953_, _11952_, _11950_);
  nand (_11954_, _10210_, _01989_);
  and (_11955_, _11954_, _10738_);
  and (_11956_, _11955_, _11953_);
  and (_11957_, _10368_, _01733_);
  or (_11958_, _11957_, _01992_);
  or (_11959_, _11958_, _11956_);
  or (_11960_, _11839_, _03377_);
  and (_11961_, _11960_, _10951_);
  and (_11962_, _11961_, _11959_);
  nor (_11963_, _05347_, _05342_);
  nor (_11964_, _11963_, _05348_);
  and (_11965_, _11964_, _10980_);
  or (_11966_, _11965_, _11962_);
  and (_11967_, _11966_, _05363_);
  or (_11968_, _06954_, _05258_);
  nor (_11969_, _05368_, _05363_);
  and (_11970_, _11969_, _11968_);
  or (_11971_, _11970_, _03098_);
  or (_11972_, _11971_, _11967_);
  nor (_11973_, _04421_, _04104_);
  nor (_11974_, _11973_, _04422_);
  or (_11975_, _11974_, _11165_);
  and (_11976_, _11975_, _03384_);
  and (_11977_, _11976_, _11972_);
  or (_11978_, _11977_, _10787_);
  or (_11979_, _10786_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_11980_, _11979_, _10970_);
  and (_11981_, _11980_, _11978_);
  not (_11982_, _10334_);
  nor (_11983_, _11982_, _01989_);
  and (_11984_, _10169_, _01989_);
  or (_11985_, _11984_, _11983_);
  and (_11986_, _11985_, _05390_);
  and (_11987_, _11986_, _10974_);
  or (_38650_, _11987_, _11981_);
  and (_11988_, _10360_, _01726_);
  and (_11989_, _10360_, _01767_);
  nand (_11990_, _08611_, _08997_);
  or (_11991_, _11990_, _04519_);
  nor (_11992_, _04646_, _04010_);
  nor (_11993_, _11992_, _04647_);
  nor (_11994_, _11993_, _03165_);
  or (_11995_, _05029_, _04550_);
  nor (_11996_, _04528_, _03964_);
  or (_11997_, _11996_, _04529_);
  and (_11998_, _11997_, _04535_);
  or (_11999_, _10360_, _01747_);
  nand (_12000_, _01747_, _06231_);
  and (_12001_, _12000_, _11999_);
  and (_12002_, _12001_, _04534_);
  or (_12003_, _12002_, _02079_);
  or (_12004_, _12003_, _11998_);
  and (_12005_, _12004_, _03165_);
  and (_12006_, _12005_, _11995_);
  or (_12007_, _12006_, _11994_);
  or (_12008_, _12007_, _03005_);
  and (_12009_, _12008_, _11991_);
  or (_12010_, _12009_, _03446_);
  nor (_12011_, _10360_, _01745_);
  nor (_12012_, _12011_, _03015_);
  and (_12013_, _12012_, _12010_);
  and (_12014_, _06655_, _03015_);
  or (_12015_, _12014_, _03024_);
  or (_12016_, _12015_, _12013_);
  nor (_12017_, _08610_, _08997_);
  or (_12018_, _12017_, _04505_);
  and (_12019_, _12018_, _12016_);
  or (_12020_, _12019_, _02052_);
  nand (_12021_, _07036_, _02052_);
  and (_12022_, _12021_, _02050_);
  and (_12023_, _12022_, _12020_);
  not (_12024_, _08998_);
  and (_12025_, _11990_, _12024_);
  and (_12026_, _12025_, _02049_);
  or (_12027_, _12026_, _12023_);
  and (_12028_, _12027_, _01750_);
  or (_12029_, _10361_, _01750_);
  nand (_12030_, _12029_, _02144_);
  or (_12031_, _12030_, _12028_);
  nand (_12032_, _07036_, _02145_);
  and (_12033_, _12032_, _12031_);
  or (_12034_, _12033_, _03041_);
  and (_12035_, _05029_, _03835_);
  nand (_12036_, _07035_, _03041_);
  or (_12037_, _12036_, _12035_);
  and (_12038_, _12037_, _12034_);
  or (_12039_, _12038_, _03040_);
  nor (_12040_, _08634_, _08610_);
  and (_12041_, _08610_, \oc8051_golden_model_1.PSW [7]);
  nor (_12042_, _12041_, _12040_);
  nand (_12043_, _12042_, _03040_);
  and (_12044_, _12043_, _04460_);
  and (_12045_, _12044_, _12039_);
  or (_12046_, _12045_, _11989_);
  and (_12047_, _12046_, _10794_);
  nor (_12048_, _03964_, _10794_);
  or (_12049_, _12048_, _02033_);
  or (_12050_, _12049_, _12047_);
  or (_12051_, _05029_, _04712_);
  and (_12052_, _12051_, _02039_);
  and (_12053_, _12052_, _12050_);
  nor (_12054_, _04716_, _03964_);
  and (_12055_, _04818_, \oc8051_golden_model_1.IP [6]);
  and (_12056_, _04833_, \oc8051_golden_model_1.PSW [6]);
  or (_12057_, _12056_, _12055_);
  and (_12058_, _04829_, \oc8051_golden_model_1.ACC [6]);
  and (_12059_, _04824_, \oc8051_golden_model_1.B [6]);
  or (_12060_, _12059_, _12058_);
  or (_12061_, _12060_, _12057_);
  and (_12062_, _04843_, \oc8051_golden_model_1.TH1 [6]);
  and (_12063_, _04902_, \oc8051_golden_model_1.DPH [6]);
  or (_12064_, _12063_, _12062_);
  and (_12065_, _04872_, \oc8051_golden_model_1.DPL [6]);
  and (_12066_, _04900_, \oc8051_golden_model_1.TMOD [6]);
  or (_12067_, _12066_, _12065_);
  or (_12068_, _12067_, _12064_);
  or (_12069_, _12068_, _12061_);
  and (_12070_, _04864_, \oc8051_golden_model_1.TCON [6]);
  and (_12071_, _04857_, \oc8051_golden_model_1.TH0 [6]);
  or (_12072_, _12071_, _12070_);
  and (_12073_, _04868_, \oc8051_golden_model_1.PCON [6]);
  and (_12074_, _04861_, \oc8051_golden_model_1.TL1 [6]);
  or (_12075_, _12074_, _12073_);
  or (_12076_, _12075_, _12072_);
  and (_12077_, _04894_, \oc8051_golden_model_1.SBUF [6]);
  and (_12078_, _04896_, \oc8051_golden_model_1.SCON [6]);
  and (_12079_, _04891_, \oc8051_golden_model_1.IE [6]);
  or (_12080_, _12079_, _12078_);
  or (_12081_, _12080_, _12077_);
  and (_12082_, _04875_, \oc8051_golden_model_1.P0INREG [6]);
  and (_12083_, _04882_, \oc8051_golden_model_1.P1INREG [6]);
  and (_12084_, _04885_, \oc8051_golden_model_1.P2INREG [6]);
  and (_12085_, _08088_, \oc8051_golden_model_1.P3INREG [6]);
  or (_12086_, _12085_, _12084_);
  or (_12087_, _12086_, _12083_);
  or (_12088_, _12087_, _12082_);
  and (_12089_, _04849_, \oc8051_golden_model_1.TL0 [6]);
  and (_12090_, _04852_, \oc8051_golden_model_1.SP [6]);
  or (_12091_, _12090_, _12089_);
  or (_12092_, _12091_, _12088_);
  or (_12093_, _12092_, _12081_);
  or (_12094_, _12093_, _12076_);
  or (_12095_, _12094_, _12069_);
  nor (_12096_, _12095_, _12054_);
  nor (_12097_, _12096_, _02039_);
  or (_12098_, _12097_, _04920_);
  or (_12099_, _12098_, _12053_);
  and (_12100_, _04920_, _02118_);
  nor (_12101_, _12100_, _01996_);
  and (_12102_, _12101_, _12099_);
  not (_12103_, _04752_);
  and (_12104_, _12103_, _01996_);
  or (_12105_, _12104_, _01718_);
  or (_12106_, _12105_, _12102_);
  and (_12107_, _10361_, _01718_);
  nor (_12108_, _12107_, _03060_);
  and (_12109_, _12108_, _12106_);
  and (_12110_, _04752_, _04010_);
  nor (_12111_, _04752_, _04010_);
  nor (_12112_, _12111_, _12110_);
  and (_12113_, _12112_, _03060_);
  or (_12114_, _12113_, _12109_);
  and (_12115_, _12114_, _04938_);
  nor (_12116_, _04010_, _06231_);
  and (_12117_, _04010_, _06231_);
  nor (_12118_, _12117_, _12116_);
  and (_12119_, _12118_, _03062_);
  or (_12120_, _12119_, _12115_);
  and (_12121_, _12120_, _04937_);
  and (_12122_, _12111_, _03064_);
  or (_12123_, _12122_, _03066_);
  or (_12124_, _12123_, _12121_);
  or (_12125_, _12116_, _04949_);
  and (_12126_, _12125_, _12124_);
  or (_12127_, _12126_, _01728_);
  and (_12128_, _10361_, _01728_);
  nor (_12129_, _12128_, _04954_);
  and (_12130_, _12129_, _12127_);
  nor (_12131_, _12110_, _04960_);
  or (_12132_, _12131_, _04959_);
  or (_12133_, _12132_, _12130_);
  nand (_12134_, _12117_, _04959_);
  and (_12135_, _12134_, _04964_);
  and (_12136_, _12135_, _12133_);
  or (_12137_, _12136_, _11988_);
  and (_12138_, _12137_, _04973_);
  not (_12139_, _04973_);
  and (_12140_, _11997_, _12139_);
  or (_12141_, _12140_, _04979_);
  or (_12142_, _12141_, _12138_);
  or (_12143_, _11997_, _03275_);
  and (_12144_, _12143_, _04984_);
  and (_12145_, _12144_, _12142_);
  nor (_12146_, _05305_, _05030_);
  or (_12147_, _12146_, _05306_);
  and (_12148_, _12147_, _03084_);
  or (_12149_, _12148_, _12145_);
  and (_12150_, _12149_, _04983_);
  nor (_12151_, _11993_, _04983_);
  or (_12152_, _12151_, _01989_);
  or (_12153_, _12152_, _12150_);
  nand (_12154_, _10202_, _01989_);
  and (_12155_, _12154_, _10738_);
  and (_12156_, _12155_, _12153_);
  and (_12157_, _10360_, _01733_);
  or (_12158_, _12157_, _01992_);
  or (_12159_, _12158_, _12156_);
  or (_12160_, _12040_, _03377_);
  and (_12161_, _12160_, _05337_);
  and (_12162_, _12161_, _12159_);
  and (_12163_, _05348_, _03964_);
  nor (_12164_, _05348_, _03964_);
  or (_12165_, _12164_, _12163_);
  and (_12166_, _12165_, _05338_);
  or (_12167_, _12166_, _03293_);
  or (_12168_, _12167_, _12162_);
  or (_12169_, _12165_, _03292_);
  and (_12170_, _12169_, _05363_);
  and (_12171_, _12170_, _12168_);
  or (_12172_, _05368_, _05029_);
  nor (_12173_, _05369_, _05363_);
  and (_12174_, _12173_, _12172_);
  or (_12175_, _12174_, _03098_);
  or (_12176_, _12175_, _12171_);
  nor (_12177_, _04422_, _04011_);
  nor (_12178_, _12177_, _04423_);
  or (_12179_, _12178_, _11165_);
  and (_12180_, _12179_, _03384_);
  and (_12181_, _12180_, _12176_);
  or (_12182_, _12181_, _10787_);
  or (_12183_, _10786_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_12184_, _12183_, _10970_);
  and (_12185_, _12184_, _12182_);
  nand (_12186_, _10163_, _01989_);
  or (_12187_, _10328_, _01989_);
  and (_12188_, _12187_, _12186_);
  and (_12189_, _12188_, _05390_);
  and (_12190_, _12189_, _10974_);
  or (_38651_, _12190_, _12185_);
  nand (_12191_, _10786_, _05377_);
  or (_12192_, _10786_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_12193_, _12192_, _10970_);
  and (_12194_, _12193_, _12191_);
  and (_12195_, _10974_, _05431_);
  or (_38652_, _12195_, _12194_);
  and (_12196_, _10781_, _03300_);
  and (_12197_, _12196_, _10784_);
  not (_12198_, _12197_);
  or (_12199_, _12198_, _10963_);
  and (_12200_, _05390_, _03437_);
  nand (_12201_, _12200_, _10967_);
  or (_12202_, _12197_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_12203_, _12202_, _12201_);
  and (_12204_, _12203_, _12199_);
  and (_12205_, _10967_, _03437_);
  and (_12206_, _12205_, _10978_);
  or (_38656_, _12206_, _12204_);
  or (_12207_, _12198_, _11168_);
  or (_12208_, _12197_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_12209_, _12208_, _12201_);
  and (_12210_, _12209_, _12207_);
  and (_12211_, _12205_, _11176_);
  or (_38657_, _12211_, _12210_);
  or (_12212_, _12198_, _11370_);
  or (_12213_, _12197_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_12214_, _12213_, _12201_);
  and (_12215_, _12214_, _12212_);
  and (_12216_, _12205_, _11378_);
  or (_38658_, _12216_, _12215_);
  or (_12217_, _12198_, _11570_);
  or (_12218_, _12197_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_12219_, _12218_, _12201_);
  and (_12220_, _12219_, _12217_);
  and (_12221_, _11577_, _05390_);
  and (_12222_, _12205_, _12221_);
  or (_38660_, _12222_, _12220_);
  or (_12223_, _12198_, _11774_);
  or (_12224_, _12197_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_12225_, _12224_, _12201_);
  and (_12226_, _12225_, _12223_);
  and (_12227_, _12205_, _11782_);
  or (_38661_, _12227_, _12226_);
  or (_12228_, _12198_, _11977_);
  or (_12229_, _12197_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_12230_, _12229_, _12201_);
  and (_12231_, _12230_, _12228_);
  and (_12232_, _12205_, _11986_);
  or (_38662_, _12232_, _12231_);
  or (_12233_, _12198_, _12181_);
  or (_12234_, _12197_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_12235_, _12234_, _12201_);
  and (_12236_, _12235_, _12233_);
  and (_12237_, _12205_, _12189_);
  or (_38663_, _12237_, _12236_);
  or (_12238_, _12198_, _05378_);
  or (_12239_, _12197_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_12240_, _12239_, _12201_);
  and (_12241_, _12240_, _12238_);
  and (_12242_, _12205_, _05431_);
  or (_38664_, _12242_, _12241_);
  not (_12243_, _03386_);
  nor (_12244_, _12243_, _03101_);
  and (_12245_, _12244_, _10784_);
  not (_12246_, _12245_);
  or (_12247_, _12246_, _10963_);
  or (_12248_, _12245_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_12249_, _05390_, _04551_);
  nand (_12250_, _12249_, _10967_);
  and (_12251_, _12250_, _12248_);
  and (_12252_, _12251_, _12247_);
  and (_12253_, _10967_, _04551_);
  and (_12254_, _12253_, _10978_);
  or (_38668_, _12254_, _12252_);
  or (_12255_, _12246_, _11168_);
  or (_12256_, _12245_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_12257_, _12256_, _12250_);
  and (_12258_, _12257_, _12255_);
  and (_12259_, _12253_, _11176_);
  or (_38669_, _12259_, _12258_);
  or (_12260_, _12246_, _11370_);
  or (_12261_, _12245_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_12262_, _12261_, _12250_);
  and (_12263_, _12262_, _12260_);
  and (_12264_, _12253_, _11378_);
  or (_38670_, _12264_, _12263_);
  or (_12265_, _12246_, _11570_);
  or (_12266_, _12245_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_12267_, _12266_, _12250_);
  and (_12268_, _12267_, _12265_);
  and (_12269_, _12253_, _12221_);
  or (_38671_, _12269_, _12268_);
  or (_12270_, _12246_, _11774_);
  or (_12271_, _12245_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_12272_, _12271_, _12250_);
  and (_12273_, _12272_, _12270_);
  and (_12274_, _12253_, _11782_);
  or (_38672_, _12274_, _12273_);
  or (_12275_, _12246_, _11977_);
  or (_12276_, _12245_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_12277_, _12276_, _12250_);
  and (_12278_, _12277_, _12275_);
  and (_12279_, _12253_, _11986_);
  or (_38674_, _12279_, _12278_);
  or (_12280_, _12246_, _12181_);
  or (_12281_, _12245_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_12282_, _12281_, _12250_);
  and (_12283_, _12282_, _12280_);
  and (_12284_, _12253_, _12189_);
  or (_38675_, _12284_, _12283_);
  or (_12285_, _12246_, _05378_);
  or (_12286_, _12245_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_12287_, _12286_, _12250_);
  and (_12288_, _12287_, _12285_);
  and (_12289_, _12253_, _05431_);
  or (_38676_, _12289_, _12288_);
  and (_12290_, _10784_, _03387_);
  or (_12291_, _12290_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_12292_, _05390_, _03105_);
  nand (_12293_, _12292_, _10967_);
  and (_12294_, _12293_, _12291_);
  not (_12295_, _12290_);
  or (_12296_, _12295_, _10963_);
  and (_12297_, _12296_, _12294_);
  and (_12298_, _10967_, _03105_);
  and (_12299_, _12298_, _10978_);
  or (_38680_, _12299_, _12297_);
  or (_12300_, _12295_, _11168_);
  or (_12301_, _12290_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_12302_, _12301_, _12293_);
  and (_12303_, _12302_, _12300_);
  and (_12304_, _12298_, _11176_);
  or (_38681_, _12304_, _12303_);
  or (_12305_, _12290_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_12306_, _12305_, _12293_);
  or (_12307_, _12295_, _11370_);
  and (_12309_, _12307_, _12306_);
  and (_12310_, _12298_, _11378_);
  or (_38682_, _12310_, _12309_);
  or (_12312_, _12295_, _11570_);
  or (_12314_, _12290_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_12315_, _12314_, _12293_);
  and (_12317_, _12315_, _12312_);
  and (_12318_, _12298_, _12221_);
  or (_38683_, _12318_, _12317_);
  or (_12320_, _12295_, _11774_);
  or (_12322_, _12290_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_12323_, _12322_, _12293_);
  and (_12325_, _12323_, _12320_);
  and (_12326_, _12298_, _11782_);
  or (_38684_, _12326_, _12325_);
  or (_12328_, _12290_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_12330_, _12328_, _12293_);
  or (_12331_, _12295_, _11977_);
  and (_12333_, _12331_, _12330_);
  and (_12334_, _12298_, _11986_);
  or (_38685_, _12334_, _12333_);
  or (_12336_, _12290_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_12338_, _12336_, _12293_);
  or (_12339_, _12295_, _12181_);
  and (_12341_, _12339_, _12338_);
  and (_12342_, _12298_, _12189_);
  or (_38686_, _12342_, _12341_);
  or (_12343_, _12290_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_12344_, _12343_, _12293_);
  or (_12345_, _12295_, _05378_);
  and (_12346_, _12345_, _12344_);
  and (_12347_, _12298_, _05431_);
  or (_38687_, _12347_, _12346_);
  not (_12348_, _05386_);
  and (_12349_, _05391_, _12348_);
  and (_12350_, _12349_, _03106_);
  not (_12351_, _12350_);
  or (_12352_, _12351_, _10978_);
  and (_12353_, _03743_, _03555_);
  and (_12354_, _12353_, _10782_);
  and (_12355_, _12354_, _10963_);
  nor (_12356_, _12354_, _02961_);
  or (_12357_, _12356_, _12350_);
  or (_12358_, _12357_, _12355_);
  and (_38692_, _12358_, _12352_);
  and (_12359_, _12350_, _11176_);
  not (_12360_, _12354_);
  or (_12361_, _12360_, _11168_);
  or (_12362_, _12354_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_12363_, _12362_, _12351_);
  and (_12364_, _12363_, _12361_);
  or (_38693_, _12364_, _12359_);
  and (_12365_, _12350_, _11378_);
  or (_12366_, _12360_, _11370_);
  or (_12367_, _12354_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_12368_, _12367_, _12351_);
  and (_12369_, _12368_, _12366_);
  or (_38694_, _12369_, _12365_);
  and (_12370_, _12350_, _12221_);
  or (_12371_, _12360_, _11570_);
  or (_12372_, _12354_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_12373_, _12372_, _12351_);
  and (_12374_, _12373_, _12371_);
  or (_38695_, _12374_, _12370_);
  or (_12375_, _12360_, _11774_);
  or (_12376_, _12354_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_12377_, _12376_, _12351_);
  and (_12378_, _12377_, _12375_);
  and (_12379_, _12350_, _11782_);
  or (_38696_, _12379_, _12378_);
  and (_12380_, _12350_, _11986_);
  or (_12381_, _12360_, _11977_);
  or (_12383_, _12354_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_12385_, _12383_, _12351_);
  and (_12386_, _12385_, _12381_);
  or (_38698_, _12386_, _12380_);
  and (_12388_, _12350_, _12189_);
  or (_12390_, _12360_, _12181_);
  or (_12391_, _12354_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_12393_, _12391_, _12351_);
  and (_12394_, _12393_, _12390_);
  or (_38699_, _12394_, _12388_);
  and (_12396_, _12350_, _05431_);
  or (_12398_, _12360_, _05378_);
  or (_12399_, _12354_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_12401_, _12399_, _12351_);
  and (_12402_, _12401_, _12398_);
  or (_38700_, _12402_, _12396_);
  and (_12404_, _12353_, _12196_);
  not (_12406_, _12404_);
  or (_12407_, _12406_, _10963_);
  and (_12409_, _12349_, _03437_);
  not (_12410_, _12409_);
  or (_12412_, _12404_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_12413_, _12412_, _12410_);
  and (_12414_, _12413_, _12407_);
  and (_12415_, _12409_, _10978_);
  or (_38703_, _12415_, _12414_);
  or (_12416_, _12406_, _11168_);
  or (_12417_, _12404_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_12418_, _12417_, _12410_);
  and (_12419_, _12418_, _12416_);
  and (_12420_, _12409_, _11176_);
  or (_38704_, _12420_, _12419_);
  or (_12421_, _12406_, _11370_);
  or (_12422_, _12404_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_12423_, _12422_, _12410_);
  and (_12424_, _12423_, _12421_);
  and (_12425_, _12409_, _11378_);
  or (_38705_, _12425_, _12424_);
  or (_12426_, _12406_, _11570_);
  or (_12427_, _12404_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_12428_, _12427_, _12410_);
  and (_12429_, _12428_, _12426_);
  and (_12430_, _12409_, _12221_);
  or (_38706_, _12430_, _12429_);
  or (_12431_, _12406_, _11774_);
  or (_12432_, _12404_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_12433_, _12432_, _12410_);
  and (_12434_, _12433_, _12431_);
  and (_12435_, _12409_, _11782_);
  or (_38708_, _12435_, _12434_);
  or (_12436_, _12406_, _11977_);
  or (_12437_, _12404_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_12438_, _12437_, _12410_);
  and (_12439_, _12438_, _12436_);
  and (_12440_, _12409_, _11986_);
  or (_38709_, _12440_, _12439_);
  or (_12441_, _12406_, _12181_);
  or (_12442_, _12404_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_12443_, _12442_, _12410_);
  and (_12444_, _12443_, _12441_);
  and (_12445_, _12409_, _12189_);
  or (_38710_, _12445_, _12444_);
  or (_12446_, _12406_, _05378_);
  or (_12447_, _12404_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_12448_, _12447_, _12410_);
  and (_12449_, _12448_, _12446_);
  and (_12450_, _12409_, _05431_);
  or (_38711_, _12450_, _12449_);
  and (_12451_, _12353_, _12244_);
  not (_12452_, _12451_);
  or (_12453_, _12452_, _10963_);
  and (_12454_, _12349_, _04551_);
  not (_12455_, _12454_);
  or (_12456_, _12451_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_12457_, _12456_, _12455_);
  and (_12458_, _12457_, _12453_);
  and (_12459_, _12454_, _10978_);
  or (_38714_, _12459_, _12458_);
  or (_12460_, _12452_, _11168_);
  or (_12461_, _12451_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_12462_, _12461_, _12455_);
  and (_12463_, _12462_, _12460_);
  and (_12464_, _12454_, _11176_);
  or (_38715_, _12464_, _12463_);
  or (_12465_, _12452_, _11370_);
  or (_12466_, _12451_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_12467_, _12466_, _12455_);
  and (_12468_, _12467_, _12465_);
  and (_12469_, _12454_, _11378_);
  or (_38716_, _12469_, _12468_);
  or (_12470_, _12452_, _11570_);
  or (_12471_, _12451_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_12472_, _12471_, _12455_);
  and (_12473_, _12472_, _12470_);
  and (_12474_, _12454_, _12221_);
  or (_38717_, _12474_, _12473_);
  or (_12475_, _12452_, _11774_);
  or (_12476_, _12451_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_12477_, _12476_, _12455_);
  and (_12478_, _12477_, _12475_);
  and (_12479_, _12454_, _11782_);
  or (_38719_, _12479_, _12478_);
  or (_12480_, _12452_, _11977_);
  or (_12481_, _12451_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_12482_, _12481_, _12455_);
  and (_12483_, _12482_, _12480_);
  and (_12484_, _12454_, _11986_);
  or (_38720_, _12484_, _12483_);
  or (_12485_, _12452_, _12181_);
  or (_12486_, _12451_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_12487_, _12486_, _12455_);
  and (_12488_, _12487_, _12485_);
  and (_12489_, _12454_, _12189_);
  or (_38721_, _12489_, _12488_);
  or (_12490_, _12452_, _05378_);
  or (_12491_, _12451_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_12492_, _12491_, _12455_);
  and (_12493_, _12492_, _12490_);
  and (_12494_, _12454_, _05431_);
  or (_38722_, _12494_, _12493_);
  and (_12495_, _12349_, _03105_);
  not (_12496_, _12495_);
  or (_12497_, _12496_, _10978_);
  and (_12498_, _12353_, _03387_);
  and (_12499_, _12498_, _10963_);
  nor (_12500_, _12498_, _02955_);
  or (_12501_, _12500_, _12495_);
  or (_12502_, _12501_, _12499_);
  and (_38726_, _12502_, _12497_);
  or (_12503_, _12498_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_12504_, _12503_, _12496_);
  not (_12505_, _12498_);
  or (_12506_, _12505_, _11168_);
  and (_12507_, _12506_, _12504_);
  and (_12508_, _12495_, _11176_);
  or (_38727_, _12508_, _12507_);
  or (_12509_, _12498_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_12510_, _12509_, _12496_);
  or (_12511_, _12505_, _11370_);
  and (_12512_, _12511_, _12510_);
  and (_12513_, _12495_, _11378_);
  or (_38728_, _12513_, _12512_);
  or (_12514_, _12498_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_12515_, _12514_, _12496_);
  or (_12516_, _12505_, _11570_);
  and (_12517_, _12516_, _12515_);
  and (_12518_, _12495_, _12221_);
  or (_38730_, _12518_, _12517_);
  or (_12519_, _12498_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_12520_, _12519_, _12496_);
  or (_12521_, _12505_, _11774_);
  and (_12522_, _12521_, _12520_);
  and (_12523_, _12495_, _11782_);
  or (_38731_, _12523_, _12522_);
  or (_12524_, _12498_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_12525_, _12524_, _12496_);
  or (_12526_, _12505_, _11977_);
  and (_12527_, _12526_, _12525_);
  and (_12528_, _12495_, _11986_);
  or (_38732_, _12528_, _12527_);
  or (_12529_, _12498_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_12530_, _12529_, _12496_);
  or (_12531_, _12505_, _12181_);
  and (_12532_, _12531_, _12530_);
  and (_12533_, _12495_, _12189_);
  or (_38733_, _12533_, _12532_);
  or (_12534_, _12498_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_12535_, _12534_, _12496_);
  or (_12536_, _12505_, _05378_);
  and (_12537_, _12536_, _12535_);
  and (_12538_, _12495_, _05431_);
  or (_38734_, _12538_, _12537_);
  and (_12539_, _10966_, _05384_);
  not (_12540_, _12539_);
  or (_12541_, _12540_, _10978_);
  and (_12542_, _10783_, _03742_);
  and (_12543_, _12542_, _10782_);
  and (_12544_, _12543_, _10963_);
  nor (_12545_, _12543_, _02978_);
  or (_12546_, _12545_, _12539_);
  or (_12547_, _12546_, _12544_);
  and (_38738_, _12547_, _12541_);
  not (_12548_, _12543_);
  or (_12549_, _12548_, _11168_);
  or (_12550_, _12543_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_12551_, _12550_, _12540_);
  and (_12552_, _12551_, _12549_);
  and (_12553_, _12539_, _11176_);
  or (_38739_, _12553_, _12552_);
  or (_12554_, _12548_, _11370_);
  or (_12555_, _12543_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_12556_, _12555_, _12540_);
  and (_12557_, _12556_, _12554_);
  and (_12558_, _12539_, _11378_);
  or (_38740_, _12558_, _12557_);
  or (_12559_, _12548_, _11570_);
  or (_12560_, _12543_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_12561_, _12560_, _12540_);
  and (_12562_, _12561_, _12559_);
  and (_12563_, _12539_, _12221_);
  or (_38741_, _12563_, _12562_);
  or (_12564_, _12548_, _11774_);
  or (_12565_, _12543_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_12566_, _12565_, _12540_);
  and (_12567_, _12566_, _12564_);
  and (_12568_, _12539_, _11782_);
  or (_38742_, _12568_, _12567_);
  or (_12569_, _12548_, _11977_);
  or (_12570_, _12543_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_12571_, _12570_, _12540_);
  and (_12572_, _12571_, _12569_);
  and (_12573_, _12539_, _11986_);
  or (_38744_, _12573_, _12572_);
  or (_12574_, _12548_, _12181_);
  or (_12575_, _12543_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_12576_, _12575_, _12540_);
  and (_12577_, _12576_, _12574_);
  and (_12578_, _12539_, _12189_);
  or (_38745_, _12578_, _12577_);
  or (_12579_, _12548_, _05378_);
  or (_12580_, _12543_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_12581_, _12580_, _12540_);
  and (_12582_, _12581_, _12579_);
  and (_12583_, _12539_, _05431_);
  or (_38746_, _12583_, _12582_);
  and (_12584_, _12542_, _12196_);
  not (_12585_, _12584_);
  or (_12586_, _12585_, _10963_);
  not (_12587_, _05388_);
  and (_12588_, _10966_, _12587_);
  and (_12589_, _12588_, _03437_);
  not (_12590_, _12589_);
  or (_12591_, _12584_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_12592_, _12591_, _12590_);
  and (_12593_, _12592_, _12586_);
  and (_12594_, _12589_, _10978_);
  or (_38749_, _12594_, _12593_);
  or (_12595_, _12585_, _11168_);
  or (_12596_, _12584_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_12597_, _12596_, _12590_);
  and (_12598_, _12597_, _12595_);
  and (_12599_, _12589_, _11176_);
  or (_38750_, _12599_, _12598_);
  or (_12600_, _12585_, _11370_);
  or (_12601_, _12584_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_12602_, _12601_, _12590_);
  and (_12603_, _12602_, _12600_);
  and (_12604_, _12589_, _11378_);
  or (_38751_, _12604_, _12603_);
  or (_12605_, _12585_, _11570_);
  or (_12606_, _12584_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_12607_, _12606_, _12590_);
  and (_12608_, _12607_, _12605_);
  and (_12609_, _12589_, _12221_);
  or (_38752_, _12609_, _12608_);
  or (_12610_, _12585_, _11774_);
  or (_12611_, _12584_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_12612_, _12611_, _12590_);
  and (_12613_, _12612_, _12610_);
  and (_12614_, _12589_, _11782_);
  or (_38754_, _12614_, _12613_);
  or (_12615_, _12585_, _11977_);
  or (_12616_, _12584_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_12617_, _12616_, _12590_);
  and (_12618_, _12617_, _12615_);
  and (_12619_, _12589_, _11986_);
  or (_38755_, _12619_, _12618_);
  or (_12620_, _12585_, _12181_);
  or (_12621_, _12584_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_12622_, _12621_, _12590_);
  and (_12623_, _12622_, _12620_);
  and (_12624_, _12589_, _12189_);
  or (_38756_, _12624_, _12623_);
  or (_12625_, _12585_, _05378_);
  or (_12626_, _12584_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_12627_, _12626_, _12590_);
  and (_12628_, _12627_, _12625_);
  and (_12629_, _12589_, _05431_);
  or (_38757_, _12629_, _12628_);
  and (_12630_, _12542_, _12244_);
  not (_12631_, _12630_);
  or (_12632_, _12631_, _10963_);
  and (_12633_, _12588_, _04551_);
  not (_12634_, _12633_);
  or (_12635_, _12630_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_12636_, _12635_, _12634_);
  and (_12637_, _12636_, _12632_);
  and (_12638_, _12633_, _10978_);
  or (_38761_, _12638_, _12637_);
  or (_12639_, _12631_, _11168_);
  or (_12640_, _12630_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_12641_, _12640_, _12634_);
  and (_12642_, _12641_, _12639_);
  and (_12643_, _12633_, _11176_);
  or (_38762_, _12643_, _12642_);
  or (_12644_, _12631_, _11370_);
  or (_12645_, _12630_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_12646_, _12645_, _12634_);
  and (_12647_, _12646_, _12644_);
  and (_12648_, _12633_, _11378_);
  or (_38763_, _12648_, _12647_);
  or (_12649_, _12631_, _11570_);
  or (_12650_, _12630_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_12651_, _12650_, _12634_);
  and (_12652_, _12651_, _12649_);
  and (_12653_, _12633_, _12221_);
  or (_38764_, _12653_, _12652_);
  or (_12654_, _12631_, _11774_);
  or (_12655_, _12630_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_12656_, _12655_, _12634_);
  and (_12657_, _12656_, _12654_);
  and (_12658_, _12633_, _11782_);
  or (_38765_, _12658_, _12657_);
  or (_12659_, _12631_, _11977_);
  or (_12660_, _12630_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_12661_, _12660_, _12634_);
  and (_12662_, _12661_, _12659_);
  and (_12663_, _12633_, _11986_);
  or (_38766_, _12663_, _12662_);
  or (_12664_, _12631_, _12181_);
  or (_12665_, _12630_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_12666_, _12665_, _12634_);
  and (_12667_, _12666_, _12664_);
  and (_12668_, _12633_, _12189_);
  or (_38767_, _12668_, _12667_);
  or (_12669_, _12631_, _05378_);
  or (_12670_, _12630_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_12671_, _12670_, _12634_);
  and (_12672_, _12671_, _12669_);
  and (_12673_, _12633_, _05431_);
  or (_38768_, _12673_, _12672_);
  nor (_12674_, _05388_, _05382_);
  nand (_12675_, _12674_, _10966_);
  nor (_12676_, _12675_, _10978_);
  and (_12677_, _12542_, _03387_);
  nand (_12678_, _12677_, _10963_);
  or (_12679_, _12677_, _02972_);
  and (_12680_, _12679_, _12675_);
  and (_12681_, _12680_, _12678_);
  nor (_38772_, _12681_, _12676_);
  and (_12682_, _12588_, _03105_);
  not (_12683_, _12682_);
  or (_12684_, _12677_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_12685_, _12684_, _12683_);
  not (_12686_, _12677_);
  or (_12687_, _12686_, _11168_);
  and (_12688_, _12687_, _12685_);
  and (_12689_, _12682_, _11176_);
  or (_38773_, _12689_, _12688_);
  or (_12690_, _12677_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_12691_, _12690_, _12683_);
  or (_12692_, _12686_, _11370_);
  and (_12693_, _12692_, _12691_);
  and (_12694_, _12682_, _11378_);
  or (_38774_, _12694_, _12693_);
  or (_12695_, _12677_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_12696_, _12695_, _12683_);
  or (_12697_, _12686_, _11570_);
  and (_12698_, _12697_, _12696_);
  and (_12699_, _12682_, _12221_);
  or (_38776_, _12699_, _12698_);
  or (_12700_, _12686_, _11774_);
  or (_12701_, _12677_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_12702_, _12701_, _12683_);
  and (_12703_, _12702_, _12700_);
  and (_12704_, _12682_, _11782_);
  or (_38777_, _12704_, _12703_);
  or (_12705_, _12686_, _11977_);
  or (_12706_, _12677_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_12707_, _12706_, _12683_);
  and (_12708_, _12707_, _12705_);
  and (_12709_, _12682_, _11986_);
  or (_38778_, _12709_, _12708_);
  or (_12710_, _12677_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_12711_, _12710_, _12683_);
  or (_12712_, _12686_, _12181_);
  and (_12713_, _12712_, _12711_);
  and (_12714_, _12682_, _12189_);
  or (_38779_, _12714_, _12713_);
  and (_12715_, _12677_, _05378_);
  or (_12716_, _12677_, _03772_);
  nand (_12717_, _12716_, _12675_);
  or (_12718_, _12717_, _12715_);
  or (_12719_, _12683_, _05431_);
  and (_38780_, _12719_, _12718_);
  not (_12720_, _03742_);
  and (_12721_, _10783_, _12720_);
  and (_12722_, _10782_, _12721_);
  not (_12723_, _12722_);
  or (_12724_, _12723_, _10963_);
  and (_12725_, _10966_, _05388_);
  and (_12726_, _12725_, _03106_);
  not (_12727_, _12726_);
  or (_12728_, _12722_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_12729_, _12728_, _12727_);
  and (_12730_, _12729_, _12724_);
  and (_12731_, _12726_, _10978_);
  or (_38783_, _12731_, _12730_);
  and (_12732_, _10782_, _03745_);
  or (_12733_, _12732_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_12734_, _12733_, _12727_);
  not (_12735_, _12732_);
  or (_12736_, _12735_, _11168_);
  and (_12737_, _12736_, _12734_);
  and (_12738_, _12726_, _11176_);
  or (_38784_, _12738_, _12737_);
  or (_12739_, _12732_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_12740_, _12739_, _12727_);
  or (_12741_, _12735_, _11370_);
  and (_12742_, _12741_, _12740_);
  and (_12743_, _12726_, _11378_);
  or (_38786_, _12743_, _12742_);
  or (_12744_, _12732_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_12745_, _12744_, _12727_);
  or (_12746_, _12735_, _11570_);
  and (_12747_, _12746_, _12745_);
  and (_12748_, _12726_, _12221_);
  or (_38787_, _12748_, _12747_);
  or (_12749_, _12732_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_12750_, _12749_, _12727_);
  or (_12751_, _12735_, _11774_);
  and (_12752_, _12751_, _12750_);
  and (_12753_, _12726_, _11782_);
  or (_38788_, _12753_, _12752_);
  or (_12754_, _12732_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_12755_, _12754_, _12727_);
  or (_12756_, _12735_, _11977_);
  and (_12757_, _12756_, _12755_);
  and (_12758_, _12726_, _11986_);
  or (_38789_, _12758_, _12757_);
  or (_12759_, _12732_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_12760_, _12759_, _12727_);
  or (_12761_, _12735_, _12181_);
  and (_12762_, _12761_, _12760_);
  and (_12763_, _12726_, _12189_);
  or (_38790_, _12763_, _12762_);
  nor (_12764_, _12722_, \oc8051_golden_model_1.IRAM[12] [7]);
  nor (_12765_, _12723_, _05378_);
  or (_12766_, _12765_, _12764_);
  nand (_12767_, _12766_, _12727_);
  or (_12768_, _12727_, _05431_);
  and (_38792_, _12768_, _12767_);
  nand (_12769_, _12196_, _12721_);
  or (_12770_, _12769_, _10963_);
  and (_12771_, _12725_, _03437_);
  not (_12772_, _12771_);
  nand (_12773_, _12769_, _02994_);
  and (_12774_, _12773_, _12772_);
  and (_12775_, _12774_, _12770_);
  and (_12776_, _12771_, _10978_);
  or (_38795_, _12776_, _12775_);
  or (_12777_, _12769_, _11168_);
  nand (_12778_, _12769_, _03152_);
  and (_12779_, _12778_, _12772_);
  and (_12780_, _12779_, _12777_);
  and (_12781_, _12771_, _11176_);
  or (_38797_, _12781_, _12780_);
  nand (_12782_, _12769_, _03616_);
  and (_12783_, _12782_, _12772_);
  or (_12784_, _12769_, _11370_);
  and (_12785_, _12784_, _12783_);
  and (_12786_, _12771_, _11378_);
  or (_38798_, _12786_, _12785_);
  nand (_12787_, _12769_, _03426_);
  and (_12788_, _12787_, _12772_);
  or (_12789_, _12769_, _11570_);
  and (_12790_, _12789_, _12788_);
  and (_12791_, _12771_, _12221_);
  or (_38799_, _12791_, _12790_);
  nand (_12792_, _12769_, _04364_);
  and (_12793_, _12792_, _12772_);
  or (_12794_, _12769_, _11774_);
  and (_12795_, _12794_, _12793_);
  and (_12796_, _12771_, _11782_);
  or (_38800_, _12796_, _12795_);
  or (_12797_, _12769_, _11977_);
  nand (_12798_, _12769_, _04049_);
  and (_12799_, _12798_, _12772_);
  and (_12800_, _12799_, _12797_);
  and (_12801_, _12771_, _11986_);
  or (_38801_, _12801_, _12800_);
  or (_12802_, _12769_, _12181_);
  nand (_12803_, _12769_, _03956_);
  and (_12804_, _12803_, _12772_);
  and (_12805_, _12804_, _12802_);
  and (_12806_, _12771_, _12189_);
  or (_38802_, _12806_, _12805_);
  nand (_12807_, _12769_, _03788_);
  and (_12808_, _12807_, _12772_);
  or (_12809_, _12769_, _05378_);
  and (_12810_, _12809_, _12808_);
  and (_12811_, _12771_, _05431_);
  or (_38803_, _12811_, _12810_);
  nand (_12812_, _12244_, _12721_);
  nor (_12813_, _12812_, _10963_);
  and (_12814_, _12725_, _04551_);
  and (_12815_, _12812_, _02988_);
  or (_12816_, _12815_, _12814_);
  nor (_12817_, _12816_, _12813_);
  and (_12818_, _12814_, _10978_);
  or (_38806_, _12818_, _12817_);
  not (_12819_, _12814_);
  and (_12820_, _12244_, _03745_);
  or (_12821_, _12820_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_12822_, _12821_, _12819_);
  not (_12823_, _12820_);
  or (_12824_, _12823_, _11168_);
  and (_12825_, _12824_, _12822_);
  and (_12826_, _12814_, _11176_);
  or (_38808_, _12826_, _12825_);
  or (_12827_, _12820_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_12828_, _12827_, _12819_);
  or (_12829_, _12823_, _11370_);
  and (_12830_, _12829_, _12828_);
  and (_12831_, _12814_, _11378_);
  or (_38809_, _12831_, _12830_);
  or (_12832_, _12820_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_12833_, _12832_, _12819_);
  or (_12834_, _12823_, _11570_);
  and (_12835_, _12834_, _12833_);
  and (_12836_, _12814_, _12221_);
  or (_38810_, _12836_, _12835_);
  or (_12837_, _12820_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_12838_, _12837_, _12819_);
  or (_12839_, _12823_, _11774_);
  and (_12840_, _12839_, _12838_);
  and (_12841_, _12814_, _11782_);
  or (_38811_, _12841_, _12840_);
  or (_12842_, _12820_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_12843_, _12842_, _12819_);
  or (_12844_, _12823_, _11977_);
  and (_12845_, _12844_, _12843_);
  and (_12846_, _12814_, _11986_);
  or (_38812_, _12846_, _12845_);
  or (_12847_, _12820_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_12848_, _12847_, _12819_);
  or (_12849_, _12823_, _12181_);
  and (_12850_, _12849_, _12848_);
  and (_12851_, _12814_, _12189_);
  or (_38814_, _12851_, _12850_);
  or (_12852_, _12820_, \oc8051_golden_model_1.IRAM[14] [7]);
  and (_12853_, _12852_, _12819_);
  or (_12854_, _12823_, _05378_);
  and (_12855_, _12854_, _12853_);
  and (_12856_, _12814_, _05431_);
  or (_38815_, _12856_, _12855_);
  nor (_12857_, _03746_, _02986_);
  and (_12858_, _10963_, _03746_);
  or (_12859_, _12858_, _12857_);
  and (_12860_, _12859_, _05393_);
  and (_12861_, _12725_, _03105_);
  and (_12862_, _10978_, _12861_);
  or (_38817_, _12862_, _12860_);
  or (_12863_, _11168_, _03747_);
  not (_12864_, _12861_);
  or (_12865_, _03746_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_12866_, _12865_, _12864_);
  and (_12867_, _12866_, _12863_);
  and (_12868_, _11176_, _12861_);
  or (_38819_, _12868_, _12867_);
  or (_12869_, _11370_, _03747_);
  or (_12870_, _03746_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_12871_, _12870_, _12864_);
  and (_12872_, _12871_, _12869_);
  and (_12873_, _11378_, _12861_);
  or (_38820_, _12873_, _12872_);
  or (_12874_, _03746_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_12875_, _12874_, _12864_);
  or (_12876_, _11570_, _03747_);
  and (_12877_, _12876_, _12875_);
  and (_12878_, _12221_, _12861_);
  or (_38821_, _12878_, _12877_);
  or (_12879_, _03746_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_12880_, _12879_, _12864_);
  or (_12881_, _11774_, _03747_);
  and (_12882_, _12881_, _12880_);
  and (_12883_, _11782_, _12861_);
  or (_38822_, _12883_, _12882_);
  or (_12884_, _03746_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_12885_, _12884_, _12864_);
  or (_12886_, _11977_, _03747_);
  and (_12887_, _12886_, _12885_);
  and (_12888_, _11986_, _12861_);
  or (_38823_, _12888_, _12887_);
  or (_12889_, _03746_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_12890_, _12889_, _12864_);
  or (_12891_, _12181_, _03747_);
  and (_12892_, _12891_, _12890_);
  and (_12893_, _12189_, _12861_);
  or (_38825_, _12893_, _12892_);
  nor (_12894_, _39632_, _06214_);
  nor (_12895_, _03847_, _06214_);
  and (_12896_, _10792_, _03847_);
  or (_12897_, _12896_, _12895_);
  and (_12898_, _12897_, _02331_);
  and (_12899_, _03847_, _03002_);
  or (_12900_, _12899_, _12895_);
  or (_12901_, _12900_, _05444_);
  nor (_12902_, _04257_, _05439_);
  or (_12903_, _12902_, _12895_);
  or (_12904_, _12903_, _03006_);
  and (_12905_, _03847_, \oc8051_golden_model_1.ACC [0]);
  or (_12906_, _12905_, _12895_);
  and (_12907_, _12906_, _02062_);
  nor (_12908_, _02062_, _06214_);
  or (_12909_, _12908_, _02158_);
  or (_12910_, _12909_, _12907_);
  and (_12911_, _12910_, _02058_);
  and (_12912_, _12911_, _12904_);
  and (_12913_, _10814_, _04478_);
  nor (_12914_, _04478_, _06214_);
  or (_12915_, _12914_, _12913_);
  and (_12916_, _12915_, _02057_);
  or (_12917_, _12916_, _12912_);
  and (_12918_, _12917_, _02519_);
  and (_12919_, _12900_, _02155_);
  or (_12920_, _12919_, _02153_);
  or (_12921_, _12920_, _12918_);
  or (_12922_, _12906_, _02549_);
  and (_12923_, _12922_, _02054_);
  and (_12924_, _12923_, _12921_);
  and (_12925_, _12895_, _02053_);
  or (_12926_, _12925_, _02046_);
  or (_12927_, _12926_, _12924_);
  or (_12928_, _12903_, _02047_);
  and (_12929_, _12928_, _12927_);
  or (_12930_, _12929_, _05474_);
  nor (_12931_, _06148_, _06146_);
  nor (_12932_, _12931_, _06149_);
  or (_12933_, _12932_, _06181_);
  and (_12934_, _12933_, _02043_);
  and (_12935_, _12934_, _12930_);
  nor (_12936_, _10798_, _06189_);
  or (_12937_, _12936_, _12914_);
  and (_12938_, _12937_, _02042_);
  or (_12939_, _12938_, _06188_);
  or (_12940_, _12939_, _12935_);
  and (_12941_, _12940_, _12901_);
  or (_12942_, _12941_, _02031_);
  and (_12943_, _05120_, _03847_);
  or (_12944_, _12895_, _02032_);
  or (_12945_, _12944_, _12943_);
  and (_12946_, _12945_, _12942_);
  or (_12947_, _12946_, _01765_);
  nor (_12948_, _10898_, _05439_);
  or (_12949_, _12895_, _02037_);
  or (_12950_, _12949_, _12948_);
  and (_12951_, _12950_, _06560_);
  and (_12952_, _12951_, _12947_);
  nand (_12953_, _06558_, _01887_);
  nor (_12954_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_12955_, _12954_, _06127_);
  or (_12956_, _06558_, _12955_);
  and (_12957_, _12956_, _06202_);
  and (_12958_, _12957_, _12953_);
  or (_12959_, _12958_, _07629_);
  or (_12960_, _12959_, _12952_);
  and (_12961_, _10914_, _03847_);
  or (_12962_, _12895_, _03059_);
  or (_12963_, _12962_, _12961_);
  and (_12964_, _03847_, _04837_);
  or (_12965_, _12964_, _12895_);
  or (_12966_, _12965_, _01995_);
  and (_12967_, _12966_, _03061_);
  and (_12968_, _12967_, _12963_);
  and (_12969_, _12968_, _12960_);
  or (_12970_, _12969_, _12898_);
  and (_12971_, _12970_, _02208_);
  nand (_12972_, _12965_, _02206_);
  nor (_12973_, _12972_, _12902_);
  or (_12974_, _12973_, _12971_);
  and (_12975_, _12974_, _03065_);
  or (_12976_, _12895_, _04257_);
  and (_12977_, _12906_, _02342_);
  and (_12978_, _12977_, _12976_);
  or (_12979_, _12978_, _02202_);
  or (_12980_, _12979_, _12975_);
  nor (_12981_, _10913_, _05439_);
  or (_12982_, _12895_, _04953_);
  or (_12983_, _12982_, _12981_);
  and (_12984_, _12983_, _04958_);
  and (_12985_, _12984_, _12980_);
  nor (_12986_, _10789_, _05439_);
  or (_12987_, _12986_, _12895_);
  and (_12988_, _12987_, _02334_);
  or (_12989_, _12988_, _02366_);
  or (_12990_, _12989_, _12985_);
  or (_12991_, _12903_, _02778_);
  and (_12992_, _12991_, _01698_);
  and (_12993_, _12992_, _12990_);
  and (_12994_, _12895_, _01697_);
  or (_12995_, _12994_, _02081_);
  or (_12996_, _12995_, _12993_);
  or (_12997_, _12903_, _02082_);
  and (_12998_, _12997_, _39632_);
  and (_12999_, _12998_, _12996_);
  or (_13000_, _12999_, _12894_);
  and (_41617_, _13000_, _39026_);
  nor (_13001_, _39632_, _06208_);
  nor (_13002_, _04478_, _06208_);
  and (_13003_, _11005_, _04478_);
  or (_13004_, _13003_, _13002_);
  or (_13005_, _13002_, _11020_);
  and (_13006_, _13005_, _13004_);
  or (_13007_, _13006_, _02047_);
  or (_13008_, _03847_, \oc8051_golden_model_1.B [1]);
  and (_13009_, _11001_, _03847_);
  not (_13010_, _13009_);
  and (_13011_, _13010_, _13008_);
  or (_13012_, _13011_, _03006_);
  nand (_13013_, _03847_, _01804_);
  and (_13014_, _13013_, _13008_);
  and (_13015_, _13014_, _02062_);
  nor (_13016_, _02062_, _06208_);
  or (_13017_, _13016_, _02158_);
  or (_13018_, _13017_, _13015_);
  and (_13019_, _13018_, _02058_);
  and (_13020_, _13019_, _13012_);
  and (_13021_, _13004_, _02057_);
  or (_13022_, _13021_, _02155_);
  or (_13023_, _13022_, _13020_);
  nor (_13024_, _03847_, _06208_);
  nor (_13025_, _05439_, _03161_);
  or (_13026_, _13025_, _13024_);
  or (_13027_, _13026_, _02519_);
  and (_13028_, _13027_, _13023_);
  or (_13029_, _13028_, _02153_);
  or (_13030_, _13014_, _02549_);
  and (_13031_, _13030_, _02054_);
  and (_13032_, _13031_, _13029_);
  and (_13033_, _10992_, _04478_);
  or (_13034_, _13033_, _13002_);
  and (_13035_, _13034_, _02053_);
  or (_13036_, _13035_, _02046_);
  or (_13037_, _13036_, _13032_);
  and (_13038_, _13037_, _13007_);
  or (_13039_, _13038_, _05474_);
  nor (_13040_, _06151_, _06094_);
  nor (_13041_, _13040_, _06152_);
  or (_13042_, _13041_, _06181_);
  and (_13043_, _13042_, _02043_);
  and (_13044_, _13043_, _13039_);
  nor (_13045_, _11038_, _06189_);
  or (_13046_, _13045_, _13002_);
  and (_13047_, _13046_, _02042_);
  or (_13048_, _13047_, _06188_);
  or (_13049_, _13048_, _13044_);
  or (_13050_, _13026_, _05444_);
  and (_13051_, _13050_, _13049_);
  or (_13052_, _13051_, _02031_);
  and (_13053_, _05075_, _03847_);
  or (_13054_, _13024_, _02032_);
  or (_13055_, _13054_, _13053_);
  and (_13056_, _13055_, _02037_);
  and (_13057_, _13056_, _13052_);
  nand (_13058_, _11096_, _03847_);
  and (_13059_, _13008_, _01765_);
  and (_13060_, _13059_, _13058_);
  or (_13061_, _13060_, _06202_);
  or (_13062_, _13061_, _13057_);
  and (_13063_, _06558_, _06524_);
  nor (_13064_, _06553_, _06552_);
  or (_13065_, _13064_, _06554_);
  nor (_13066_, _13065_, _06558_);
  or (_13067_, _13066_, _13063_);
  or (_13068_, _13067_, _06560_);
  and (_13069_, _13068_, _01995_);
  and (_13070_, _13069_, _13062_);
  nand (_13071_, _03847_, _02893_);
  and (_13072_, _13008_, _01994_);
  and (_13073_, _13072_, _13071_);
  or (_13074_, _13073_, _13070_);
  and (_13075_, _13074_, _03059_);
  or (_13076_, _10989_, _05439_);
  and (_13077_, _13008_, _02210_);
  and (_13078_, _13077_, _13076_);
  or (_13079_, _13078_, _13075_);
  and (_13080_, _13079_, _03061_);
  or (_13081_, _11113_, _05439_);
  and (_13082_, _13008_, _02331_);
  and (_13083_, _13082_, _13081_);
  or (_13084_, _13083_, _13080_);
  and (_13085_, _13084_, _02208_);
  or (_13086_, _10988_, _05439_);
  and (_13087_, _13008_, _02206_);
  and (_13088_, _13087_, _13086_);
  or (_13089_, _13088_, _13085_);
  and (_13090_, _13089_, _03065_);
  or (_13091_, _13024_, _04209_);
  and (_13092_, _13014_, _02342_);
  and (_13093_, _13092_, _13091_);
  or (_13094_, _13093_, _13090_);
  and (_13095_, _13094_, _02335_);
  or (_13096_, _13013_, _04209_);
  and (_13097_, _13008_, _02334_);
  and (_13098_, _13097_, _13096_);
  or (_13099_, _13098_, _02366_);
  or (_13100_, _13071_, _04209_);
  and (_13101_, _13008_, _02202_);
  and (_13102_, _13101_, _13100_);
  or (_13103_, _13102_, _13099_);
  or (_13104_, _13103_, _13095_);
  or (_13105_, _13011_, _02778_);
  and (_13106_, _13105_, _01698_);
  and (_13107_, _13106_, _13104_);
  and (_13108_, _13034_, _01697_);
  or (_13109_, _13108_, _02081_);
  or (_13110_, _13109_, _13107_);
  or (_13111_, _13024_, _02082_);
  or (_13112_, _13111_, _13009_);
  and (_13113_, _13112_, _39632_);
  and (_13114_, _13113_, _13110_);
  or (_13115_, _13114_, _13001_);
  and (_41618_, _13115_, _39026_);
  nor (_13116_, _39632_, _06222_);
  nor (_13117_, _03847_, _06222_);
  nor (_13118_, _05439_, _03624_);
  or (_13119_, _13118_, _13117_);
  or (_13120_, _13119_, _05444_);
  nor (_13121_, _04478_, _06222_);
  and (_13122_, _11194_, _04478_);
  or (_13123_, _13122_, _13121_);
  or (_13124_, _13121_, _11223_);
  and (_13125_, _13124_, _13123_);
  or (_13126_, _13125_, _02047_);
  nor (_13127_, _11199_, _05439_);
  or (_13128_, _13127_, _13117_);
  or (_13129_, _13128_, _03006_);
  and (_13130_, _03847_, \oc8051_golden_model_1.ACC [2]);
  or (_13131_, _13130_, _13117_);
  and (_13132_, _13131_, _02062_);
  nor (_13133_, _02062_, _06222_);
  or (_13134_, _13133_, _02158_);
  or (_13135_, _13134_, _13132_);
  and (_13136_, _13135_, _02058_);
  and (_13137_, _13136_, _13129_);
  and (_13138_, _13123_, _02057_);
  or (_13139_, _13138_, _02155_);
  or (_13140_, _13139_, _13137_);
  or (_13141_, _13119_, _02519_);
  and (_13142_, _13141_, _13140_);
  or (_13143_, _13142_, _02153_);
  or (_13144_, _13131_, _02549_);
  and (_13145_, _13144_, _02054_);
  and (_13146_, _13145_, _13143_);
  and (_13147_, _11192_, _04478_);
  or (_13148_, _13147_, _13121_);
  and (_13149_, _13148_, _02053_);
  or (_13150_, _13149_, _02046_);
  or (_13151_, _13150_, _13146_);
  and (_13152_, _13151_, _13126_);
  or (_13153_, _13152_, _05474_);
  nor (_13154_, _06154_, _06049_);
  nor (_13155_, _13154_, _06155_);
  or (_13156_, _13155_, _06181_);
  and (_13157_, _13156_, _02043_);
  and (_13158_, _13157_, _13153_);
  nor (_13159_, _11241_, _06189_);
  or (_13160_, _13159_, _13121_);
  and (_13161_, _13160_, _02042_);
  or (_13162_, _13161_, _06188_);
  or (_13163_, _13162_, _13158_);
  and (_13164_, _13163_, _13120_);
  or (_13165_, _13164_, _02031_);
  and (_13166_, _05211_, _03847_);
  or (_13167_, _13117_, _02032_);
  or (_13168_, _13167_, _13166_);
  and (_13169_, _13168_, _13165_);
  or (_13170_, _13169_, _01765_);
  nor (_13171_, _11298_, _05439_);
  or (_13172_, _13117_, _02037_);
  or (_13173_, _13172_, _13171_);
  and (_13174_, _13173_, _06560_);
  and (_13175_, _13174_, _13170_);
  not (_13176_, _06558_);
  or (_13177_, _13176_, _06514_);
  nor (_13178_, _06554_, _06525_);
  not (_13179_, _13178_);
  and (_13180_, _13179_, _06517_);
  nor (_13181_, _13179_, _06517_);
  nor (_13182_, _13181_, _13180_);
  or (_13183_, _13182_, _06558_);
  and (_13184_, _13183_, _06202_);
  and (_13185_, _13184_, _13177_);
  or (_13186_, _13185_, _07629_);
  or (_13187_, _13186_, _13175_);
  and (_13188_, _11189_, _03847_);
  or (_13189_, _13117_, _03059_);
  or (_13190_, _13189_, _13188_);
  and (_13191_, _03847_, _04866_);
  or (_13192_, _13191_, _13117_);
  or (_13193_, _13192_, _01995_);
  and (_13194_, _13193_, _03061_);
  and (_13195_, _13194_, _13190_);
  and (_13196_, _13195_, _13187_);
  and (_13197_, _11315_, _03847_);
  or (_13198_, _13197_, _13117_);
  and (_13199_, _13198_, _02331_);
  or (_13200_, _13199_, _13196_);
  and (_13201_, _13200_, _02208_);
  or (_13202_, _13117_, _04309_);
  and (_13203_, _13192_, _02206_);
  and (_13204_, _13203_, _13202_);
  or (_13205_, _13204_, _13201_);
  and (_13206_, _13205_, _03065_);
  and (_13207_, _13131_, _02342_);
  and (_13208_, _13207_, _13202_);
  or (_13209_, _13208_, _02202_);
  or (_13210_, _13209_, _13206_);
  nor (_13211_, _11187_, _05439_);
  or (_13212_, _13117_, _04953_);
  or (_13213_, _13212_, _13211_);
  and (_13214_, _13213_, _04958_);
  and (_13215_, _13214_, _13210_);
  nor (_13216_, _11314_, _05439_);
  or (_13217_, _13216_, _13117_);
  and (_13218_, _13217_, _02334_);
  or (_13219_, _13218_, _02366_);
  or (_13220_, _13219_, _13215_);
  or (_13221_, _13128_, _02778_);
  and (_13222_, _13221_, _01698_);
  and (_13223_, _13222_, _13220_);
  and (_13224_, _13148_, _01697_);
  or (_13225_, _13224_, _02081_);
  or (_13226_, _13225_, _13223_);
  and (_13227_, _11367_, _03847_);
  or (_13228_, _13117_, _02082_);
  or (_13229_, _13228_, _13227_);
  and (_13230_, _13229_, _39632_);
  and (_13231_, _13230_, _13226_);
  or (_13232_, _13231_, _13116_);
  and (_41619_, _13232_, _39026_);
  nor (_13233_, _39632_, _06223_);
  nor (_13234_, _03847_, _06223_);
  nor (_13235_, _05439_, _03434_);
  or (_13236_, _13235_, _13234_);
  or (_13237_, _13236_, _05444_);
  nor (_13238_, _04478_, _06223_);
  and (_13239_, _11398_, _04478_);
  or (_13240_, _13239_, _13238_);
  or (_13241_, _13238_, _11415_);
  and (_13242_, _13241_, _13240_);
  or (_13243_, _13242_, _02047_);
  nor (_13244_, _11394_, _05439_);
  or (_13245_, _13244_, _13234_);
  or (_13246_, _13245_, _03006_);
  and (_13247_, _03847_, \oc8051_golden_model_1.ACC [3]);
  or (_13248_, _13247_, _13234_);
  and (_13249_, _13248_, _02062_);
  nor (_13250_, _02062_, _06223_);
  or (_13251_, _13250_, _02158_);
  or (_13252_, _13251_, _13249_);
  and (_13253_, _13252_, _02058_);
  and (_13254_, _13253_, _13246_);
  and (_13255_, _13240_, _02057_);
  or (_13256_, _13255_, _02155_);
  or (_13257_, _13256_, _13254_);
  or (_13258_, _13236_, _02519_);
  and (_13259_, _13258_, _13257_);
  or (_13260_, _13259_, _02153_);
  or (_13261_, _13248_, _02549_);
  and (_13262_, _13261_, _02054_);
  and (_13263_, _13262_, _13260_);
  and (_13264_, _11408_, _04478_);
  or (_13265_, _13264_, _13238_);
  and (_13266_, _13265_, _02053_);
  or (_13267_, _13266_, _02046_);
  or (_13268_, _13267_, _13263_);
  and (_13269_, _13268_, _13243_);
  or (_13270_, _13269_, _05474_);
  nor (_13271_, _06157_, _05991_);
  nor (_13272_, _13271_, _06158_);
  or (_13273_, _13272_, _06181_);
  and (_13274_, _13273_, _02043_);
  and (_13275_, _13274_, _13270_);
  nor (_13276_, _11433_, _06189_);
  or (_13277_, _13276_, _13238_);
  and (_13278_, _13277_, _02042_);
  or (_13279_, _13278_, _06188_);
  or (_13280_, _13279_, _13275_);
  and (_13281_, _13280_, _13237_);
  or (_13282_, _13281_, _02031_);
  and (_13283_, _05166_, _03847_);
  or (_13284_, _13234_, _02032_);
  or (_13285_, _13284_, _13283_);
  and (_13286_, _13285_, _13282_);
  or (_13287_, _13286_, _01765_);
  nor (_13288_, _11490_, _05439_);
  or (_13289_, _13234_, _02037_);
  or (_13290_, _13289_, _13288_);
  and (_13291_, _13290_, _06560_);
  and (_13292_, _13291_, _13287_);
  nor (_13293_, _13180_, _06516_);
  nor (_13294_, _13293_, _06509_);
  and (_13295_, _13293_, _06509_);
  or (_13296_, _13295_, _13294_);
  or (_13297_, _13296_, _06558_);
  or (_13298_, _13176_, _06506_);
  and (_13299_, _13298_, _06202_);
  and (_13300_, _13299_, _13297_);
  or (_13301_, _13300_, _07629_);
  or (_13302_, _13301_, _13292_);
  and (_13303_, _11505_, _03847_);
  or (_13304_, _13234_, _03059_);
  or (_13305_, _13304_, _13303_);
  and (_13306_, _03847_, _04719_);
  or (_13307_, _13306_, _13234_);
  or (_13308_, _13307_, _01995_);
  and (_13309_, _13308_, _03061_);
  and (_13310_, _13309_, _13305_);
  and (_13311_, _13310_, _13302_);
  and (_13312_, _11511_, _03847_);
  or (_13313_, _13312_, _13234_);
  and (_13314_, _13313_, _02331_);
  or (_13315_, _13314_, _13311_);
  and (_13316_, _13315_, _02208_);
  or (_13317_, _13234_, _04153_);
  and (_13318_, _13307_, _02206_);
  and (_13319_, _13318_, _13317_);
  or (_13320_, _13319_, _13316_);
  and (_13321_, _13320_, _03065_);
  and (_13322_, _13248_, _02342_);
  and (_13323_, _13322_, _13317_);
  or (_13324_, _13323_, _02202_);
  or (_13325_, _13324_, _13321_);
  nor (_13326_, _11503_, _05439_);
  or (_13327_, _13234_, _04953_);
  or (_13328_, _13327_, _13326_);
  and (_13329_, _13328_, _04958_);
  and (_13330_, _13329_, _13325_);
  nor (_13331_, _11510_, _05439_);
  or (_13332_, _13331_, _13234_);
  and (_13333_, _13332_, _02334_);
  or (_13334_, _13333_, _02366_);
  or (_13335_, _13334_, _13330_);
  or (_13336_, _13245_, _02778_);
  and (_13337_, _13336_, _01698_);
  and (_13338_, _13337_, _13335_);
  and (_13339_, _13265_, _01697_);
  or (_13340_, _13339_, _02081_);
  or (_13341_, _13340_, _13338_);
  and (_13342_, _11567_, _03847_);
  or (_13343_, _13234_, _02082_);
  or (_13344_, _13343_, _13342_);
  and (_13345_, _13344_, _39632_);
  and (_13346_, _13345_, _13341_);
  or (_13347_, _13346_, _13233_);
  and (_41620_, _13347_, _39026_);
  nor (_13348_, _39632_, _06224_);
  nor (_13349_, _03847_, _06224_);
  nor (_13350_, _11704_, _05439_);
  or (_13351_, _13350_, _13349_);
  and (_13352_, _13351_, _01765_);
  nor (_13353_, _04478_, _06224_);
  and (_13354_, _11595_, _04478_);
  or (_13355_, _13354_, _13353_);
  and (_13356_, _13355_, _02053_);
  nor (_13357_, _04372_, _05439_);
  or (_13358_, _13357_, _13349_);
  or (_13359_, _13358_, _02519_);
  nor (_13360_, _11611_, _05439_);
  or (_13361_, _13360_, _13349_);
  or (_13362_, _13361_, _03006_);
  and (_13363_, _03847_, \oc8051_golden_model_1.ACC [4]);
  or (_13364_, _13363_, _13349_);
  and (_13365_, _13364_, _02062_);
  nor (_13366_, _02062_, _06224_);
  or (_13367_, _13366_, _02158_);
  or (_13368_, _13367_, _13365_);
  and (_13369_, _13368_, _02058_);
  and (_13370_, _13369_, _13362_);
  and (_13371_, _11597_, _04478_);
  or (_13372_, _13371_, _13353_);
  and (_13373_, _13372_, _02057_);
  or (_13374_, _13373_, _02155_);
  or (_13375_, _13374_, _13370_);
  and (_13376_, _13375_, _13359_);
  or (_13377_, _13376_, _02153_);
  or (_13378_, _13364_, _02549_);
  and (_13379_, _13378_, _02054_);
  and (_13380_, _13379_, _13377_);
  or (_13381_, _13380_, _13356_);
  and (_13382_, _13381_, _02047_);
  or (_13383_, _13353_, _11628_);
  and (_13384_, _13383_, _02046_);
  and (_13385_, _13384_, _13372_);
  or (_13386_, _13385_, _05474_);
  or (_13387_, _13386_, _13382_);
  nor (_13388_, _06162_, _06160_);
  nor (_13389_, _13388_, _06163_);
  or (_13390_, _13389_, _06181_);
  and (_13391_, _13390_, _02043_);
  and (_13392_, _13391_, _13387_);
  nor (_13393_, _11646_, _06189_);
  or (_13394_, _13393_, _13353_);
  and (_13395_, _13394_, _02042_);
  or (_13396_, _13395_, _06188_);
  or (_13397_, _13396_, _13392_);
  or (_13398_, _13358_, _05444_);
  and (_13399_, _13398_, _13397_);
  or (_13400_, _13399_, _02031_);
  and (_13401_, _05303_, _03847_);
  or (_13402_, _13349_, _02032_);
  or (_13403_, _13402_, _13401_);
  and (_13404_, _13403_, _02037_);
  and (_13405_, _13404_, _13400_);
  or (_13406_, _13405_, _13352_);
  and (_13407_, _13406_, _06560_);
  or (_13408_, _13176_, _06498_);
  nor (_13409_, _13293_, _06508_);
  or (_13410_, _13409_, _06507_);
  nand (_13411_, _13410_, _06547_);
  or (_13412_, _13410_, _06547_);
  and (_13413_, _13412_, _13411_);
  or (_13414_, _13413_, _06558_);
  and (_13415_, _13414_, _06202_);
  and (_13416_, _13415_, _13408_);
  or (_13417_, _13416_, _07629_);
  or (_13418_, _13417_, _13407_);
  and (_13419_, _11592_, _03847_);
  or (_13420_, _13349_, _03059_);
  or (_13421_, _13420_, _13419_);
  and (_13422_, _04831_, _03847_);
  or (_13423_, _13422_, _13349_);
  or (_13424_, _13423_, _01995_);
  and (_13425_, _13424_, _03061_);
  and (_13426_, _13425_, _13421_);
  and (_13427_, _13426_, _13418_);
  and (_13428_, _11588_, _03847_);
  or (_13429_, _13428_, _13349_);
  and (_13430_, _13429_, _02331_);
  or (_13431_, _13430_, _13427_);
  and (_13432_, _13431_, _02208_);
  or (_13433_, _13349_, _04420_);
  and (_13434_, _13423_, _02206_);
  and (_13435_, _13434_, _13433_);
  or (_13436_, _13435_, _13432_);
  and (_13437_, _13436_, _03065_);
  and (_13438_, _13364_, _02342_);
  and (_13439_, _13438_, _13433_);
  or (_13440_, _13439_, _02202_);
  or (_13441_, _13440_, _13437_);
  nor (_13442_, _11590_, _05439_);
  or (_13443_, _13349_, _04953_);
  or (_13444_, _13443_, _13442_);
  and (_13445_, _13444_, _04958_);
  and (_13446_, _13445_, _13441_);
  nor (_13447_, _11587_, _05439_);
  or (_13448_, _13447_, _13349_);
  and (_13449_, _13448_, _02334_);
  or (_13450_, _13449_, _02366_);
  or (_13451_, _13450_, _13446_);
  or (_13452_, _13361_, _02778_);
  and (_13453_, _13452_, _01698_);
  and (_13454_, _13453_, _13451_);
  and (_13455_, _13355_, _01697_);
  or (_13456_, _13455_, _02081_);
  or (_13457_, _13456_, _13454_);
  and (_13458_, _11771_, _03847_);
  or (_13459_, _13349_, _02082_);
  or (_13460_, _13459_, _13458_);
  and (_13461_, _13460_, _39632_);
  and (_13462_, _13461_, _13457_);
  or (_13463_, _13462_, _13348_);
  and (_41621_, _13463_, _39026_);
  nor (_13464_, _39632_, _06225_);
  nor (_13465_, _03847_, _06225_);
  nor (_13466_, _11900_, _05439_);
  or (_13467_, _13466_, _13465_);
  and (_13468_, _13467_, _01765_);
  nor (_13469_, _04057_, _05439_);
  or (_13470_, _13469_, _13465_);
  or (_13471_, _13470_, _05444_);
  or (_13472_, _13470_, _02519_);
  nor (_13473_, _11804_, _05439_);
  or (_13474_, _13473_, _13465_);
  or (_13475_, _13474_, _03006_);
  and (_13476_, _03847_, \oc8051_golden_model_1.ACC [5]);
  or (_13477_, _13476_, _13465_);
  and (_13478_, _13477_, _02062_);
  nor (_13479_, _02062_, _06225_);
  or (_13480_, _13479_, _02158_);
  or (_13481_, _13480_, _13478_);
  and (_13482_, _13481_, _02058_);
  and (_13483_, _13482_, _13475_);
  nor (_13484_, _04478_, _06225_);
  and (_13485_, _11789_, _04478_);
  or (_13486_, _13485_, _13484_);
  and (_13487_, _13486_, _02057_);
  or (_13488_, _13487_, _02155_);
  or (_13489_, _13488_, _13483_);
  and (_13490_, _13489_, _13472_);
  or (_13491_, _13490_, _02153_);
  or (_13492_, _13477_, _02549_);
  and (_13493_, _13492_, _02054_);
  and (_13494_, _13493_, _13491_);
  and (_13495_, _11816_, _04478_);
  or (_13496_, _13495_, _13484_);
  and (_13497_, _13496_, _02053_);
  or (_13498_, _13497_, _13494_);
  and (_13499_, _13498_, _02047_);
  or (_13500_, _13484_, _11823_);
  and (_13501_, _13500_, _02046_);
  and (_13502_, _13501_, _13486_);
  or (_13503_, _13502_, _05474_);
  or (_13504_, _13503_, _13499_);
  or (_13505_, _05744_, _05746_);
  and (_13506_, _13505_, _06164_);
  nor (_13507_, _13506_, _06165_);
  or (_13508_, _13507_, _06181_);
  and (_13509_, _13508_, _02043_);
  and (_13510_, _13509_, _13504_);
  nor (_13511_, _11841_, _06189_);
  or (_13512_, _13511_, _13484_);
  and (_13513_, _13512_, _02042_);
  or (_13514_, _13513_, _06188_);
  or (_13515_, _13514_, _13510_);
  and (_13516_, _13515_, _13471_);
  or (_13517_, _13516_, _02031_);
  and (_13518_, _05258_, _03847_);
  or (_13519_, _13465_, _02032_);
  or (_13520_, _13519_, _13518_);
  and (_13521_, _13520_, _02037_);
  and (_13522_, _13521_, _13517_);
  or (_13523_, _13522_, _13468_);
  and (_13524_, _13523_, _06560_);
  not (_13525_, _06536_);
  and (_13526_, _13411_, _13525_);
  nor (_13527_, _13526_, _06548_);
  and (_13528_, _13526_, _06548_);
  or (_13529_, _13528_, _13527_);
  nor (_13530_, _06558_, _06560_);
  and (_13531_, _13530_, _13529_);
  and (_13532_, _06490_, _06202_);
  and (_13533_, _13532_, _06558_);
  or (_13534_, _13533_, _07629_);
  or (_13535_, _13534_, _13531_);
  or (_13536_, _13535_, _13524_);
  and (_13537_, _11915_, _03847_);
  or (_13538_, _13465_, _03059_);
  or (_13539_, _13538_, _13537_);
  and (_13540_, _04827_, _03847_);
  or (_13541_, _13540_, _13465_);
  or (_13542_, _13541_, _01995_);
  and (_13543_, _13542_, _03061_);
  and (_13544_, _13543_, _13539_);
  and (_13545_, _13544_, _13536_);
  and (_13546_, _11786_, _03847_);
  or (_13547_, _13546_, _13465_);
  and (_13548_, _13547_, _02331_);
  or (_13549_, _13548_, _13545_);
  and (_13550_, _13549_, _02208_);
  or (_13551_, _13465_, _04104_);
  and (_13552_, _13541_, _02206_);
  and (_13553_, _13552_, _13551_);
  or (_13554_, _13553_, _13550_);
  and (_13555_, _13554_, _03065_);
  and (_13556_, _13477_, _02342_);
  and (_13557_, _13556_, _13551_);
  or (_13558_, _13557_, _02202_);
  or (_13559_, _13558_, _13555_);
  nor (_13560_, _11913_, _05439_);
  or (_13561_, _13465_, _04953_);
  or (_13562_, _13561_, _13560_);
  and (_13563_, _13562_, _04958_);
  and (_13564_, _13563_, _13559_);
  nor (_13565_, _11785_, _05439_);
  or (_13566_, _13565_, _13465_);
  and (_13567_, _13566_, _02334_);
  or (_13568_, _13567_, _02366_);
  or (_13569_, _13568_, _13564_);
  or (_13570_, _13474_, _02778_);
  and (_13571_, _13570_, _01698_);
  and (_13572_, _13571_, _13569_);
  and (_13573_, _13496_, _01697_);
  or (_13574_, _13573_, _02081_);
  or (_13575_, _13574_, _13572_);
  and (_13576_, _11974_, _03847_);
  or (_13577_, _13465_, _02082_);
  or (_13578_, _13577_, _13576_);
  and (_13579_, _13578_, _39632_);
  and (_13580_, _13579_, _13575_);
  or (_13581_, _13580_, _13464_);
  and (_41622_, _13581_, _39026_);
  nor (_13582_, _39632_, _06475_);
  nor (_13583_, _03847_, _06475_);
  nor (_13584_, _12096_, _05439_);
  or (_13585_, _13584_, _13583_);
  and (_13586_, _13585_, _01765_);
  nor (_13587_, _03964_, _05439_);
  or (_13588_, _13587_, _13583_);
  or (_13589_, _13588_, _05444_);
  or (_13590_, _13588_, _02519_);
  nor (_13591_, _11993_, _05439_);
  or (_13592_, _13591_, _13583_);
  or (_13593_, _13592_, _03006_);
  and (_13594_, _03847_, \oc8051_golden_model_1.ACC [6]);
  or (_13595_, _13594_, _13583_);
  and (_13596_, _13595_, _02062_);
  nor (_13597_, _02062_, _06475_);
  or (_13598_, _13597_, _02158_);
  or (_13599_, _13598_, _13596_);
  and (_13600_, _13599_, _02058_);
  and (_13601_, _13600_, _13593_);
  nor (_13602_, _04478_, _06475_);
  and (_13603_, _11990_, _04478_);
  or (_13604_, _13603_, _13602_);
  and (_13605_, _13604_, _02057_);
  or (_13606_, _13605_, _02155_);
  or (_13607_, _13606_, _13601_);
  and (_13608_, _13607_, _13590_);
  or (_13609_, _13608_, _02153_);
  or (_13610_, _13595_, _02549_);
  and (_13611_, _13610_, _02054_);
  and (_13612_, _13611_, _13609_);
  and (_13613_, _12017_, _04478_);
  or (_13614_, _13613_, _13602_);
  and (_13615_, _13614_, _02053_);
  or (_13616_, _13615_, _13612_);
  and (_13617_, _13616_, _02047_);
  or (_13618_, _13602_, _12024_);
  and (_13619_, _13618_, _02046_);
  and (_13620_, _13619_, _13604_);
  or (_13621_, _13620_, _05474_);
  or (_13622_, _13621_, _13617_);
  not (_13623_, _06180_);
  or (_13624_, _06179_, _06166_);
  and (_13625_, _13624_, _13623_);
  or (_13626_, _13625_, _06181_);
  and (_13627_, _13626_, _02043_);
  and (_13628_, _13627_, _13622_);
  nor (_13629_, _12042_, _06189_);
  or (_13630_, _13629_, _13602_);
  and (_13631_, _13630_, _02042_);
  or (_13632_, _13631_, _06188_);
  or (_13633_, _13632_, _13628_);
  and (_13634_, _13633_, _13589_);
  or (_13635_, _13634_, _02031_);
  and (_13636_, _05029_, _03847_);
  or (_13637_, _13583_, _02032_);
  or (_13638_, _13637_, _13636_);
  and (_13639_, _13638_, _02037_);
  and (_13640_, _13639_, _13635_);
  or (_13641_, _13640_, _13586_);
  and (_13642_, _13641_, _06560_);
  nor (_13643_, _13526_, _06491_);
  or (_13644_, _13643_, _06492_);
  or (_13645_, _13644_, _06545_);
  nand (_13646_, _13644_, _06545_);
  and (_13647_, _13646_, _13645_);
  or (_13648_, _13647_, _06558_);
  or (_13649_, _13176_, _06481_);
  and (_13650_, _13649_, _06202_);
  and (_13651_, _13650_, _13648_);
  or (_13652_, _13651_, _07629_);
  or (_13653_, _13652_, _13642_);
  and (_13654_, _12112_, _03847_);
  or (_13655_, _13583_, _03059_);
  or (_13656_, _13655_, _13654_);
  and (_13657_, _12103_, _03847_);
  or (_13658_, _13657_, _13583_);
  or (_13659_, _13658_, _01995_);
  and (_13660_, _13659_, _03061_);
  and (_13661_, _13660_, _13656_);
  and (_13662_, _13661_, _13653_);
  and (_13663_, _12118_, _03847_);
  or (_13664_, _13663_, _13583_);
  and (_13665_, _13664_, _02331_);
  or (_13666_, _13665_, _13662_);
  and (_13667_, _13666_, _02208_);
  or (_13668_, _13583_, _04011_);
  and (_13669_, _13658_, _02206_);
  and (_13670_, _13669_, _13668_);
  or (_13671_, _13670_, _13667_);
  and (_13672_, _13671_, _03065_);
  and (_13673_, _13595_, _02342_);
  and (_13674_, _13673_, _13668_);
  or (_13675_, _13674_, _02202_);
  or (_13676_, _13675_, _13672_);
  nor (_13677_, _12110_, _05439_);
  or (_13678_, _13583_, _04953_);
  or (_13679_, _13678_, _13677_);
  and (_13680_, _13679_, _04958_);
  and (_13681_, _13680_, _13676_);
  nor (_13682_, _12117_, _05439_);
  or (_13683_, _13682_, _13583_);
  and (_13684_, _13683_, _02334_);
  or (_13685_, _13684_, _02366_);
  or (_13686_, _13685_, _13681_);
  or (_13687_, _13592_, _02778_);
  and (_13688_, _13687_, _01698_);
  and (_13689_, _13688_, _13686_);
  and (_13690_, _13614_, _01697_);
  or (_13691_, _13690_, _02081_);
  or (_13692_, _13691_, _13689_);
  and (_13693_, _12178_, _03847_);
  or (_13694_, _13583_, _02082_);
  or (_13695_, _13694_, _13693_);
  and (_13696_, _13695_, _39632_);
  and (_13697_, _13696_, _13692_);
  or (_13698_, _13697_, _13582_);
  and (_41623_, _13698_, _39026_);
  nor (_13699_, _39632_, _01887_);
  nand (_13700_, _07533_, _04939_);
  nand (_13701_, _08874_, _02085_);
  and (_13702_, _13701_, _08458_);
  and (_13703_, _02236_, _01737_);
  nor (_13704_, _06611_, _02745_);
  nand (_13705_, _07338_, _08918_);
  nor (_13706_, _09037_, _02138_);
  nor (_13707_, _13706_, _10130_);
  and (_13708_, _02497_, _01727_);
  nor (_13709_, _13708_, _02895_);
  nand (_13710_, _02129_, _01727_);
  and (_13711_, _13710_, _13709_);
  not (_13712_, _13711_);
  and (_13713_, _13712_, _06637_);
  nor (_13714_, _03841_, _01887_);
  and (_13715_, _10914_, _03841_);
  nor (_13716_, _13715_, _13714_);
  nand (_13717_, _13716_, _02210_);
  nand (_13718_, _02027_, _01775_);
  nor (_13719_, _10898_, _06736_);
  nor (_13720_, _13719_, _13714_);
  nor (_13721_, _13720_, _02037_);
  and (_13722_, _03841_, _03002_);
  nor (_13723_, _13722_, _13714_);
  nand (_13724_, _13723_, _06188_);
  nand (_13725_, _07002_, _06815_);
  or (_13726_, _06820_, _03002_);
  nor (_13727_, _02552_, _02079_);
  or (_13728_, _13727_, _05120_);
  or (_13729_, _06852_, _03002_);
  nor (_13730_, _06855_, _01887_);
  and (_13731_, _06855_, _01887_);
  nor (_13732_, _13731_, _13730_);
  nand (_13733_, _13732_, _06859_);
  and (_13734_, _13733_, _13729_);
  or (_13735_, _13734_, _02160_);
  nand (_13736_, _07094_, _02160_);
  and (_13737_, _13736_, _10299_);
  and (_13738_, _13737_, _13735_);
  or (_13739_, _13738_, _02079_);
  and (_13740_, _13739_, _03006_);
  and (_13741_, _13740_, _13728_);
  nor (_13742_, _04257_, _06736_);
  nor (_13743_, _13742_, _13714_);
  nor (_13744_, _13743_, _03006_);
  or (_13745_, _13744_, _02057_);
  or (_13746_, _13745_, _13741_);
  nor (_13747_, _04483_, _01887_);
  and (_13748_, _10814_, _04483_);
  nor (_13749_, _13748_, _13747_);
  nand (_13750_, _13749_, _02057_);
  and (_13751_, _13750_, _02519_);
  and (_13752_, _13751_, _13746_);
  nor (_13753_, _13723_, _02519_);
  or (_13754_, _13753_, _06821_);
  or (_13755_, _13754_, _13752_);
  and (_13756_, _13755_, _13726_);
  or (_13757_, _13756_, _02582_);
  or (_13758_, _05120_, _06884_);
  and (_13759_, _13758_, _02549_);
  and (_13760_, _13759_, _13757_);
  nor (_13761_, _07094_, _02549_);
  or (_13762_, _13761_, _06888_);
  or (_13763_, _13762_, _13760_);
  nand (_13764_, _06888_, _06283_);
  and (_13765_, _13764_, _13763_);
  or (_13766_, _13765_, _02053_);
  or (_13767_, _13714_, _02054_);
  and (_13768_, _13767_, _02047_);
  and (_13769_, _13768_, _13766_);
  nor (_13770_, _13743_, _02047_);
  or (_13771_, _13770_, _05474_);
  or (_13772_, _13771_, _13769_);
  not (_13773_, _06127_);
  nand (_13774_, _13773_, _05474_);
  and (_13775_, _13774_, _06816_);
  and (_13776_, _13775_, _13772_);
  nor (_13777_, _06924_, _06816_);
  or (_13778_, _13777_, _06815_);
  or (_13779_, _13778_, _13776_);
  and (_13780_, _13779_, _13725_);
  or (_13781_, _13780_, _02186_);
  nand (_13782_, _07186_, _02186_);
  and (_13783_, _13782_, _06741_);
  and (_13784_, _13783_, _13781_);
  nor (_13785_, _06792_, _06741_);
  or (_13786_, _13785_, _01876_);
  or (_13787_, _13786_, _13784_);
  nand (_13788_, _02027_, _01876_);
  and (_13789_, _13788_, _02043_);
  and (_13790_, _13789_, _13787_);
  nor (_13791_, _10798_, _07215_);
  nor (_13792_, _13791_, _13747_);
  nor (_13793_, _13792_, _02043_);
  or (_13794_, _13793_, _06188_);
  or (_13795_, _13794_, _13790_);
  and (_13796_, _13795_, _13724_);
  or (_13797_, _13796_, _02031_);
  and (_13798_, _05120_, _03841_);
  nor (_13799_, _13798_, _13714_);
  nand (_13800_, _13799_, _02031_);
  and (_13801_, _13800_, _02037_);
  and (_13802_, _13801_, _13797_);
  or (_13803_, _13802_, _13721_);
  and (_13804_, _13803_, _06560_);
  or (_13805_, _13530_, _01775_);
  or (_13806_, _13805_, _13804_);
  and (_13807_, _13806_, _13718_);
  or (_13808_, _13807_, _01994_);
  and (_13809_, _03841_, _04837_);
  nor (_13810_, _13809_, _13714_);
  nand (_13811_, _13810_, _01994_);
  and (_13812_, _13811_, _07240_);
  and (_13813_, _13812_, _13808_);
  nor (_13814_, _07240_, _02027_);
  or (_13815_, _13814_, _07248_);
  nor (_13816_, _13815_, _13813_);
  and (_13817_, _03020_, _01887_);
  nor (_13818_, _13817_, _06637_);
  nor (_13819_, _07251_, _13818_);
  or (_13820_, _07260_, _07256_);
  or (_13821_, _13820_, _13819_);
  or (_13822_, _13821_, _13816_);
  and (_13823_, _13820_, _13818_);
  nor (_13824_, _13823_, _07263_);
  nand (_13825_, _13824_, _13822_);
  nor (_13826_, _05120_, \oc8051_golden_model_1.ACC [0]);
  nor (_13827_, _07468_, _13826_);
  or (_13828_, _13827_, _07264_);
  and (_13829_, _13828_, _13825_);
  or (_13830_, _13829_, _02329_);
  or (_13831_, _10792_, _02330_);
  and (_13832_, _13831_, _07281_);
  and (_13833_, _13832_, _13830_);
  and (_13834_, _06734_, _08919_);
  or (_13835_, _13834_, _02210_);
  or (_13836_, _13835_, _13833_);
  and (_13837_, _13836_, _13717_);
  or (_13838_, _13837_, _02331_);
  or (_13839_, _13714_, _03061_);
  and (_13840_, _13839_, _13711_);
  and (_13841_, _13840_, _13838_);
  or (_13842_, _13841_, _13713_);
  and (_13843_, _13842_, _07305_);
  and (_13844_, _07468_, _07304_);
  or (_13845_, _13844_, _02340_);
  or (_13846_, _13845_, _13843_);
  or (_13847_, _10791_, _02341_);
  and (_13848_, _13847_, _07313_);
  and (_13849_, _13848_, _13846_);
  and (_13850_, _07312_, _07553_);
  or (_13851_, _13850_, _13849_);
  and (_13852_, _13851_, _02208_);
  and (_13853_, _06732_, _05332_);
  nor (_13854_, _13810_, _13742_);
  and (_13855_, _13854_, _02206_);
  or (_13856_, _13855_, _13853_);
  or (_13857_, _13856_, _13852_);
  nand (_13858_, _13853_, _13817_);
  nand (_13859_, _13858_, _13857_);
  nor (_13860_, _13859_, _13707_);
  not (_13861_, _13707_);
  nor (_13862_, _13861_, _13817_);
  or (_13863_, _13862_, _10128_);
  or (_13864_, _13863_, _13860_);
  nor (_13865_, _13817_, _02719_);
  or (_13866_, _13865_, _10129_);
  and (_13867_, _13866_, _13864_);
  nor (_13868_, _13817_, _07327_);
  or (_13869_, _13868_, _07331_);
  or (_13870_, _13869_, _13867_);
  nand (_13871_, _13826_, _07331_);
  and (_13872_, _13871_, _02337_);
  and (_13873_, _13872_, _13870_);
  nand (_13874_, _10789_, _07341_);
  and (_13875_, _13874_, _07340_);
  or (_13876_, _13875_, _13873_);
  and (_13877_, _13876_, _13705_);
  or (_13878_, _13877_, _02202_);
  nor (_13879_, _10913_, _06736_);
  nor (_13880_, _13879_, _13714_);
  nand (_13881_, _13880_, _02202_);
  and (_13882_, _13881_, _06729_);
  and (_13883_, _13882_, _13878_);
  nor (_13884_, _06924_, _06729_);
  or (_13885_, _13884_, _06727_);
  or (_13886_, _13885_, _13883_);
  nor (_13887_, _06924_, _06654_);
  or (_13888_, _13887_, _02731_);
  and (_13889_, _13888_, _13886_);
  nor (_13890_, _07002_, _07356_);
  or (_13891_, _13890_, _02345_);
  or (_13892_, _13891_, _13889_);
  nand (_13893_, _07186_, _02345_);
  and (_13894_, _13893_, _07417_);
  and (_13895_, _13894_, _13892_);
  nor (_13896_, _07417_, _06792_);
  or (_13897_, _13896_, _07415_);
  or (_13898_, _13897_, _13895_);
  nor (_13899_, _09038_, _02499_);
  and (_13900_, _07415_, _06707_);
  nor (_13901_, _13900_, _13899_);
  and (_13902_, _13901_, _13898_);
  and (_13903_, _13899_, _13818_);
  nor (_13904_, _13903_, _13902_);
  nand (_13905_, _13904_, _13704_);
  or (_13906_, _13704_, _13818_);
  nand (_13907_, _13906_, _13905_);
  nor (_13908_, _13907_, _13703_);
  and (_13909_, _13703_, _13827_);
  nor (_13910_, _13909_, _13908_);
  nor (_13911_, _13910_, _02748_);
  and (_13912_, _13827_, _02748_);
  or (_13913_, _13912_, _13911_);
  or (_13914_, _13913_, _02085_);
  and (_13915_, _13914_, _13702_);
  and (_13916_, _07487_, _08919_);
  or (_13917_, _13916_, _07533_);
  or (_13918_, _13917_, _13915_);
  and (_13919_, _13918_, _13700_);
  or (_13920_, _13919_, _02366_);
  nand (_13921_, _13743_, _02366_);
  and (_13922_, _13921_, _07576_);
  and (_13923_, _13922_, _13920_);
  nor (_13924_, _07580_, _01887_);
  nor (_13925_, _13924_, _07581_);
  or (_13926_, _13925_, _13923_);
  nand (_13927_, _07580_, _01804_);
  and (_13928_, _13927_, _01698_);
  and (_13929_, _13928_, _13926_);
  and (_13930_, _13714_, _01697_);
  or (_13931_, _13930_, _02081_);
  or (_13932_, _13931_, _13929_);
  nand (_13933_, _13743_, _02081_);
  and (_13934_, _13933_, _07600_);
  and (_13935_, _13934_, _13932_);
  nor (_13936_, _07606_, _01887_);
  nor (_13937_, _13936_, _10751_);
  or (_13938_, _13937_, _13935_);
  nand (_13939_, _07606_, _01804_);
  and (_13940_, _13939_, _39632_);
  and (_13941_, _13940_, _13938_);
  or (_13942_, _13941_, _13699_);
  and (_41625_, _13942_, _39026_);
  nor (_13943_, _39632_, _01804_);
  and (_13944_, _07424_, _06786_);
  nor (_13945_, _13944_, _07425_);
  or (_13946_, _13945_, _07417_);
  nand (_13947_, _07466_, _07331_);
  not (_13948_, _10131_);
  nand (_13949_, _13948_, _06635_);
  or (_13950_, _07465_, _07305_);
  nor (_13951_, _03841_, _01804_);
  and (_13952_, _10989_, _03841_);
  nor (_13953_, _13952_, _13951_);
  nand (_13954_, _13953_, _02210_);
  or (_13955_, _11113_, _02330_);
  and (_13956_, _13955_, _07281_);
  nand (_13957_, _02859_, _01775_);
  nor (_13958_, _06736_, _03161_);
  nor (_13959_, _13958_, _13951_);
  nand (_13960_, _13959_, _06188_);
  nand (_13961_, _06821_, _03161_);
  nor (_13962_, _06825_, \oc8051_golden_model_1.PSW [6]);
  nor (_13963_, _13962_, \oc8051_golden_model_1.ACC [1]);
  and (_13964_, _13962_, \oc8051_golden_model_1.ACC [1]);
  nor (_13965_, _13964_, _13963_);
  nand (_13966_, _13965_, _06823_);
  or (_13967_, _13727_, _05075_);
  nand (_13968_, _06853_, _03161_);
  or (_13969_, _06855_, \oc8051_golden_model_1.ACC [1]);
  nand (_13970_, _06855_, \oc8051_golden_model_1.ACC [1]);
  nand (_13971_, _13970_, _13969_);
  nand (_13972_, _13971_, _06859_);
  and (_13973_, _13972_, _13968_);
  or (_13974_, _13973_, _02160_);
  nand (_13975_, _07082_, _02160_);
  and (_13976_, _13975_, _10299_);
  and (_13977_, _13976_, _13974_);
  or (_13978_, _13977_, _02079_);
  and (_13979_, _13978_, _03006_);
  and (_13980_, _13979_, _13967_);
  nor (_13981_, _03841_, \oc8051_golden_model_1.ACC [1]);
  and (_13982_, _11001_, _03841_);
  nor (_13983_, _13982_, _13981_);
  and (_13984_, _13983_, _02158_);
  or (_13985_, _13984_, _06823_);
  or (_13986_, _13985_, _13980_);
  and (_13987_, _13986_, _13966_);
  or (_13988_, _13987_, _02057_);
  nor (_13989_, _04483_, _01804_);
  and (_13990_, _11005_, _04483_);
  nor (_13991_, _13990_, _13989_);
  nand (_13992_, _13991_, _02057_);
  and (_13993_, _13992_, _02519_);
  and (_13994_, _13993_, _13988_);
  nor (_13995_, _13959_, _02519_);
  or (_13996_, _13995_, _06821_);
  or (_13997_, _13996_, _13994_);
  and (_13998_, _13997_, _13961_);
  or (_13999_, _13998_, _02582_);
  or (_14000_, _05075_, _06884_);
  and (_14001_, _14000_, _02549_);
  and (_14002_, _14001_, _13999_);
  nor (_14003_, _07082_, _02549_);
  or (_14004_, _14003_, _06888_);
  or (_14005_, _14004_, _14002_);
  nand (_14006_, _06888_, _06277_);
  and (_14007_, _14006_, _14005_);
  or (_14008_, _14007_, _02053_);
  and (_14009_, _10992_, _04483_);
  nor (_14010_, _14009_, _13989_);
  nand (_14011_, _14010_, _02053_);
  and (_14012_, _14011_, _02047_);
  and (_14013_, _14012_, _14008_);
  and (_14014_, _13990_, _11020_);
  nor (_14015_, _14014_, _13989_);
  nor (_14016_, _14015_, _02047_);
  or (_14017_, _14016_, _05474_);
  or (_14018_, _14017_, _14013_);
  and (_14019_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_14020_, _14019_, _06520_);
  nor (_14021_, _14020_, _06128_);
  or (_14022_, _14021_, _06181_);
  and (_14023_, _14022_, _06816_);
  and (_14024_, _14023_, _14018_);
  not (_14025_, _07191_);
  and (_14026_, _14025_, _03002_);
  nor (_14027_, _14026_, _07190_);
  and (_14028_, _14027_, _06636_);
  nor (_14029_, _14027_, _06636_);
  or (_14030_, _14029_, _14028_);
  and (_14031_, _14030_, _06817_);
  or (_14032_, _14031_, _06815_);
  or (_14033_, _14032_, _14024_);
  and (_14034_, _14025_, _05120_);
  nor (_14035_, _14034_, _07190_);
  and (_14036_, _14035_, _07467_);
  nor (_14037_, _14035_, _07467_);
  or (_14038_, _14037_, _14036_);
  or (_14039_, _14038_, _06941_);
  and (_14040_, _14039_, _02191_);
  and (_14041_, _14040_, _14033_);
  nor (_14042_, _07196_, _02191_);
  or (_14043_, _14042_, _14041_);
  and (_14044_, _14043_, _06741_);
  nor (_14045_, _07191_, _02027_);
  nor (_14046_, _14045_, _07190_);
  and (_14047_, _14046_, _07552_);
  nor (_14048_, _14046_, _07552_);
  nor (_14049_, _14048_, _14047_);
  nor (_14050_, _14049_, _06741_);
  or (_14051_, _14050_, _01876_);
  or (_14052_, _14051_, _14044_);
  nand (_14053_, _02859_, _01876_);
  and (_14054_, _14053_, _02043_);
  and (_14055_, _14054_, _14052_);
  nor (_14056_, _11038_, _07215_);
  nor (_14057_, _14056_, _13989_);
  nor (_14058_, _14057_, _02043_);
  or (_14059_, _14058_, _06188_);
  or (_14060_, _14059_, _14055_);
  and (_14061_, _14060_, _13960_);
  or (_14062_, _14061_, _02031_);
  and (_14063_, _05075_, _03841_);
  nor (_14064_, _14063_, _13951_);
  nand (_14065_, _14064_, _02031_);
  and (_14066_, _14065_, _02037_);
  and (_14067_, _14066_, _14062_);
  nor (_14068_, _11096_, _06736_);
  nor (_14069_, _14068_, _13951_);
  nor (_14070_, _14069_, _02037_);
  or (_14071_, _14070_, _06202_);
  or (_14072_, _14071_, _14067_);
  nand (_14073_, _06468_, _06202_);
  and (_14074_, _14073_, _14072_);
  or (_14075_, _14074_, _01775_);
  and (_14076_, _14075_, _13957_);
  or (_14077_, _14076_, _01994_);
  and (_14078_, _03841_, _02893_);
  nor (_14079_, _14078_, _13981_);
  or (_14080_, _14079_, _01995_);
  and (_14081_, _14080_, _07240_);
  nand (_14082_, _14081_, _14077_);
  or (_14083_, _07240_, _02859_);
  and (_14084_, _14083_, _07251_);
  and (_14085_, _14084_, _14082_);
  nor (_14086_, _07251_, _06636_);
  not (_14087_, _07258_);
  nand (_14088_, _14087_, _07253_);
  or (_14089_, _14088_, _14086_);
  nor (_14090_, _14089_, _14085_);
  and (_14091_, _14088_, _06636_);
  or (_14092_, _14091_, _07259_);
  or (_14093_, _14092_, _14090_);
  and (_14094_, _02132_, _01721_);
  not (_14095_, _14094_);
  or (_14096_, _06636_, _14095_);
  and (_14097_, _14096_, _14093_);
  or (_14098_, _14097_, _07263_);
  or (_14099_, _07467_, _07264_);
  and (_14100_, _14099_, _14098_);
  or (_14101_, _14100_, _02329_);
  and (_14102_, _14101_, _13956_);
  and (_14103_, _06734_, _07552_);
  or (_14104_, _14103_, _02210_);
  or (_14105_, _14104_, _14102_);
  and (_14106_, _14105_, _13954_);
  or (_14107_, _14106_, _02331_);
  or (_14108_, _13951_, _03061_);
  and (_14109_, _14108_, _13711_);
  and (_14110_, _14109_, _14107_);
  and (_14111_, _13712_, _06634_);
  or (_14112_, _14111_, _07304_);
  or (_14113_, _14112_, _14110_);
  and (_14114_, _14113_, _13950_);
  or (_14115_, _14114_, _02340_);
  or (_14116_, _11111_, _02341_);
  and (_14117_, _14116_, _07313_);
  and (_14118_, _14117_, _14115_);
  and (_14119_, _07312_, _07550_);
  or (_14120_, _14119_, _14118_);
  and (_14121_, _14120_, _02208_);
  and (_14122_, _10988_, _03841_);
  nor (_14123_, _14122_, _13951_);
  nor (_14124_, _14123_, _02208_);
  or (_14125_, _14124_, _13948_);
  or (_14126_, _14125_, _14121_);
  and (_14127_, _14126_, _13949_);
  or (_14128_, _14127_, _10128_);
  nor (_14129_, _06635_, _02719_);
  or (_14130_, _14129_, _10129_);
  and (_14131_, _14130_, _14128_);
  nor (_14132_, _06635_, _07327_);
  or (_14133_, _14132_, _07331_);
  or (_14134_, _14133_, _14131_);
  and (_14135_, _14134_, _13947_);
  or (_14136_, _14135_, _02336_);
  nand (_14137_, _11112_, _02336_);
  and (_14138_, _14137_, _07341_);
  and (_14139_, _14138_, _14136_);
  nor (_14140_, _07341_, _07551_);
  or (_14141_, _14140_, _02202_);
  or (_14142_, _14141_, _14139_);
  nor (_14143_, _10987_, _06736_);
  or (_14144_, _14143_, _13951_);
  or (_14145_, _14144_, _04953_);
  and (_14146_, _14145_, _06730_);
  and (_14147_, _14146_, _14142_);
  and (_14148_, _06711_, _06706_);
  nor (_14149_, _14148_, _06712_);
  and (_14150_, _14149_, _07348_);
  or (_14151_, _14150_, _06654_);
  or (_14152_, _14151_, _14147_);
  and (_14153_, _07365_, _07000_);
  nor (_14154_, _14153_, _07366_);
  or (_14155_, _14154_, _07356_);
  and (_14156_, _14155_, _02346_);
  and (_14157_, _14156_, _14152_);
  and (_14158_, _07396_, _07394_);
  nor (_14159_, _14158_, _07397_);
  or (_14160_, _14159_, _07384_);
  and (_14161_, _14160_, _07386_);
  or (_14162_, _14161_, _14157_);
  and (_14163_, _14162_, _13946_);
  or (_14164_, _14163_, _07415_);
  nand (_14165_, _07415_, _01887_);
  and (_14166_, _14165_, _06614_);
  and (_14167_, _14166_, _14164_);
  nor (_14168_, _06637_, _06636_);
  nor (_14169_, _14168_, _06638_);
  and (_14170_, _14169_, _09155_);
  or (_14171_, _14170_, _06609_);
  or (_14172_, _14171_, _14167_);
  nor (_14173_, _07468_, _07467_);
  nor (_14174_, _14173_, _07469_);
  or (_14175_, _14174_, _07448_);
  and (_14176_, _14175_, _02087_);
  and (_14177_, _14176_, _14172_);
  and (_14178_, _07512_, _07189_);
  nor (_14179_, _14178_, _07513_);
  or (_14180_, _14179_, _07487_);
  and (_14181_, _14180_, _07489_);
  or (_14182_, _14181_, _14177_);
  nor (_14183_, _07553_, _07552_);
  nor (_14184_, _14183_, _07554_);
  or (_14185_, _14184_, _08458_);
  and (_14186_, _14185_, _07534_);
  and (_14187_, _14186_, _14182_);
  and (_14188_, _07533_, \oc8051_golden_model_1.ACC [0]);
  or (_14189_, _14188_, _02366_);
  or (_14190_, _14189_, _14187_);
  or (_14191_, _13983_, _02778_);
  and (_14192_, _14191_, _07576_);
  and (_14193_, _14192_, _14190_);
  nor (_14194_, _07607_, _07582_);
  nor (_14195_, _14194_, _07576_);
  or (_14196_, _14195_, _07580_);
  or (_14197_, _14196_, _14193_);
  nand (_14198_, _07580_, _06383_);
  and (_14199_, _14198_, _01698_);
  and (_14200_, _14199_, _14197_);
  nor (_14201_, _14010_, _01698_);
  or (_14202_, _14201_, _02081_);
  or (_14203_, _14202_, _14200_);
  nor (_14204_, _13982_, _13951_);
  nand (_14205_, _14204_, _02081_);
  and (_14206_, _14205_, _07600_);
  and (_14207_, _14206_, _14203_);
  and (_14208_, _14194_, _07599_);
  or (_14209_, _14208_, _07606_);
  or (_14210_, _14209_, _14207_);
  nand (_14211_, _07606_, _06383_);
  and (_14212_, _14211_, _39632_);
  and (_14213_, _14212_, _14210_);
  or (_14214_, _14213_, _13943_);
  and (_41626_, _14214_, _39026_);
  nor (_14215_, _39632_, _06383_);
  and (_14216_, _06639_, _06633_);
  nor (_14217_, _14216_, _06640_);
  nor (_14218_, _05442_, _02499_);
  nand (_14219_, _14218_, _14217_);
  nand (_14220_, _07338_, _07547_);
  nor (_14221_, _02134_, _10130_);
  and (_14222_, _13712_, _06630_);
  nor (_14223_, _03841_, _06383_);
  and (_14224_, _11189_, _03841_);
  nor (_14225_, _14224_, _14223_);
  nand (_14226_, _14225_, _02210_);
  or (_14227_, _14087_, _06632_);
  nand (_14228_, _02452_, _01775_);
  nor (_14229_, _06736_, _03624_);
  nor (_14230_, _14229_, _14223_);
  nand (_14231_, _14230_, _06188_);
  nand (_14232_, _06821_, _03624_);
  nand (_14233_, _13962_, \oc8051_golden_model_1.ACC [2]);
  and (_14234_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_14235_, _14234_, _06824_);
  or (_14236_, _14235_, _13962_);
  and (_14237_, _14236_, _14233_);
  nand (_14238_, _14237_, _06823_);
  nand (_14239_, _06853_, _03624_);
  or (_14240_, _06855_, \oc8051_golden_model_1.ACC [2]);
  nand (_14241_, _06855_, \oc8051_golden_model_1.ACC [2]);
  nand (_14242_, _14241_, _14240_);
  nand (_14243_, _14242_, _06859_);
  and (_14244_, _14243_, _14239_);
  or (_14245_, _14244_, _02160_);
  nand (_14246_, _07068_, _02160_);
  and (_14247_, _14246_, _10299_);
  and (_14248_, _14247_, _14245_);
  or (_14249_, _14248_, _02079_);
  or (_14250_, _13727_, _05211_);
  and (_14251_, _14250_, _14249_);
  and (_14252_, _14251_, _03006_);
  nor (_14253_, _11199_, _06736_);
  nor (_14254_, _14253_, _14223_);
  nor (_14255_, _14254_, _03006_);
  or (_14256_, _14255_, _06823_);
  or (_14257_, _14256_, _14252_);
  and (_14258_, _14257_, _14238_);
  or (_14259_, _14258_, _02057_);
  nor (_14260_, _04483_, _06383_);
  and (_14261_, _11194_, _04483_);
  nor (_14262_, _14261_, _14260_);
  nand (_14263_, _14262_, _02057_);
  and (_14264_, _14263_, _02519_);
  and (_14265_, _14264_, _14259_);
  nor (_14266_, _14230_, _02519_);
  or (_14267_, _14266_, _06821_);
  or (_14268_, _14267_, _14265_);
  and (_14269_, _14268_, _14232_);
  or (_14270_, _14269_, _02582_);
  or (_14271_, _05211_, _06884_);
  and (_14272_, _14271_, _02549_);
  and (_14273_, _14272_, _14270_);
  nor (_14274_, _07068_, _02549_);
  or (_14275_, _14274_, _06888_);
  or (_14276_, _14275_, _14273_);
  nand (_14277_, _06888_, _06231_);
  and (_14278_, _14277_, _14276_);
  or (_14279_, _14278_, _02053_);
  and (_14280_, _11192_, _04483_);
  nor (_14281_, _14280_, _14260_);
  nand (_14282_, _14281_, _02053_);
  and (_14283_, _14282_, _02047_);
  and (_14284_, _14283_, _14279_);
  and (_14285_, _14261_, _11223_);
  nor (_14286_, _14285_, _14260_);
  nor (_14287_, _14286_, _02047_);
  or (_14288_, _14287_, _05474_);
  or (_14289_, _14288_, _14284_);
  nor (_14290_, _06130_, _06128_);
  nor (_14291_, _14290_, _06131_);
  or (_14292_, _14291_, _06181_);
  and (_14293_, _14292_, _14289_);
  or (_14294_, _14293_, _06817_);
  and (_14295_, _03161_, \oc8051_golden_model_1.ACC [1]);
  and (_14296_, _03002_, _01887_);
  nor (_14297_, _14296_, _06636_);
  nor (_14298_, _14297_, _14295_);
  nor (_14299_, _06632_, _14298_);
  and (_14300_, _06632_, _14298_);
  nor (_14301_, _14300_, _14299_);
  nor (_14302_, _13818_, _06636_);
  not (_14303_, _14302_);
  or (_14304_, _14303_, _14301_);
  and (_14305_, _14304_, \oc8051_golden_model_1.PSW [7]);
  nor (_14306_, _14301_, \oc8051_golden_model_1.PSW [7]);
  or (_14307_, _14306_, _14305_);
  nand (_14308_, _14303_, _14301_);
  and (_14309_, _14308_, _14307_);
  nand (_14310_, _14309_, _06817_);
  and (_14311_, _14310_, _06941_);
  and (_14312_, _14311_, _14294_);
  nor (_14313_, _05075_, _01804_);
  not (_14314_, _14313_);
  and (_14315_, _05120_, _01887_);
  or (_14316_, _14315_, _07467_);
  and (_14317_, _14316_, _14314_);
  nor (_14318_, _07463_, _14317_);
  and (_14319_, _07463_, _14317_);
  nor (_14320_, _14319_, _14318_);
  nor (_14321_, _13827_, _07467_);
  and (_14322_, _14321_, \oc8051_golden_model_1.PSW [7]);
  not (_14323_, _14322_);
  nor (_14324_, _14323_, _14320_);
  and (_14325_, _14323_, _14320_);
  nor (_14326_, _14325_, _14324_);
  nor (_14327_, _14326_, _06941_);
  or (_14328_, _14327_, _02186_);
  or (_14329_, _14328_, _14312_);
  nor (_14330_, _08873_, _07187_);
  or (_14331_, _14330_, _07188_);
  and (_14332_, _07509_, _14331_);
  nor (_14333_, _07509_, _14331_);
  nor (_14334_, _14333_, _14332_);
  and (_14335_, _08875_, \oc8051_golden_model_1.PSW [7]);
  not (_14336_, _14335_);
  nor (_14337_, _14336_, _14334_);
  and (_14338_, _14336_, _14334_);
  nor (_14339_, _14338_, _14337_);
  nand (_14340_, _14339_, _02186_);
  and (_14341_, _14340_, _06741_);
  and (_14342_, _14341_, _14329_);
  nor (_14343_, _02027_, \oc8051_golden_model_1.ACC [0]);
  nor (_14344_, _14343_, _07552_);
  nor (_14345_, _14344_, _08886_);
  nor (_14346_, _07548_, _14345_);
  and (_14347_, _07548_, _14345_);
  nor (_14348_, _14347_, _14346_);
  and (_14349_, _08920_, \oc8051_golden_model_1.PSW [7]);
  and (_14350_, _14349_, _14348_);
  nor (_14351_, _14349_, _14348_);
  or (_14352_, _14351_, _14350_);
  nor (_14353_, _14352_, _06741_);
  or (_14354_, _14353_, _01876_);
  or (_14355_, _14354_, _14342_);
  nand (_14356_, _02452_, _01876_);
  and (_14357_, _14356_, _02043_);
  and (_14358_, _14357_, _14355_);
  nor (_14359_, _11241_, _07215_);
  nor (_14360_, _14359_, _14260_);
  nor (_14361_, _14360_, _02043_);
  or (_14362_, _14361_, _06188_);
  or (_14363_, _14362_, _14358_);
  and (_14364_, _14363_, _14231_);
  or (_14365_, _14364_, _02031_);
  and (_14366_, _05211_, _03841_);
  nor (_14367_, _14366_, _14223_);
  nand (_14368_, _14367_, _02031_);
  and (_14369_, _14368_, _02037_);
  and (_14370_, _14369_, _14365_);
  nor (_14371_, _11298_, _06736_);
  nor (_14372_, _14371_, _14223_);
  nor (_14373_, _14372_, _02037_);
  or (_14374_, _14373_, _06202_);
  or (_14375_, _14374_, _14370_);
  or (_14376_, _06398_, _06560_);
  and (_14377_, _14376_, _14375_);
  or (_14378_, _14377_, _01775_);
  and (_14379_, _14378_, _14228_);
  or (_14380_, _14379_, _01994_);
  and (_14381_, _03841_, _04866_);
  nor (_14382_, _14381_, _14223_);
  nand (_14383_, _14382_, _01994_);
  and (_14384_, _14383_, _07240_);
  and (_14385_, _14384_, _14380_);
  nor (_14386_, _07240_, _02452_);
  or (_14387_, _14386_, _07248_);
  or (_14388_, _14387_, _14385_);
  or (_14389_, _07251_, _06632_);
  and (_14390_, _14389_, _07253_);
  and (_14391_, _14390_, _14388_);
  and (_14392_, _07256_, _06632_);
  or (_14393_, _14392_, _07258_);
  or (_14394_, _14393_, _14391_);
  and (_14395_, _14394_, _14227_);
  or (_14396_, _14395_, _14094_);
  and (_14397_, _02236_, _01721_);
  not (_14398_, _14397_);
  or (_14399_, _06632_, _14095_);
  and (_14400_, _14399_, _14398_);
  and (_14401_, _14400_, _14396_);
  or (_14402_, _07463_, _01598_);
  and (_14403_, _14402_, _07263_);
  or (_14404_, _14403_, _14401_);
  not (_14405_, _02696_);
  or (_14406_, _07463_, _14405_);
  and (_14407_, _14406_, _14404_);
  or (_14408_, _14407_, _02329_);
  or (_14409_, _11315_, _02330_);
  and (_14410_, _14409_, _07281_);
  and (_14411_, _14410_, _14408_);
  and (_14412_, _06734_, _07548_);
  or (_14413_, _14412_, _02210_);
  or (_14414_, _14413_, _14411_);
  and (_14415_, _14414_, _14226_);
  or (_14416_, _14415_, _02331_);
  or (_14417_, _14223_, _03061_);
  and (_14418_, _14417_, _13711_);
  and (_14419_, _14418_, _14416_);
  or (_14420_, _14419_, _14222_);
  and (_14421_, _14420_, _07305_);
  and (_14422_, _07461_, _07304_);
  or (_14423_, _14422_, _02340_);
  or (_14424_, _14423_, _14421_);
  or (_14425_, _11313_, _02341_);
  and (_14426_, _14425_, _07313_);
  and (_14427_, _14426_, _14424_);
  and (_14428_, _07312_, _07546_);
  or (_14429_, _14428_, _14427_);
  and (_14430_, _14429_, _02208_);
  or (_14431_, _14382_, _11314_);
  or (_14432_, _14431_, _02208_);
  nor (_14433_, _06732_, _02905_);
  nand (_14434_, _14433_, _14432_);
  or (_14435_, _14434_, _14430_);
  not (_14436_, _06631_);
  or (_14437_, _14433_, _14436_);
  nand (_14438_, _14437_, _14435_);
  nor (_14439_, _14438_, _14221_);
  and (_14440_, _14221_, _14436_);
  or (_14441_, _14440_, _07331_);
  or (_14442_, _14441_, _14439_);
  nand (_14443_, _07462_, _07331_);
  and (_14444_, _14443_, _02337_);
  and (_14445_, _14444_, _14442_);
  nand (_14446_, _11314_, _07341_);
  and (_14447_, _14446_, _07340_);
  or (_14448_, _14447_, _14445_);
  and (_14449_, _14448_, _14220_);
  or (_14450_, _14449_, _02202_);
  nor (_14451_, _11187_, _06736_);
  nor (_14452_, _14451_, _14223_);
  nand (_14453_, _14452_, _02202_);
  and (_14454_, _14453_, _06730_);
  and (_14455_, _14454_, _14450_);
  and (_14456_, _06713_, _06699_);
  nor (_14457_, _14456_, _06714_);
  and (_14458_, _14457_, _07348_);
  nor (_14459_, _14458_, _14455_);
  nor (_14460_, _14459_, _06654_);
  and (_14461_, _07367_, _06983_);
  nor (_14462_, _14461_, _07368_);
  and (_14463_, _14462_, _06654_);
  or (_14464_, _14463_, _02345_);
  or (_14465_, _14464_, _14460_);
  and (_14466_, _07398_, _07168_);
  nor (_14467_, _14466_, _07399_);
  or (_14468_, _14467_, _02346_);
  and (_14469_, _14468_, _07417_);
  and (_14470_, _14469_, _14465_);
  and (_14471_, _07426_, _06779_);
  nor (_14472_, _14471_, _07427_);
  and (_14473_, _14472_, _07384_);
  or (_14474_, _14473_, _07415_);
  or (_14475_, _14474_, _14470_);
  not (_14476_, _14218_);
  nand (_14477_, _07415_, _01804_);
  and (_14478_, _14477_, _14476_);
  nand (_14479_, _14478_, _14475_);
  and (_14480_, _14479_, _14219_);
  nor (_14481_, _14480_, _02747_);
  and (_14482_, _14217_, _02747_);
  or (_14483_, _14482_, _06609_);
  or (_14484_, _14483_, _14481_);
  and (_14485_, _07470_, _07464_);
  nor (_14486_, _14485_, _07471_);
  or (_14487_, _14486_, _07448_);
  and (_14488_, _14487_, _02087_);
  and (_14489_, _14488_, _14484_);
  and (_14490_, _07514_, _07509_);
  nor (_14491_, _14490_, _07515_);
  and (_14492_, _14491_, _02085_);
  or (_14493_, _14492_, _07487_);
  or (_14494_, _14493_, _14489_);
  and (_14495_, _07555_, _07549_);
  nor (_14496_, _14495_, _07556_);
  or (_14497_, _14496_, _08458_);
  and (_14498_, _14497_, _07534_);
  and (_14499_, _14498_, _14494_);
  and (_14500_, _07533_, \oc8051_golden_model_1.ACC [1]);
  or (_14501_, _14500_, _02366_);
  or (_14502_, _14501_, _14499_);
  nand (_14503_, _14254_, _02366_);
  and (_14504_, _14503_, _07576_);
  and (_14505_, _14504_, _14502_);
  and (_14506_, _06824_, _01887_);
  nor (_14507_, _07582_, _06383_);
  or (_14508_, _14507_, _14506_);
  and (_14509_, _14508_, _07575_);
  or (_14510_, _14509_, _07580_);
  or (_14511_, _14510_, _14505_);
  nand (_14512_, _07580_, _06377_);
  and (_14513_, _14512_, _01698_);
  and (_14514_, _14513_, _14511_);
  nor (_14515_, _14281_, _01698_);
  or (_14516_, _14515_, _02081_);
  or (_14517_, _14516_, _14514_);
  and (_14518_, _11367_, _03841_);
  nor (_14519_, _14518_, _14223_);
  nand (_14520_, _14519_, _02081_);
  and (_14521_, _14520_, _07600_);
  and (_14522_, _14521_, _14517_);
  and (_14523_, _07607_, \oc8051_golden_model_1.ACC [2]);
  nor (_14524_, _07607_, \oc8051_golden_model_1.ACC [2]);
  nor (_14525_, _14524_, _14523_);
  nor (_14526_, _14525_, _07606_);
  nor (_14527_, _14526_, _10751_);
  or (_14528_, _14527_, _14522_);
  nand (_14529_, _07606_, _06377_);
  and (_14530_, _14529_, _39632_);
  and (_14531_, _14530_, _14528_);
  or (_14532_, _14531_, _14215_);
  and (_41627_, _14532_, _39026_);
  nor (_14533_, _39632_, _06377_);
  nor (_14534_, _06627_, _06629_);
  nor (_14535_, _06641_, _14534_);
  and (_14536_, _06641_, _14534_);
  nor (_14537_, _14536_, _14535_);
  nand (_14538_, _14537_, _09155_);
  nor (_14539_, _03841_, _06377_);
  nor (_14540_, _11503_, _06736_);
  nor (_14541_, _14540_, _14539_);
  nor (_14542_, _14541_, _04953_);
  nand (_14543_, _13948_, _06629_);
  and (_14544_, _11505_, _03841_);
  nor (_14545_, _14544_, _14539_);
  nand (_14546_, _14545_, _02210_);
  and (_14547_, _02239_, _01721_);
  not (_14548_, _14547_);
  and (_14549_, _02137_, _01773_);
  and (_14550_, _14549_, _01721_);
  nor (_14551_, _14550_, _02902_);
  and (_14552_, _14551_, _14548_);
  or (_14553_, _14552_, _14534_);
  nand (_14554_, _01983_, _01775_);
  nor (_14555_, _06736_, _03434_);
  nor (_14556_, _14555_, _14539_);
  nand (_14557_, _14556_, _06188_);
  and (_14558_, _14320_, \oc8051_golden_model_1.PSW [7]);
  nor (_14559_, _14321_, _06707_);
  or (_14560_, _14559_, _14558_);
  nor (_14561_, _05211_, _06383_);
  nor (_14562_, _14318_, _14561_);
  nor (_14563_, _07459_, _07457_);
  not (_14564_, _14563_);
  nand (_14565_, _14564_, _14562_);
  or (_14566_, _14564_, _14562_);
  and (_14567_, _14566_, _14565_);
  or (_14568_, _14567_, _06707_);
  nand (_14569_, _14567_, _06707_);
  and (_14570_, _14569_, _14568_);
  and (_14571_, _14570_, _14560_);
  nor (_14572_, _14570_, _14560_);
  or (_14573_, _14572_, _14571_);
  nand (_14574_, _14573_, _06815_);
  nor (_14575_, _04483_, _06377_);
  and (_14576_, _11398_, _04483_);
  and (_14577_, _14576_, _11415_);
  nor (_14578_, _14577_, _14575_);
  nor (_14579_, _14578_, _02047_);
  nand (_14580_, _06821_, _03434_);
  or (_14581_, _13727_, _05166_);
  nand (_14582_, _06853_, _03434_);
  or (_14583_, _06855_, \oc8051_golden_model_1.ACC [3]);
  nand (_14584_, _06855_, \oc8051_golden_model_1.ACC [3]);
  nand (_14585_, _14584_, _14583_);
  nand (_14586_, _14585_, _06859_);
  and (_14587_, _14586_, _14582_);
  or (_14588_, _14587_, _02160_);
  nand (_14589_, _07056_, _02160_);
  and (_14590_, _14589_, _10299_);
  and (_14591_, _14590_, _14588_);
  or (_14592_, _14591_, _02079_);
  and (_14593_, _14592_, _03006_);
  and (_14594_, _14593_, _14581_);
  nor (_14595_, _11394_, _06736_);
  nor (_14596_, _14595_, _14539_);
  nor (_14597_, _14596_, _03006_);
  or (_14598_, _14597_, _06823_);
  or (_14599_, _14598_, _14594_);
  not (_14600_, \oc8051_golden_model_1.PSW [6]);
  nor (_14601_, _06824_, _14600_);
  nor (_14602_, _14601_, \oc8051_golden_model_1.ACC [3]);
  nor (_14603_, _14602_, _06825_);
  not (_14604_, _14603_);
  nand (_14605_, _14604_, _06823_);
  and (_14606_, _14605_, _14599_);
  or (_14607_, _14606_, _02057_);
  nor (_14608_, _14576_, _14575_);
  nand (_14609_, _14608_, _02057_);
  and (_14610_, _14609_, _02519_);
  and (_14611_, _14610_, _14607_);
  nor (_14612_, _14556_, _02519_);
  or (_14613_, _14612_, _06821_);
  or (_14614_, _14613_, _14611_);
  and (_14615_, _14614_, _14580_);
  or (_14616_, _14615_, _02582_);
  or (_14617_, _05166_, _06884_);
  and (_14618_, _14617_, _02549_);
  and (_14619_, _14618_, _14616_);
  nor (_14620_, _07056_, _02549_);
  or (_14621_, _14620_, _06888_);
  or (_14622_, _14621_, _14619_);
  nand (_14623_, _06888_, _04939_);
  and (_14624_, _14623_, _14622_);
  or (_14625_, _14624_, _02053_);
  and (_14626_, _11408_, _04483_);
  nor (_14627_, _14626_, _14575_);
  nand (_14628_, _14627_, _02053_);
  and (_14629_, _14628_, _02047_);
  and (_14630_, _14629_, _14625_);
  or (_14631_, _14630_, _14579_);
  and (_14632_, _14631_, _06181_);
  nor (_14633_, _06133_, _06131_);
  nor (_14634_, _14633_, _06134_);
  nand (_14635_, _14634_, _05474_);
  nand (_14636_, _14635_, _09041_);
  or (_14637_, _14636_, _14632_);
  and (_14638_, _03624_, \oc8051_golden_model_1.ACC [2]);
  nor (_14639_, _14299_, _14638_);
  nor (_14640_, _14534_, _14639_);
  and (_14641_, _14534_, _14639_);
  nor (_14642_, _14641_, _14640_);
  and (_14643_, _14642_, \oc8051_golden_model_1.PSW [7]);
  nor (_14644_, _14642_, \oc8051_golden_model_1.PSW [7]);
  nor (_14645_, _14644_, _14643_);
  and (_14646_, _14645_, _14305_);
  nor (_14647_, _14645_, _14305_);
  or (_14648_, _14647_, _14646_);
  nor (_14649_, _14648_, _02625_);
  or (_14650_, _14649_, _06816_);
  and (_14651_, _14650_, _14637_);
  nor (_14652_, _14648_, _02626_);
  or (_14653_, _14652_, _06815_);
  or (_14654_, _14653_, _14651_);
  and (_14655_, _14654_, _14574_);
  or (_14656_, _14655_, _02186_);
  nor (_14657_, _14332_, _07507_);
  nor (_14658_, _08849_, _14657_);
  and (_14659_, _08849_, _14657_);
  or (_14660_, _14659_, _14658_);
  not (_14661_, _14337_);
  and (_14662_, _14661_, _14660_);
  and (_14663_, _08876_, \oc8051_golden_model_1.PSW [7]);
  nor (_14664_, _14663_, _14662_);
  nand (_14665_, _14664_, _02186_);
  and (_14666_, _14665_, _06741_);
  and (_14667_, _14666_, _14656_);
  and (_14668_, _02452_, \oc8051_golden_model_1.ACC [2]);
  nor (_14669_, _14346_, _14668_);
  nor (_14670_, _08883_, _14669_);
  and (_14671_, _08883_, _14669_);
  nor (_14672_, _14671_, _14670_);
  not (_14673_, _14349_);
  nor (_14674_, _14673_, _14348_);
  not (_14675_, _14674_);
  or (_14676_, _14675_, _14672_);
  nand (_14677_, _14675_, _14672_);
  and (_14678_, _14677_, _14676_);
  nor (_14679_, _14678_, _06741_);
  or (_14680_, _14679_, _01876_);
  or (_14681_, _14680_, _14667_);
  nand (_14682_, _01983_, _01876_);
  and (_14683_, _14682_, _02043_);
  and (_14684_, _14683_, _14681_);
  nor (_14685_, _11433_, _07215_);
  nor (_14686_, _14685_, _14575_);
  nor (_14687_, _14686_, _02043_);
  or (_14688_, _14687_, _06188_);
  or (_14689_, _14688_, _14684_);
  and (_14690_, _14689_, _14557_);
  or (_14691_, _14690_, _02031_);
  and (_14692_, _05166_, _03841_);
  nor (_14693_, _14692_, _14539_);
  nand (_14694_, _14693_, _02031_);
  and (_14695_, _14694_, _02037_);
  and (_14696_, _14695_, _14691_);
  nor (_14697_, _11490_, _06736_);
  nor (_14698_, _14697_, _14539_);
  nor (_14699_, _14698_, _02037_);
  or (_14700_, _14699_, _06202_);
  or (_14701_, _14700_, _14696_);
  or (_14702_, _06344_, _06560_);
  and (_14703_, _14702_, _14701_);
  or (_14704_, _14703_, _01775_);
  and (_14705_, _14704_, _14554_);
  or (_14706_, _14705_, _01994_);
  and (_14707_, _03841_, _04719_);
  nor (_14708_, _14707_, _14539_);
  nand (_14709_, _14708_, _01994_);
  and (_14710_, _14709_, _07240_);
  and (_14711_, _14710_, _14706_);
  or (_14712_, _07240_, _01983_);
  nand (_14713_, _14712_, _14552_);
  or (_14714_, _14713_, _14711_);
  and (_14715_, _14714_, _14553_);
  or (_14716_, _14715_, _07258_);
  or (_14717_, _14087_, _14534_);
  and (_14718_, _14717_, _14095_);
  and (_14719_, _14718_, _14716_);
  and (_14720_, _07259_, _14534_);
  or (_14721_, _14720_, _07263_);
  or (_14722_, _14721_, _14719_);
  or (_14723_, _14563_, _07264_);
  and (_14724_, _14723_, _14722_);
  or (_14725_, _14724_, _02329_);
  or (_14726_, _11511_, _02330_);
  and (_14727_, _14726_, _07281_);
  and (_14728_, _14727_, _14725_);
  and (_14729_, _06734_, _08883_);
  or (_14730_, _14729_, _02210_);
  or (_14731_, _14730_, _14728_);
  and (_14732_, _14731_, _14546_);
  or (_14733_, _14732_, _02331_);
  not (_14734_, _02904_);
  and (_14735_, _13709_, _14734_);
  or (_14736_, _14539_, _03061_);
  and (_14737_, _14736_, _14735_);
  and (_14738_, _14737_, _14733_);
  and (_14739_, _02133_, _01727_);
  or (_14740_, _14739_, _02702_);
  or (_14741_, _14740_, _06627_);
  and (_14742_, _14741_, _13712_);
  or (_14743_, _14742_, _14738_);
  not (_14744_, _14740_);
  or (_14745_, _14744_, _06627_);
  and (_14746_, _14745_, _07305_);
  and (_14747_, _14746_, _14743_);
  and (_14748_, _07459_, _07304_);
  or (_14749_, _14748_, _02340_);
  or (_14750_, _14749_, _14747_);
  or (_14751_, _11509_, _02341_);
  and (_14752_, _14751_, _07313_);
  and (_14753_, _14752_, _14750_);
  and (_14754_, _07312_, _07544_);
  or (_14755_, _14754_, _14753_);
  and (_14756_, _14755_, _02208_);
  or (_14757_, _14708_, _11510_);
  nor (_14758_, _14757_, _02208_);
  or (_14759_, _14758_, _13948_);
  or (_14760_, _14759_, _14756_);
  and (_14761_, _14760_, _14543_);
  or (_14762_, _14761_, _10128_);
  nor (_14763_, _06629_, _02719_);
  or (_14764_, _14763_, _10129_);
  and (_14765_, _14764_, _14762_);
  nor (_14766_, _06629_, _07327_);
  or (_14767_, _14766_, _07331_);
  or (_14768_, _14767_, _14765_);
  nand (_14769_, _07457_, _07331_);
  and (_14770_, _14769_, _02337_);
  and (_14771_, _14770_, _14768_);
  nand (_14772_, _11510_, _07341_);
  and (_14773_, _14772_, _07340_);
  or (_14774_, _14773_, _14771_);
  nand (_14775_, _07338_, _07545_);
  and (_14776_, _14775_, _04953_);
  and (_14777_, _14776_, _14774_);
  or (_14778_, _14777_, _14542_);
  and (_14779_, _14778_, _06730_);
  and (_14780_, _06715_, _06693_);
  nor (_14781_, _14780_, _06716_);
  and (_14782_, _14781_, _07348_);
  or (_14783_, _14782_, _06654_);
  or (_14784_, _14783_, _14779_);
  and (_14785_, _07369_, _06978_);
  nor (_14786_, _14785_, _07370_);
  or (_14787_, _14786_, _07356_);
  and (_14788_, _14787_, _02346_);
  and (_14789_, _14788_, _14784_);
  and (_14790_, _07400_, _07162_);
  nor (_14791_, _14790_, _07401_);
  or (_14792_, _14791_, _07384_);
  and (_14793_, _14792_, _07386_);
  or (_14794_, _14793_, _14789_);
  and (_14795_, _07428_, _06774_);
  nor (_14796_, _14795_, _07429_);
  or (_14797_, _14796_, _07417_);
  and (_14798_, _14797_, _07416_);
  and (_14799_, _14798_, _14794_);
  nand (_14800_, _07415_, \oc8051_golden_model_1.ACC [2]);
  nand (_14801_, _14800_, _06614_);
  or (_14802_, _14801_, _14799_);
  and (_14803_, _14802_, _14538_);
  or (_14804_, _14803_, _06609_);
  nor (_14805_, _07472_, _14563_);
  and (_14806_, _07472_, _14563_);
  nor (_14807_, _14806_, _14805_);
  nand (_14808_, _14807_, _06609_);
  and (_14809_, _14808_, _02087_);
  and (_14810_, _14809_, _14804_);
  nor (_14811_, _07516_, _08849_);
  and (_14812_, _07516_, _08849_);
  nor (_14813_, _14812_, _14811_);
  and (_14814_, _14813_, _02085_);
  or (_14815_, _14814_, _07487_);
  or (_14816_, _14815_, _14810_);
  nor (_14817_, _07557_, _08883_);
  and (_14818_, _07557_, _08883_);
  nor (_14819_, _14818_, _14817_);
  nand (_14820_, _14819_, _07487_);
  and (_14821_, _14820_, _07534_);
  and (_14822_, _14821_, _14816_);
  and (_14823_, _07533_, \oc8051_golden_model_1.ACC [2]);
  or (_14824_, _14823_, _02366_);
  or (_14825_, _14824_, _14822_);
  nand (_14826_, _14596_, _02366_);
  and (_14827_, _14826_, _07576_);
  and (_14828_, _14827_, _14825_);
  nor (_14829_, _14506_, _06377_);
  or (_14830_, _14829_, _07583_);
  and (_14831_, _14830_, _07575_);
  or (_14832_, _14831_, _07580_);
  or (_14833_, _14832_, _14828_);
  nand (_14834_, _07580_, _06283_);
  and (_14835_, _14834_, _01698_);
  and (_14836_, _14835_, _14833_);
  nor (_14837_, _14627_, _01698_);
  or (_14838_, _14837_, _02081_);
  or (_14839_, _14838_, _14836_);
  and (_14840_, _11567_, _03841_);
  nor (_14841_, _14840_, _14539_);
  nand (_14842_, _14841_, _02081_);
  and (_14843_, _14842_, _07600_);
  and (_14844_, _14843_, _14839_);
  or (_14845_, _14523_, \oc8051_golden_model_1.ACC [3]);
  and (_14846_, _14845_, _07608_);
  and (_14847_, _14846_, _07599_);
  or (_14848_, _14847_, _07606_);
  or (_14849_, _14848_, _14844_);
  nand (_14850_, _07606_, _06283_);
  and (_14851_, _14850_, _39632_);
  and (_14852_, _14851_, _14849_);
  or (_14853_, _14852_, _14533_);
  and (_41628_, _14853_, _39026_);
  nor (_14854_, _39632_, _06283_);
  nand (_14855_, _07533_, _06377_);
  nand (_14856_, _07338_, _07542_);
  nand (_14857_, _13948_, _06624_);
  nor (_14858_, _07298_, _02702_);
  not (_14859_, _14858_);
  and (_14860_, _14859_, _06623_);
  nor (_14861_, _14550_, _10141_);
  not (_14862_, _14861_);
  nand (_14863_, _14862_, _06625_);
  nand (_14864_, _02825_, _01775_);
  nor (_14865_, _03841_, _06283_);
  nor (_14866_, _04372_, _06736_);
  nor (_14867_, _14866_, _14865_);
  nand (_14868_, _14867_, _06188_);
  nand (_14869_, _06821_, _04372_);
  nor (_14870_, _06825_, \oc8051_golden_model_1.ACC [4]);
  nor (_14871_, _14870_, _06831_);
  not (_14872_, _14871_);
  nand (_14873_, _14872_, _06823_);
  nor (_14874_, _07126_, _06847_);
  or (_14875_, _05303_, _06849_);
  nand (_14876_, _06853_, _04372_);
  or (_14877_, _06855_, \oc8051_golden_model_1.ACC [4]);
  nand (_14878_, _06855_, \oc8051_golden_model_1.ACC [4]);
  nand (_14879_, _14878_, _14877_);
  nand (_14880_, _14879_, _06859_);
  and (_14881_, _14880_, _14876_);
  and (_14882_, _14881_, _06847_);
  and (_14883_, _14882_, _14875_);
  or (_14884_, _14883_, _14874_);
  and (_14885_, _14884_, _06846_);
  nor (_14886_, _11611_, _06736_);
  nor (_14887_, _14886_, _14865_);
  nor (_14888_, _14887_, _03006_);
  or (_14889_, _14888_, _06823_);
  or (_14890_, _14889_, _14885_);
  and (_14891_, _14890_, _14873_);
  or (_14892_, _14891_, _02057_);
  nor (_14893_, _04483_, _06283_);
  and (_14894_, _11597_, _04483_);
  nor (_14895_, _14894_, _14893_);
  nand (_14896_, _14895_, _02057_);
  and (_14897_, _14896_, _02519_);
  and (_14898_, _14897_, _14892_);
  nor (_14899_, _14867_, _02519_);
  or (_14900_, _14899_, _06821_);
  or (_14901_, _14900_, _14898_);
  and (_14902_, _14901_, _14869_);
  or (_14903_, _14902_, _02582_);
  or (_14904_, _05303_, _06884_);
  and (_14905_, _14904_, _02549_);
  and (_14906_, _14905_, _14903_);
  nor (_14907_, _07126_, _02549_);
  or (_14908_, _14907_, _06888_);
  or (_14909_, _14908_, _14906_);
  nand (_14910_, _06888_, _01887_);
  and (_14911_, _14910_, _14909_);
  or (_14912_, _14911_, _02053_);
  and (_14913_, _11595_, _04483_);
  nor (_14914_, _14913_, _14893_);
  nand (_14915_, _14914_, _02053_);
  and (_14916_, _14915_, _02047_);
  and (_14917_, _14916_, _14912_);
  and (_14918_, _14894_, _11628_);
  nor (_14919_, _14918_, _14893_);
  nor (_14920_, _14919_, _02047_);
  or (_14921_, _14920_, _05474_);
  or (_14922_, _14921_, _14917_);
  nor (_14923_, _06136_, _06134_);
  nor (_14924_, _14923_, _06137_);
  or (_14925_, _14924_, _06181_);
  and (_14926_, _14925_, _14922_);
  or (_14927_, _14926_, _06817_);
  or (_14928_, _14646_, _14643_);
  nor (_14929_, _03434_, \oc8051_golden_model_1.ACC [3]);
  nand (_14930_, _03434_, \oc8051_golden_model_1.ACC [3]);
  and (_14931_, _14930_, _14639_);
  or (_14932_, _14931_, _14929_);
  nor (_14933_, _06625_, _14932_);
  and (_14934_, _06625_, _14932_);
  nor (_14935_, _14934_, _14933_);
  and (_14936_, _14935_, \oc8051_golden_model_1.PSW [7]);
  nor (_14937_, _14935_, \oc8051_golden_model_1.PSW [7]);
  nor (_14938_, _14937_, _14936_);
  and (_14939_, _14938_, _14928_);
  nor (_14940_, _14938_, _14928_);
  nor (_14941_, _14940_, _14939_);
  and (_14942_, _14941_, _06941_);
  or (_14943_, _14942_, _10153_);
  and (_14944_, _14943_, _14927_);
  not (_14945_, _14571_);
  and (_14946_, _14945_, _14568_);
  and (_14947_, _05166_, _06377_);
  or (_14948_, _05166_, _06377_);
  and (_14949_, _14948_, _14562_);
  or (_14950_, _14949_, _14947_);
  nor (_14951_, _07456_, _14950_);
  not (_14952_, _14951_);
  nand (_14953_, _07456_, _14950_);
  and (_14954_, _14953_, _14952_);
  nand (_14955_, _14954_, \oc8051_golden_model_1.PSW [7]);
  or (_14956_, _14954_, \oc8051_golden_model_1.PSW [7]);
  nand (_14957_, _14956_, _14955_);
  or (_14958_, _14957_, _14946_);
  and (_14959_, _14957_, _14946_);
  not (_14960_, _14959_);
  and (_14961_, _14960_, _14958_);
  and (_14962_, _14961_, _06815_);
  or (_14963_, _14962_, _02186_);
  or (_14964_, _14963_, _14944_);
  nor (_14965_, _14657_, _08847_);
  or (_14966_, _14965_, _08848_);
  and (_14967_, _07504_, _14966_);
  nor (_14968_, _07504_, _14966_);
  nor (_14969_, _14968_, _14967_);
  not (_14970_, _14663_);
  nor (_14971_, _14970_, _14969_);
  and (_14972_, _14970_, _14969_);
  nor (_14973_, _14972_, _14971_);
  nand (_14974_, _14973_, _02186_);
  and (_14975_, _14974_, _06741_);
  and (_14976_, _14975_, _14964_);
  nor (_14977_, _08921_, _06707_);
  nor (_14978_, _14669_, _08893_);
  nor (_14979_, _14978_, _08892_);
  nor (_14980_, _07543_, _14979_);
  and (_14981_, _07543_, _14979_);
  nor (_14982_, _14981_, _14980_);
  and (_14983_, _14982_, \oc8051_golden_model_1.PSW [7]);
  nor (_14984_, _14982_, \oc8051_golden_model_1.PSW [7]);
  nor (_14985_, _14984_, _14983_);
  and (_14986_, _14985_, _14977_);
  nor (_14987_, _14985_, _14977_);
  nor (_14988_, _14987_, _14986_);
  and (_14989_, _14988_, _06740_);
  or (_14990_, _14989_, _01876_);
  or (_14991_, _14990_, _14976_);
  nand (_14992_, _02825_, _01876_);
  and (_14993_, _14992_, _02043_);
  and (_14994_, _14993_, _14991_);
  nor (_14995_, _11646_, _07215_);
  nor (_14996_, _14995_, _14893_);
  nor (_14997_, _14996_, _02043_);
  or (_14998_, _14997_, _06188_);
  or (_14999_, _14998_, _14994_);
  and (_15000_, _14999_, _14868_);
  or (_15001_, _15000_, _02031_);
  and (_15002_, _05303_, _03841_);
  nor (_15003_, _15002_, _14865_);
  nand (_15004_, _15003_, _02031_);
  and (_15005_, _15004_, _02037_);
  and (_15006_, _15005_, _15001_);
  nor (_15007_, _11704_, _06736_);
  nor (_15008_, _15007_, _14865_);
  nor (_15009_, _15008_, _02037_);
  or (_15010_, _15009_, _06202_);
  or (_15011_, _15010_, _15006_);
  or (_15012_, _06292_, _06560_);
  and (_15013_, _15012_, _15011_);
  or (_15014_, _15013_, _01775_);
  nand (_15015_, _15014_, _14864_);
  and (_15016_, _15015_, _01995_);
  and (_15017_, _04831_, _03841_);
  nor (_15018_, _15017_, _14865_);
  and (_15019_, _15018_, _01994_);
  or (_15020_, _15019_, _07239_);
  or (_15021_, _15020_, _15016_);
  or (_15022_, _07240_, _02825_);
  and (_15023_, _15022_, _14548_);
  and (_15024_, _15023_, _15021_);
  nor (_15025_, _06625_, _14548_);
  or (_15026_, _15025_, _14862_);
  or (_15027_, _15026_, _15024_);
  and (_15028_, _15027_, _14863_);
  and (_15029_, _02691_, _01629_);
  or (_15030_, _15029_, _07258_);
  nor (_15031_, _15030_, _15028_);
  and (_15032_, _15030_, _06625_);
  or (_15033_, _15032_, _07259_);
  or (_15034_, _15033_, _15031_);
  nand (_15035_, _07259_, _06626_);
  and (_15036_, _15035_, _07264_);
  and (_15037_, _15036_, _15034_);
  and (_15038_, _07456_, _07263_);
  or (_15039_, _15038_, _02329_);
  or (_15040_, _15039_, _15037_);
  or (_15041_, _11588_, _02330_);
  and (_15042_, _15041_, _15040_);
  and (_15043_, _15042_, _07281_);
  and (_15044_, _06734_, _07543_);
  or (_15045_, _15044_, _02210_);
  or (_15046_, _15045_, _15043_);
  and (_15047_, _11592_, _03841_);
  nor (_15048_, _15047_, _14865_);
  nand (_15049_, _15048_, _02210_);
  and (_15050_, _15049_, _03061_);
  and (_15051_, _15050_, _15046_);
  and (_15052_, _14865_, _02331_);
  or (_15053_, _15052_, _07292_);
  or (_15054_, _15053_, _15051_);
  or (_15055_, _07295_, _06623_);
  and (_15056_, _15055_, _14858_);
  and (_15057_, _15056_, _15054_);
  or (_15058_, _15057_, _14860_);
  and (_15059_, _15058_, _07305_);
  and (_15060_, _07454_, _07304_);
  or (_15061_, _15060_, _02340_);
  or (_15062_, _15061_, _15059_);
  or (_15063_, _11586_, _02341_);
  and (_15064_, _15063_, _07313_);
  and (_15065_, _15064_, _15062_);
  and (_15066_, _07312_, _07541_);
  or (_15067_, _15066_, _15065_);
  and (_15068_, _15067_, _02208_);
  or (_15069_, _15018_, _11587_);
  nor (_15070_, _15069_, _02208_);
  or (_15071_, _15070_, _13948_);
  or (_15072_, _15071_, _15068_);
  and (_15073_, _15072_, _14857_);
  or (_15074_, _15073_, _10128_);
  nor (_15075_, _06624_, _02719_);
  or (_15076_, _15075_, _10129_);
  and (_15077_, _15076_, _15074_);
  nor (_15078_, _06624_, _07327_);
  or (_15079_, _15078_, _07331_);
  or (_15080_, _15079_, _15077_);
  nand (_15081_, _07455_, _07331_);
  and (_15082_, _15081_, _02337_);
  and (_15083_, _15082_, _15080_);
  nand (_15084_, _11587_, _07341_);
  and (_15085_, _15084_, _07340_);
  or (_15086_, _15085_, _15083_);
  and (_15087_, _15086_, _14856_);
  or (_15088_, _15087_, _02202_);
  nor (_15089_, _11590_, _06736_);
  nor (_15090_, _15089_, _14865_);
  nand (_15091_, _15090_, _02202_);
  and (_15092_, _15091_, _06730_);
  and (_15093_, _15092_, _15088_);
  and (_15094_, _06717_, _06684_);
  nor (_15095_, _15094_, _06718_);
  and (_15096_, _15095_, _07348_);
  or (_15097_, _15096_, _06654_);
  or (_15098_, _15097_, _15093_);
  and (_15099_, _07371_, _06969_);
  nor (_15100_, _15099_, _07372_);
  or (_15101_, _15100_, _07356_);
  and (_15102_, _15101_, _02346_);
  and (_15103_, _15102_, _15098_);
  and (_15104_, _07402_, _07155_);
  nor (_15105_, _15104_, _07403_);
  or (_15106_, _15105_, _07384_);
  and (_15107_, _15106_, _07386_);
  or (_15108_, _15107_, _15103_);
  and (_15109_, _07430_, _06768_);
  nor (_15110_, _15109_, _07431_);
  or (_15111_, _15110_, _07417_);
  and (_15112_, _15111_, _15108_);
  or (_15113_, _15112_, _07415_);
  nand (_15114_, _07415_, _06377_);
  and (_15115_, _15114_, _06614_);
  and (_15116_, _15115_, _15113_);
  and (_15117_, _06643_, _06626_);
  nor (_15118_, _15117_, _06644_);
  and (_15119_, _15118_, _09155_);
  or (_15120_, _15119_, _06609_);
  or (_15121_, _15120_, _15116_);
  nor (_15122_, _07474_, _07456_);
  nor (_15123_, _15122_, _07475_);
  or (_15124_, _15123_, _07448_);
  and (_15125_, _15124_, _15121_);
  or (_15126_, _15125_, _02085_);
  nor (_15127_, _07520_, _07505_);
  nor (_15128_, _15127_, _07521_);
  or (_15129_, _15128_, _02087_);
  and (_15130_, _15129_, _08458_);
  and (_15131_, _15130_, _15126_);
  nor (_15132_, _07559_, _07543_);
  nor (_15133_, _15132_, _07560_);
  and (_15134_, _15133_, _07487_);
  or (_15135_, _15134_, _07533_);
  or (_15136_, _15135_, _15131_);
  and (_15137_, _15136_, _14855_);
  or (_15138_, _15137_, _02366_);
  nand (_15139_, _14887_, _02366_);
  and (_15140_, _15139_, _07576_);
  and (_15141_, _15140_, _15138_);
  and (_15142_, _07583_, _06283_);
  nor (_15143_, _07583_, _06283_);
  nor (_15144_, _15143_, _15142_);
  not (_15145_, _15144_);
  nor (_15146_, _15145_, _07580_);
  nor (_15147_, _15146_, _07581_);
  or (_15148_, _15147_, _15141_);
  nand (_15149_, _07580_, _06277_);
  and (_15150_, _15149_, _01698_);
  and (_15151_, _15150_, _15148_);
  nor (_15152_, _14914_, _01698_);
  or (_15153_, _15152_, _02081_);
  or (_15154_, _15153_, _15151_);
  and (_15155_, _11771_, _03841_);
  nor (_15156_, _15155_, _14865_);
  nand (_15157_, _15156_, _02081_);
  and (_15158_, _15157_, _07600_);
  and (_15159_, _15158_, _15154_);
  and (_15160_, _07608_, _06283_);
  nor (_15161_, _15160_, _07609_);
  nor (_15162_, _15161_, _07606_);
  nor (_15163_, _15162_, _10751_);
  or (_15164_, _15163_, _15159_);
  nand (_15165_, _07606_, _06277_);
  and (_15166_, _15165_, _39632_);
  and (_15167_, _15166_, _15164_);
  or (_15168_, _15167_, _14854_);
  and (_41629_, _15168_, _39026_);
  nor (_15169_, _39632_, _06277_);
  nor (_15170_, _06622_, _06621_);
  not (_15171_, _15170_);
  nor (_15172_, _06645_, _15171_);
  and (_15173_, _06645_, _15171_);
  nor (_15174_, _15173_, _15172_);
  or (_15175_, _15174_, _06614_);
  and (_15176_, _06719_, _06676_);
  nor (_15177_, _15176_, _06720_);
  or (_15178_, _15177_, _06730_);
  not (_15179_, _10132_);
  nand (_15180_, _15179_, _06622_);
  or (_15181_, _07452_, _07305_);
  nor (_15182_, _03841_, _06277_);
  and (_15183_, _11915_, _03841_);
  nor (_15184_, _15183_, _15182_);
  nand (_15185_, _15184_, _02210_);
  not (_15186_, _02695_);
  nand (_15187_, _02410_, _01775_);
  nor (_15188_, _04057_, _06736_);
  nor (_15189_, _15188_, _15182_);
  nand (_15190_, _15189_, _06188_);
  nor (_15191_, _05303_, _06283_);
  nor (_15192_, _14951_, _15191_);
  nor (_15193_, _07453_, _07452_);
  not (_15194_, _15193_);
  nand (_15195_, _15194_, _15192_);
  or (_15196_, _15194_, _15192_);
  and (_15197_, _15196_, _15195_);
  or (_15198_, _15197_, _06707_);
  nand (_15199_, _15197_, _06707_);
  nand (_15200_, _15199_, _15198_);
  and (_15201_, _14958_, _14955_);
  or (_15202_, _15201_, _15200_);
  and (_15203_, _15201_, _15200_);
  not (_15204_, _15203_);
  and (_15205_, _15204_, _15202_);
  or (_15206_, _15205_, _06941_);
  nor (_15207_, _04483_, _06277_);
  and (_15208_, _11789_, _04483_);
  and (_15209_, _15208_, _11823_);
  nor (_15210_, _15209_, _15207_);
  nor (_15211_, _15210_, _02047_);
  nand (_15212_, _06821_, _04057_);
  and (_15213_, _08711_, _06833_);
  nor (_15214_, _08711_, _06833_);
  nor (_15215_, _15214_, _15213_);
  nand (_15216_, _15215_, _06823_);
  nor (_15217_, _07115_, _06847_);
  or (_15218_, _05258_, _06849_);
  nand (_15219_, _06853_, _04057_);
  or (_15220_, _06855_, \oc8051_golden_model_1.ACC [5]);
  nand (_15221_, _06855_, \oc8051_golden_model_1.ACC [5]);
  nand (_15222_, _15221_, _15220_);
  nand (_15223_, _15222_, _06859_);
  and (_15224_, _15223_, _15219_);
  and (_15225_, _15224_, _06847_);
  and (_15226_, _15225_, _15218_);
  or (_15227_, _15226_, _15217_);
  and (_15228_, _15227_, _06846_);
  nor (_15229_, _11804_, _06736_);
  nor (_15230_, _15229_, _15182_);
  nor (_15231_, _15230_, _03006_);
  or (_15232_, _15231_, _06823_);
  or (_15233_, _15232_, _15228_);
  and (_15234_, _15233_, _15216_);
  or (_15235_, _15234_, _02057_);
  nor (_15236_, _15208_, _15207_);
  nand (_15237_, _15236_, _02057_);
  and (_15238_, _15237_, _02519_);
  and (_15239_, _15238_, _15235_);
  nor (_15240_, _15189_, _02519_);
  or (_15241_, _15240_, _06821_);
  or (_15242_, _15241_, _15239_);
  and (_15243_, _15242_, _15212_);
  or (_15244_, _15243_, _02582_);
  or (_15245_, _05258_, _06884_);
  and (_15246_, _15245_, _02549_);
  and (_15247_, _15246_, _15244_);
  nor (_15248_, _07115_, _02549_);
  or (_15249_, _15248_, _06888_);
  or (_15250_, _15249_, _15247_);
  nand (_15251_, _06888_, _01804_);
  and (_15252_, _15251_, _15250_);
  or (_15253_, _15252_, _02053_);
  and (_15254_, _11816_, _04483_);
  nor (_15255_, _15254_, _15207_);
  nand (_15256_, _15255_, _02053_);
  and (_15257_, _15256_, _02047_);
  and (_15258_, _15257_, _15253_);
  or (_15259_, _15258_, _15211_);
  and (_15260_, _15259_, _06181_);
  nor (_15261_, _06139_, _06137_);
  nor (_15262_, _15261_, _06140_);
  nand (_15263_, _15262_, _05474_);
  nand (_15264_, _15263_, _09041_);
  or (_15265_, _15264_, _15260_);
  and (_15266_, _04372_, \oc8051_golden_model_1.ACC [4]);
  nor (_15267_, _14933_, _15266_);
  and (_15268_, _15171_, _15267_);
  nor (_15269_, _15171_, _15267_);
  nor (_15270_, _15269_, _15268_);
  nor (_15271_, _15270_, _06707_);
  and (_15272_, _15270_, _06707_);
  nor (_15273_, _15272_, _15271_);
  nor (_15274_, _14939_, _14936_);
  not (_15275_, _15274_);
  and (_15276_, _15275_, _15273_);
  nor (_15277_, _15275_, _15273_);
  nor (_15278_, _15277_, _15276_);
  and (_15279_, _15278_, _02626_);
  or (_15280_, _15279_, _06816_);
  and (_15281_, _15280_, _15265_);
  and (_15282_, _15278_, _02625_);
  or (_15283_, _15282_, _06815_);
  or (_15284_, _15283_, _15281_);
  and (_15285_, _15284_, _15206_);
  or (_15286_, _15285_, _02186_);
  nor (_15287_, _14967_, _07502_);
  nor (_15288_, _07500_, _15287_);
  and (_15289_, _07500_, _15287_);
  or (_15290_, _15289_, _15288_);
  not (_15291_, _14971_);
  nor (_15292_, _15291_, _15290_);
  and (_15293_, _15291_, _15290_);
  nor (_15294_, _15293_, _15292_);
  nand (_15295_, _15294_, _02186_);
  and (_15296_, _15295_, _06741_);
  and (_15297_, _15296_, _15286_);
  and (_15298_, _02825_, \oc8051_golden_model_1.ACC [4]);
  nor (_15299_, _14980_, _15298_);
  nor (_15300_, _07540_, _15299_);
  and (_15301_, _07540_, _15299_);
  or (_15302_, _15301_, _15300_);
  and (_15303_, _15302_, \oc8051_golden_model_1.PSW [7]);
  nor (_15304_, _15302_, \oc8051_golden_model_1.PSW [7]);
  nor (_15305_, _15304_, _15303_);
  nor (_15306_, _14986_, _14983_);
  not (_15307_, _15306_);
  and (_15308_, _15307_, _15305_);
  nor (_15309_, _15307_, _15305_);
  nor (_15310_, _15309_, _15308_);
  and (_15311_, _15310_, _06740_);
  or (_15312_, _15311_, _01876_);
  or (_15313_, _15312_, _15297_);
  nand (_15314_, _02410_, _01876_);
  and (_15315_, _15314_, _02043_);
  and (_15316_, _15315_, _15313_);
  nor (_15317_, _11841_, _07215_);
  nor (_15318_, _15317_, _15207_);
  nor (_15319_, _15318_, _02043_);
  or (_15320_, _15319_, _06188_);
  or (_15321_, _15320_, _15316_);
  and (_15322_, _15321_, _15190_);
  or (_15323_, _15322_, _02031_);
  and (_15324_, _05258_, _03841_);
  nor (_15325_, _15324_, _15182_);
  nand (_15326_, _15325_, _02031_);
  and (_15327_, _15326_, _02037_);
  and (_15328_, _15327_, _15323_);
  nor (_15329_, _11900_, _06736_);
  nor (_15330_, _15329_, _15182_);
  nor (_15331_, _15330_, _02037_);
  or (_15332_, _15331_, _06202_);
  or (_15333_, _15332_, _15328_);
  or (_15334_, _06262_, _06560_);
  and (_15335_, _15334_, _15333_);
  or (_15336_, _15335_, _01775_);
  nand (_15337_, _15336_, _15187_);
  and (_15338_, _15337_, _01995_);
  and (_15339_, _04827_, _03841_);
  nor (_15340_, _15339_, _15182_);
  and (_15341_, _15340_, _01994_);
  or (_15342_, _15341_, _07239_);
  or (_15343_, _15342_, _15338_);
  or (_15344_, _07240_, _02410_);
  and (_15345_, _15344_, _14548_);
  and (_15346_, _15345_, _15343_);
  nor (_15347_, _15170_, _14548_);
  or (_15348_, _15347_, _15346_);
  and (_15349_, _15348_, _15186_);
  nor (_15350_, _15170_, _15186_);
  and (_15351_, _02247_, _01721_);
  or (_15352_, _10142_, _15351_);
  or (_15353_, _15352_, _15030_);
  or (_15354_, _15353_, _15350_);
  nor (_15355_, _15354_, _15349_);
  and (_15356_, _15353_, _15170_);
  or (_15357_, _15356_, _07259_);
  or (_15358_, _15357_, _15355_);
  or (_15359_, _15170_, _14095_);
  and (_15360_, _15359_, _14398_);
  and (_15361_, _15360_, _15358_);
  or (_15362_, _15193_, _01598_);
  and (_15363_, _15362_, _07263_);
  or (_15364_, _15363_, _15361_);
  or (_15365_, _15193_, _14405_);
  and (_15366_, _15365_, _15364_);
  or (_15367_, _15366_, _02329_);
  or (_15368_, _11786_, _02330_);
  and (_15369_, _15368_, _07281_);
  and (_15370_, _15369_, _15367_);
  nor (_15371_, _07281_, _07540_);
  or (_15372_, _15371_, _02210_);
  or (_15373_, _15372_, _15370_);
  and (_15374_, _15373_, _15185_);
  or (_15375_, _15374_, _02331_);
  or (_15376_, _15182_, _03061_);
  and (_15377_, _15376_, _13709_);
  and (_15378_, _15377_, _15375_);
  nor (_15379_, _06621_, _02904_);
  nor (_15380_, _15379_, _14735_);
  or (_15381_, _15380_, _15378_);
  or (_15382_, _13710_, _06621_);
  and (_15383_, _15382_, _14744_);
  and (_15384_, _15383_, _15381_);
  and (_15385_, _14740_, _06621_);
  or (_15386_, _15385_, _07304_);
  or (_15387_, _15386_, _15384_);
  and (_15388_, _15387_, _15181_);
  or (_15389_, _15388_, _02340_);
  or (_15390_, _11784_, _02341_);
  and (_15391_, _15390_, _07313_);
  and (_15392_, _15391_, _15389_);
  and (_15393_, _07312_, _07538_);
  or (_15394_, _15393_, _15392_);
  and (_15395_, _15394_, _02208_);
  or (_15396_, _15340_, _11785_);
  nor (_15397_, _15396_, _02208_);
  or (_15398_, _15397_, _15179_);
  or (_15399_, _15398_, _15395_);
  and (_15400_, _15399_, _15180_);
  or (_15401_, _15400_, _07331_);
  nand (_15402_, _07453_, _07331_);
  and (_15403_, _15402_, _02337_);
  and (_15404_, _15403_, _15401_);
  nand (_15405_, _11785_, _07341_);
  and (_15406_, _15405_, _07340_);
  or (_15407_, _15406_, _15404_);
  nand (_15408_, _07338_, _07539_);
  and (_15409_, _15408_, _04953_);
  and (_15410_, _15409_, _15407_);
  nor (_15411_, _11913_, _06736_);
  nor (_15412_, _15411_, _15182_);
  nor (_15413_, _15412_, _04953_);
  or (_15414_, _15413_, _07348_);
  or (_15415_, _15414_, _15410_);
  and (_15416_, _15415_, _15178_);
  or (_15417_, _15416_, _06654_);
  and (_15418_, _07373_, _06967_);
  nor (_15419_, _15418_, _07374_);
  or (_15420_, _15419_, _07356_);
  and (_15421_, _15420_, _02346_);
  and (_15422_, _15421_, _15417_);
  and (_15423_, _07404_, _07153_);
  nor (_15424_, _15423_, _07405_);
  or (_15425_, _15424_, _07384_);
  and (_15426_, _15425_, _07386_);
  or (_15427_, _15426_, _15422_);
  and (_15428_, _07432_, _06763_);
  nor (_15429_, _15428_, _07433_);
  or (_15430_, _15429_, _07417_);
  and (_15431_, _15430_, _07416_);
  and (_15432_, _15431_, _15427_);
  and (_15433_, _07415_, \oc8051_golden_model_1.ACC [4]);
  or (_15434_, _15433_, _06610_);
  or (_15435_, _15434_, _06613_);
  or (_15436_, _15435_, _15432_);
  and (_15437_, _15436_, _15175_);
  or (_15438_, _15437_, _06609_);
  nor (_15439_, _07476_, _15194_);
  and (_15440_, _07476_, _15194_);
  nor (_15441_, _15440_, _15439_);
  or (_15442_, _15441_, _07448_);
  and (_15443_, _15442_, _02087_);
  and (_15444_, _15443_, _15438_);
  and (_15445_, _07522_, _07500_);
  nor (_15446_, _15445_, _07523_);
  and (_15447_, _15446_, _02085_);
  or (_15448_, _15447_, _07487_);
  or (_15449_, _15448_, _15444_);
  and (_15450_, _07561_, _07540_);
  nor (_15451_, _15450_, _07562_);
  or (_15452_, _15451_, _08458_);
  and (_15453_, _15452_, _07534_);
  and (_15454_, _15453_, _15449_);
  and (_15455_, _07533_, \oc8051_golden_model_1.ACC [4]);
  or (_15456_, _15455_, _02366_);
  or (_15457_, _15456_, _15454_);
  nand (_15458_, _15230_, _02366_);
  and (_15459_, _15458_, _07576_);
  and (_15460_, _15459_, _15457_);
  nor (_15461_, _15142_, _06277_);
  or (_15462_, _15461_, _07584_);
  and (_15463_, _15462_, _07575_);
  or (_15464_, _15463_, _07580_);
  or (_15465_, _15464_, _15460_);
  nand (_15466_, _07580_, _06231_);
  and (_15467_, _15466_, _01698_);
  and (_15468_, _15467_, _15465_);
  nor (_15469_, _15255_, _01698_);
  or (_15470_, _15469_, _02081_);
  or (_15471_, _15470_, _15468_);
  and (_15472_, _11974_, _03841_);
  nor (_15473_, _15472_, _15182_);
  nand (_15474_, _15473_, _02081_);
  and (_15475_, _15474_, _07600_);
  and (_15476_, _15475_, _15471_);
  nor (_15477_, _07609_, \oc8051_golden_model_1.ACC [5]);
  nor (_15478_, _15477_, _07610_);
  and (_15479_, _15478_, _07599_);
  or (_15480_, _15479_, _07606_);
  or (_15481_, _15480_, _15476_);
  nand (_15482_, _07606_, _06231_);
  and (_15483_, _15482_, _39632_);
  and (_15484_, _15483_, _15481_);
  or (_15485_, _15484_, _15169_);
  and (_41630_, _15485_, _39026_);
  nor (_15486_, _39632_, _06231_);
  nand (_15487_, _07338_, _07536_);
  nand (_15488_, _13948_, _06619_);
  or (_15489_, _13708_, _02904_);
  or (_15490_, _15489_, _14740_);
  and (_15491_, _15490_, _06618_);
  nand (_15492_, _02118_, _01775_);
  nor (_15493_, _03841_, _06231_);
  nor (_15494_, _03964_, _06736_);
  nor (_15495_, _15494_, _15493_);
  nand (_15496_, _15495_, _06188_);
  nor (_15497_, _15287_, _07498_);
  or (_15498_, _15497_, _07499_);
  and (_15499_, _15498_, _07496_);
  nor (_15500_, _15498_, _07496_);
  nor (_15501_, _15500_, _15499_);
  not (_15502_, _15292_);
  and (_15503_, _15502_, _15501_);
  nor (_15504_, _15502_, _15501_);
  nor (_15505_, _15504_, _15503_);
  nand (_15506_, _15505_, _02186_);
  and (_15507_, _15506_, _06741_);
  or (_15508_, _05258_, _06277_);
  and (_15509_, _05258_, _06277_);
  or (_15510_, _15192_, _15509_);
  and (_15511_, _15510_, _15508_);
  nor (_15512_, _15511_, _07451_);
  and (_15513_, _15511_, _07451_);
  nor (_15514_, _15513_, _15512_);
  and (_15515_, _15202_, _15198_);
  and (_15516_, _15515_, \oc8051_golden_model_1.PSW [7]);
  or (_15517_, _15516_, _15514_);
  nand (_15518_, _15516_, _15514_);
  and (_15519_, _15518_, _15517_);
  and (_15520_, _15519_, _06815_);
  nand (_15521_, _06821_, _03964_);
  not (_15522_, _06835_);
  nor (_15523_, _15214_, _15522_);
  and (_15524_, _08710_, _06836_);
  nor (_15525_, _15524_, _15523_);
  nand (_15526_, _15525_, _06823_);
  nor (_15527_, _07036_, _06847_);
  or (_15528_, _05029_, _06849_);
  nor (_15529_, _06852_, _03964_);
  and (_15530_, _06855_, _06231_);
  nor (_15531_, _06855_, _06231_);
  or (_15532_, _15531_, _02552_);
  or (_15533_, _15532_, _15530_);
  and (_15534_, _15533_, _06852_);
  or (_15535_, _15534_, _15529_);
  and (_15536_, _15535_, _06847_);
  and (_15537_, _15536_, _15528_);
  or (_15538_, _15537_, _15527_);
  and (_15539_, _15538_, _06846_);
  nor (_15540_, _11993_, _06736_);
  nor (_15541_, _15540_, _15493_);
  nor (_15542_, _15541_, _03006_);
  or (_15543_, _15542_, _06823_);
  or (_15544_, _15543_, _15539_);
  and (_15545_, _15544_, _15526_);
  or (_15546_, _15545_, _02057_);
  nor (_15547_, _04483_, _06231_);
  and (_15548_, _11990_, _04483_);
  nor (_15549_, _15548_, _15547_);
  nand (_15550_, _15549_, _02057_);
  and (_15551_, _15550_, _02519_);
  and (_15552_, _15551_, _15546_);
  nor (_15553_, _15495_, _02519_);
  or (_15554_, _15553_, _06821_);
  or (_15555_, _15554_, _15552_);
  and (_15556_, _15555_, _15521_);
  or (_15557_, _15556_, _02582_);
  or (_15558_, _05029_, _06884_);
  and (_15559_, _15558_, _02549_);
  and (_15560_, _15559_, _15557_);
  nor (_15561_, _07036_, _02549_);
  or (_15562_, _15561_, _06888_);
  or (_15563_, _15562_, _15560_);
  nand (_15564_, _06888_, _06383_);
  and (_15565_, _15564_, _15563_);
  or (_15566_, _15565_, _02053_);
  and (_15567_, _12017_, _04483_);
  nor (_15568_, _15567_, _15547_);
  nand (_15569_, _15568_, _02053_);
  and (_15570_, _15569_, _02047_);
  and (_15571_, _15570_, _15566_);
  and (_15572_, _15548_, _12024_);
  nor (_15573_, _15572_, _15547_);
  nor (_15574_, _15573_, _02047_);
  or (_15575_, _15574_, _05474_);
  or (_15576_, _15575_, _15571_);
  nor (_15577_, _06142_, _06140_);
  nor (_15578_, _15577_, _06143_);
  or (_15579_, _15578_, _06181_);
  and (_15580_, _15579_, _15576_);
  or (_15581_, _15580_, _06817_);
  nand (_15582_, _04057_, \oc8051_golden_model_1.ACC [5]);
  nor (_15583_, _04057_, \oc8051_golden_model_1.ACC [5]);
  or (_15584_, _15267_, _15583_);
  and (_15585_, _15584_, _15582_);
  nor (_15586_, _15585_, _06620_);
  and (_15587_, _15585_, _06620_);
  nor (_15588_, _15587_, _15586_);
  nor (_15589_, _15276_, _15271_);
  and (_15590_, _15589_, \oc8051_golden_model_1.PSW [7]);
  or (_15591_, _15590_, _15588_);
  nand (_15592_, _15590_, _15588_);
  and (_15593_, _15592_, _15591_);
  or (_15594_, _15593_, _06816_);
  and (_15595_, _15594_, _06941_);
  and (_15596_, _15595_, _15581_);
  or (_15597_, _15596_, _02186_);
  or (_15598_, _15597_, _15520_);
  and (_15599_, _15598_, _15507_);
  nor (_15600_, _15299_, _08905_);
  nor (_15601_, _15600_, _08904_);
  nor (_15602_, _15601_, _07537_);
  and (_15603_, _15601_, _07537_);
  nor (_15604_, _15603_, _15602_);
  nor (_15605_, _15308_, _15303_);
  and (_15606_, _15605_, \oc8051_golden_model_1.PSW [7]);
  nor (_15607_, _15606_, _15604_);
  and (_15608_, _15606_, _15604_);
  nor (_15609_, _15608_, _15607_);
  and (_15610_, _15609_, _06740_);
  or (_15611_, _15610_, _01876_);
  or (_15612_, _15611_, _15599_);
  nand (_15613_, _02118_, _01876_);
  and (_15614_, _15613_, _02043_);
  and (_15615_, _15614_, _15612_);
  nor (_15616_, _12042_, _07215_);
  nor (_15617_, _15616_, _15547_);
  nor (_15618_, _15617_, _02043_);
  or (_15619_, _15618_, _06188_);
  or (_15620_, _15619_, _15615_);
  and (_15621_, _15620_, _15496_);
  or (_15622_, _15621_, _02031_);
  and (_15623_, _05029_, _03841_);
  nor (_15624_, _15623_, _15493_);
  nand (_15625_, _15624_, _02031_);
  and (_15626_, _15625_, _02037_);
  and (_15627_, _15626_, _15622_);
  nor (_15628_, _12096_, _06736_);
  nor (_15629_, _15628_, _15493_);
  nor (_15630_, _15629_, _02037_);
  or (_15631_, _15630_, _06202_);
  or (_15632_, _15631_, _15627_);
  not (_15633_, _06232_);
  and (_15634_, _06236_, _15633_);
  or (_15635_, _15634_, _06560_);
  and (_15636_, _15635_, _15632_);
  or (_15637_, _15636_, _01775_);
  and (_15638_, _15637_, _15492_);
  or (_15639_, _15638_, _01994_);
  and (_15640_, _12103_, _03841_);
  nor (_15641_, _15640_, _15493_);
  nand (_15642_, _15641_, _01994_);
  and (_15643_, _15642_, _07240_);
  and (_15644_, _15643_, _15639_);
  nor (_15645_, _14547_, _02695_);
  or (_15646_, _07240_, _02118_);
  nand (_15647_, _15646_, _15645_);
  or (_15648_, _15647_, _15644_);
  nor (_15649_, _15645_, _06620_);
  nor (_15650_, _15649_, _15351_);
  and (_15651_, _15650_, _15648_);
  and (_15652_, _06620_, _15351_);
  or (_15653_, _15652_, _02693_);
  or (_15654_, _15653_, _15651_);
  or (_15655_, _06620_, _02694_);
  and (_15656_, _15655_, _15654_);
  and (_15657_, _02599_, _01721_);
  nor (_15658_, _10141_, _15657_);
  and (_15659_, _15658_, _14087_);
  and (_15660_, _15659_, _15656_);
  not (_15661_, _06620_);
  nor (_15662_, _15659_, _15661_);
  nor (_15663_, _15662_, _15660_);
  nand (_15664_, _15663_, _14095_);
  nand (_15665_, _07259_, _15661_);
  and (_15666_, _15665_, _07264_);
  and (_15667_, _15666_, _15664_);
  and (_15668_, _07451_, _07263_);
  or (_15669_, _15668_, _02329_);
  or (_15670_, _15669_, _15667_);
  or (_15671_, _12118_, _02330_);
  and (_15672_, _15671_, _15670_);
  and (_15673_, _15672_, _07281_);
  and (_15674_, _06734_, _07537_);
  or (_15676_, _15674_, _02210_);
  or (_15677_, _15676_, _15673_);
  and (_15678_, _12112_, _03841_);
  nor (_15679_, _15678_, _15493_);
  nand (_15680_, _15679_, _02210_);
  and (_15681_, _15680_, _03061_);
  and (_15682_, _15681_, _15677_);
  and (_15683_, _15493_, _02331_);
  or (_15684_, _15683_, _02895_);
  or (_15685_, _15684_, _15682_);
  not (_15687_, _13708_);
  and (_15688_, _15687_, _06618_);
  or (_15689_, _15688_, _13709_);
  and (_15690_, _15689_, _13710_);
  and (_15691_, _15690_, _15685_);
  or (_15692_, _15691_, _15491_);
  and (_15693_, _15692_, _07305_);
  and (_15694_, _07449_, _07304_);
  or (_15695_, _15694_, _02340_);
  or (_15696_, _15695_, _15693_);
  or (_15698_, _12116_, _02341_);
  and (_15699_, _15698_, _07313_);
  and (_15700_, _15699_, _15696_);
  and (_15701_, _07312_, _07535_);
  or (_15702_, _15701_, _15700_);
  and (_15703_, _15702_, _02208_);
  or (_15704_, _15641_, _12117_);
  nor (_15705_, _15704_, _02208_);
  or (_15706_, _15705_, _13948_);
  or (_15707_, _15706_, _15703_);
  and (_15709_, _15707_, _15488_);
  or (_15710_, _15709_, _10128_);
  nor (_15711_, _06619_, _02719_);
  or (_15712_, _15711_, _10129_);
  and (_15713_, _15712_, _15710_);
  nor (_15714_, _06619_, _07327_);
  or (_15715_, _15714_, _07331_);
  or (_15716_, _15715_, _15713_);
  nand (_15717_, _07450_, _07331_);
  and (_15718_, _15717_, _02337_);
  and (_15720_, _15718_, _15716_);
  nand (_15721_, _12117_, _07341_);
  and (_15722_, _15721_, _07340_);
  or (_15723_, _15722_, _15720_);
  and (_15724_, _15723_, _15487_);
  or (_15725_, _15724_, _02202_);
  nor (_15726_, _12110_, _06736_);
  nor (_15727_, _15726_, _15493_);
  nand (_15728_, _15727_, _02202_);
  and (_15729_, _15728_, _06730_);
  and (_15731_, _15729_, _15725_);
  and (_15732_, _06721_, _06669_);
  nor (_15733_, _15732_, _06722_);
  and (_15734_, _15733_, _07348_);
  or (_15735_, _15734_, _06654_);
  or (_15736_, _15735_, _15731_);
  and (_15737_, _07375_, _07358_);
  nor (_15738_, _15737_, _07376_);
  or (_15739_, _15738_, _07356_);
  and (_15740_, _15739_, _02346_);
  and (_15742_, _15740_, _15736_);
  and (_15743_, _07406_, _07388_);
  nor (_15744_, _15743_, _07407_);
  and (_15745_, _15744_, _02345_);
  or (_15746_, _15745_, _07384_);
  or (_15747_, _15746_, _15742_);
  and (_15748_, _07434_, _06757_);
  nor (_15749_, _15748_, _07435_);
  or (_15750_, _15749_, _07417_);
  and (_15751_, _15750_, _15747_);
  or (_15753_, _15751_, _07415_);
  nand (_15754_, _07415_, _06277_);
  and (_15755_, _15754_, _06614_);
  and (_15756_, _15755_, _15753_);
  nor (_15757_, _06647_, _06620_);
  nor (_15758_, _15757_, _06648_);
  and (_15759_, _15758_, _09155_);
  or (_15760_, _15759_, _06609_);
  or (_15761_, _15760_, _15756_);
  nor (_15762_, _07478_, _07451_);
  nor (_15764_, _15762_, _07479_);
  or (_15765_, _15764_, _07448_);
  and (_15766_, _15765_, _02087_);
  and (_15767_, _15766_, _15761_);
  and (_15768_, _07524_, _07496_);
  nor (_15769_, _15768_, _07525_);
  or (_15770_, _15769_, _07487_);
  and (_15771_, _15770_, _07489_);
  or (_15772_, _15771_, _15767_);
  nor (_15773_, _07563_, _07537_);
  nor (_15775_, _15773_, _07564_);
  or (_15776_, _15775_, _08458_);
  and (_15777_, _15776_, _07534_);
  and (_15778_, _15777_, _15772_);
  and (_15779_, _07533_, \oc8051_golden_model_1.ACC [5]);
  or (_15780_, _15779_, _02366_);
  or (_15781_, _15780_, _15778_);
  nand (_15782_, _15541_, _02366_);
  and (_15783_, _15782_, _07576_);
  and (_15784_, _15783_, _15781_);
  nor (_15786_, _07584_, _06231_);
  or (_15787_, _15786_, _07585_);
  and (_15788_, _15787_, _07575_);
  or (_15789_, _15788_, _07580_);
  or (_15790_, _15789_, _15784_);
  nand (_15791_, _07580_, _04939_);
  and (_15792_, _15791_, _01698_);
  and (_15793_, _15792_, _15790_);
  nor (_15794_, _15568_, _01698_);
  or (_15795_, _15794_, _02081_);
  or (_15797_, _15795_, _15793_);
  and (_15798_, _12178_, _03841_);
  nor (_15799_, _15798_, _15493_);
  nand (_15800_, _15799_, _02081_);
  and (_15801_, _15800_, _07600_);
  and (_15802_, _15801_, _15797_);
  nor (_15803_, _07610_, \oc8051_golden_model_1.ACC [6]);
  nor (_15804_, _15803_, _07611_);
  nor (_15805_, _15804_, _07606_);
  nor (_15806_, _15805_, _10751_);
  or (_15808_, _15806_, _15802_);
  nand (_15809_, _07606_, _04939_);
  and (_15810_, _15809_, _39632_);
  and (_15811_, _15810_, _15808_);
  or (_15812_, _15811_, _15486_);
  and (_41632_, _15812_, _39026_);
  not (_15813_, \oc8051_golden_model_1.DPL [0]);
  nor (_15814_, _39632_, _15813_);
  nor (_15815_, _04180_, _15813_);
  and (_15816_, _04180_, _03002_);
  or (_15818_, _15816_, _15815_);
  or (_15819_, _15818_, _05444_);
  and (_15820_, _03896_, \oc8051_golden_model_1.ACC [0]);
  or (_15821_, _15820_, _15815_);
  or (_15822_, _15821_, _02549_);
  nor (_15823_, _04257_, _07625_);
  or (_15824_, _15823_, _15815_);
  or (_15825_, _15824_, _03006_);
  and (_15826_, _15821_, _02062_);
  nor (_15827_, _02062_, _15813_);
  or (_15829_, _15827_, _02158_);
  or (_15830_, _15829_, _15826_);
  and (_15831_, _15830_, _02519_);
  and (_15832_, _15831_, _15825_);
  and (_15833_, _15818_, _02155_);
  or (_15834_, _15833_, _02153_);
  or (_15835_, _15834_, _15832_);
  and (_15836_, _15835_, _15822_);
  or (_15837_, _15836_, _07648_);
  nand (_15838_, _07648_, \oc8051_golden_model_1.DPL [0]);
  and (_15840_, _15838_, _07633_);
  and (_15841_, _15840_, _15837_);
  nor (_15842_, _02679_, _07633_);
  or (_15843_, _15842_, _06188_);
  or (_15844_, _15843_, _15841_);
  and (_15845_, _15844_, _15819_);
  or (_15846_, _15845_, _02031_);
  or (_15847_, _15815_, _02032_);
  and (_15848_, _05120_, _03896_);
  or (_15849_, _15848_, _15847_);
  and (_15851_, _15849_, _15846_);
  or (_15852_, _15851_, _01765_);
  nor (_15853_, _10898_, _07675_);
  or (_15854_, _15853_, _15815_);
  or (_15855_, _15854_, _02037_);
  and (_15856_, _15855_, _01995_);
  and (_15857_, _15856_, _15852_);
  and (_15858_, _03896_, _04837_);
  or (_15859_, _15858_, _15815_);
  and (_15860_, _15859_, _01994_);
  or (_15862_, _15860_, _02210_);
  or (_15863_, _15862_, _15857_);
  and (_15864_, _10914_, _03896_);
  or (_15865_, _15864_, _15815_);
  or (_15866_, _15865_, _03059_);
  and (_15867_, _15866_, _15863_);
  or (_15868_, _15867_, _02331_);
  and (_15869_, _10792_, _04180_);
  or (_15870_, _15815_, _03061_);
  or (_15871_, _15870_, _15869_);
  and (_15873_, _15871_, _02208_);
  and (_15874_, _15873_, _15868_);
  nand (_15875_, _15859_, _02206_);
  nor (_15876_, _15875_, _15823_);
  or (_15877_, _15876_, _15874_);
  and (_15878_, _15877_, _03065_);
  or (_15879_, _15815_, _04257_);
  and (_15880_, _15821_, _02342_);
  and (_15881_, _15880_, _15879_);
  or (_15882_, _15881_, _02202_);
  or (_15884_, _15882_, _15878_);
  nor (_15885_, _10913_, _07625_);
  or (_15886_, _15815_, _04953_);
  or (_15887_, _15886_, _15885_);
  and (_15888_, _15887_, _04958_);
  and (_15889_, _15888_, _15884_);
  not (_15890_, _02458_);
  nor (_15891_, _10789_, _07625_);
  or (_15892_, _15891_, _15815_);
  and (_15893_, _15892_, _02334_);
  or (_15895_, _15893_, _15890_);
  or (_15896_, _15895_, _15889_);
  or (_15897_, _15824_, _02458_);
  and (_15898_, _15897_, _39632_);
  and (_15899_, _15898_, _15896_);
  or (_15900_, _15899_, _15814_);
  and (_41633_, _15900_, _39026_);
  and (_15901_, _39633_, \oc8051_golden_model_1.DPL [1]);
  or (_15902_, _10988_, _07625_);
  or (_15903_, _04180_, \oc8051_golden_model_1.DPL [1]);
  and (_15905_, _15903_, _02206_);
  and (_15906_, _15905_, _15902_);
  or (_15907_, _11113_, _07625_);
  and (_15908_, _15903_, _02331_);
  and (_15909_, _15908_, _15907_);
  and (_15910_, _07625_, \oc8051_golden_model_1.DPL [1]);
  nor (_15911_, _07625_, _03161_);
  or (_15912_, _15911_, _15910_);
  or (_15913_, _15912_, _05444_);
  nor (_15914_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_15916_, _15914_, _07653_);
  and (_15917_, _15916_, _07648_);
  and (_15918_, _11001_, _04180_);
  not (_15919_, _15918_);
  and (_15920_, _15919_, _15903_);
  or (_15921_, _15920_, _03006_);
  nand (_15922_, _04180_, _01804_);
  and (_15923_, _15922_, _15903_);
  and (_15924_, _15923_, _02062_);
  and (_15925_, _02063_, \oc8051_golden_model_1.DPL [1]);
  or (_15927_, _15925_, _02158_);
  or (_15928_, _15927_, _15924_);
  and (_15929_, _15928_, _02519_);
  and (_15930_, _15929_, _15921_);
  and (_15931_, _15912_, _02155_);
  or (_15932_, _15931_, _02153_);
  or (_15933_, _15932_, _15930_);
  or (_15934_, _15923_, _02549_);
  and (_15935_, _15934_, _07649_);
  and (_15936_, _15935_, _15933_);
  or (_15938_, _15936_, _15917_);
  and (_15939_, _15938_, _07633_);
  nor (_15940_, _02893_, _07633_);
  or (_15941_, _15940_, _06188_);
  or (_15942_, _15941_, _15939_);
  and (_15943_, _15942_, _15913_);
  or (_15944_, _15943_, _02031_);
  and (_15945_, _05075_, _03896_);
  or (_15946_, _15910_, _02032_);
  or (_15947_, _15946_, _15945_);
  and (_15949_, _15947_, _02037_);
  and (_15950_, _15949_, _15944_);
  and (_15951_, _15903_, _01765_);
  nand (_15952_, _11096_, _04180_);
  and (_15953_, _15952_, _15951_);
  or (_15954_, _15953_, _15950_);
  and (_15955_, _15954_, _02212_);
  and (_15956_, _15903_, _01994_);
  nand (_15957_, _04180_, _02893_);
  and (_15958_, _15957_, _15956_);
  and (_15960_, _15903_, _02210_);
  or (_15961_, _10989_, _07625_);
  and (_15962_, _15961_, _15960_);
  or (_15963_, _15962_, _15958_);
  or (_15964_, _15963_, _15955_);
  and (_15965_, _15964_, _03061_);
  or (_15966_, _15965_, _15909_);
  and (_15967_, _15966_, _02208_);
  or (_15968_, _15967_, _15906_);
  and (_15969_, _15968_, _03065_);
  or (_15971_, _15910_, _04209_);
  and (_15972_, _15923_, _02342_);
  and (_15973_, _15972_, _15971_);
  or (_15974_, _15973_, _15969_);
  and (_15975_, _15974_, _02335_);
  or (_15976_, _15922_, _04209_);
  and (_15977_, _15903_, _02334_);
  and (_15978_, _15977_, _15976_);
  or (_15979_, _15978_, _02366_);
  or (_15980_, _15957_, _04209_);
  and (_15982_, _15903_, _02202_);
  and (_15983_, _15982_, _15980_);
  or (_15984_, _15983_, _15979_);
  or (_15985_, _15984_, _15975_);
  or (_15986_, _15920_, _02778_);
  and (_15987_, _15986_, _15985_);
  or (_15988_, _15987_, _02081_);
  or (_15989_, _15910_, _02082_);
  or (_15990_, _15989_, _15918_);
  and (_15991_, _15990_, _39632_);
  and (_15993_, _15991_, _15988_);
  or (_15994_, _15993_, _15901_);
  and (_41634_, _15994_, _39026_);
  not (_15995_, \oc8051_golden_model_1.DPL [2]);
  nor (_15996_, _39632_, _15995_);
  nor (_15997_, _04180_, _15995_);
  nor (_15998_, _11314_, _07625_);
  or (_15999_, _15998_, _15997_);
  and (_16000_, _15999_, _02334_);
  and (_16001_, _11315_, _04180_);
  or (_16003_, _16001_, _15997_);
  and (_16004_, _16003_, _02331_);
  nor (_16005_, _07625_, _03624_);
  or (_16006_, _16005_, _15997_);
  or (_16007_, _16006_, _05444_);
  or (_16008_, _16006_, _02519_);
  nor (_16009_, _11199_, _07625_);
  or (_16010_, _16009_, _15997_);
  and (_16011_, _16010_, _02158_);
  nor (_16012_, _02062_, _15995_);
  and (_16014_, _04180_, \oc8051_golden_model_1.ACC [2]);
  or (_16015_, _16014_, _15997_);
  and (_16016_, _16015_, _02062_);
  or (_16017_, _16016_, _16012_);
  and (_16018_, _16017_, _03006_);
  or (_16019_, _16018_, _02155_);
  or (_16020_, _16019_, _16011_);
  and (_16021_, _16020_, _16008_);
  or (_16022_, _16021_, _02153_);
  or (_16023_, _16015_, _02549_);
  and (_16024_, _16023_, _07649_);
  and (_16025_, _16024_, _16022_);
  nor (_16026_, _07653_, \oc8051_golden_model_1.DPL [2]);
  nor (_16027_, _16026_, _07654_);
  and (_16028_, _16027_, _07648_);
  or (_16029_, _16028_, _16025_);
  and (_16030_, _16029_, _07633_);
  nor (_16031_, _02494_, _07633_);
  or (_16032_, _16031_, _06188_);
  or (_16033_, _16032_, _16030_);
  and (_16036_, _16033_, _16007_);
  or (_16037_, _16036_, _02031_);
  or (_16038_, _15997_, _02032_);
  and (_16039_, _05211_, _03896_);
  or (_16040_, _16039_, _16038_);
  and (_16041_, _16040_, _02037_);
  and (_16042_, _16041_, _16037_);
  nor (_16043_, _11298_, _07675_);
  or (_16044_, _16043_, _15997_);
  and (_16045_, _16044_, _01765_);
  or (_16047_, _16045_, _16042_);
  or (_16048_, _16047_, _07629_);
  and (_16049_, _11189_, _04180_);
  or (_16050_, _15997_, _03059_);
  or (_16051_, _16050_, _16049_);
  and (_16052_, _03896_, _04866_);
  or (_16053_, _16052_, _15997_);
  or (_16054_, _16053_, _01995_);
  and (_16055_, _16054_, _03061_);
  and (_16056_, _16055_, _16051_);
  and (_16058_, _16056_, _16048_);
  or (_16059_, _16058_, _16004_);
  and (_16060_, _16059_, _02208_);
  or (_16061_, _15997_, _04309_);
  and (_16062_, _16053_, _02206_);
  and (_16063_, _16062_, _16061_);
  or (_16064_, _16063_, _16060_);
  and (_16065_, _16064_, _03065_);
  and (_16066_, _16015_, _02342_);
  and (_16067_, _16066_, _16061_);
  or (_16069_, _16067_, _02202_);
  or (_16070_, _16069_, _16065_);
  nor (_16071_, _11187_, _07625_);
  or (_16072_, _15997_, _04953_);
  or (_16073_, _16072_, _16071_);
  and (_16074_, _16073_, _04958_);
  and (_16075_, _16074_, _16070_);
  or (_16076_, _16075_, _16000_);
  and (_16077_, _16076_, _02778_);
  and (_16078_, _16010_, _02366_);
  or (_16080_, _16078_, _02081_);
  or (_16081_, _16080_, _16077_);
  and (_16082_, _11367_, _04180_);
  or (_16083_, _15997_, _02082_);
  or (_16084_, _16083_, _16082_);
  and (_16085_, _16084_, _39632_);
  and (_16086_, _16085_, _16081_);
  or (_16087_, _16086_, _15996_);
  and (_41636_, _16087_, _39026_);
  not (_16088_, \oc8051_golden_model_1.DPL [3]);
  nor (_16090_, _39632_, _16088_);
  nor (_16091_, _04180_, _16088_);
  nor (_16092_, _11510_, _07625_);
  or (_16093_, _16092_, _16091_);
  and (_16094_, _16093_, _02334_);
  and (_16095_, _11511_, _04180_);
  or (_16096_, _16095_, _16091_);
  and (_16097_, _16096_, _02331_);
  nor (_16098_, _07625_, _03434_);
  or (_16099_, _16098_, _16091_);
  or (_16101_, _16099_, _05444_);
  nor (_16102_, _11394_, _07625_);
  or (_16103_, _16102_, _16091_);
  or (_16104_, _16103_, _03006_);
  and (_16105_, _03896_, \oc8051_golden_model_1.ACC [3]);
  or (_16106_, _16105_, _16091_);
  and (_16107_, _16106_, _02062_);
  nor (_16108_, _02062_, _16088_);
  or (_16109_, _16108_, _02158_);
  or (_16110_, _16109_, _16107_);
  and (_16112_, _16110_, _02519_);
  and (_16113_, _16112_, _16104_);
  and (_16114_, _16099_, _02155_);
  or (_16115_, _16114_, _02153_);
  or (_16116_, _16115_, _16113_);
  or (_16117_, _16106_, _02549_);
  and (_16118_, _16117_, _07649_);
  and (_16119_, _16118_, _16116_);
  nor (_16120_, _07654_, \oc8051_golden_model_1.DPL [3]);
  nor (_16121_, _16120_, _07655_);
  and (_16123_, _16121_, _07648_);
  or (_16124_, _16123_, _16119_);
  and (_16125_, _16124_, _07633_);
  nor (_16126_, _02324_, _07633_);
  or (_16127_, _16126_, _06188_);
  or (_16128_, _16127_, _16125_);
  and (_16129_, _16128_, _16101_);
  or (_16130_, _16129_, _02031_);
  or (_16131_, _16091_, _02032_);
  and (_16132_, _05166_, _03896_);
  or (_16134_, _16132_, _16131_);
  and (_16135_, _16134_, _02037_);
  and (_16136_, _16135_, _16130_);
  nor (_16137_, _11490_, _07675_);
  or (_16138_, _16137_, _16091_);
  and (_16139_, _16138_, _01765_);
  or (_16140_, _16139_, _16136_);
  or (_16141_, _16140_, _07629_);
  and (_16142_, _11505_, _04180_);
  or (_16143_, _16091_, _03059_);
  or (_16145_, _16143_, _16142_);
  and (_16146_, _03896_, _04719_);
  or (_16147_, _16146_, _16091_);
  or (_16148_, _16147_, _01995_);
  and (_16149_, _16148_, _03061_);
  and (_16150_, _16149_, _16145_);
  and (_16151_, _16150_, _16141_);
  or (_16152_, _16151_, _16097_);
  and (_16153_, _16152_, _02208_);
  or (_16154_, _16091_, _04153_);
  and (_16156_, _16147_, _02206_);
  and (_16157_, _16156_, _16154_);
  or (_16158_, _16157_, _16153_);
  and (_16159_, _16158_, _03065_);
  and (_16160_, _16106_, _02342_);
  and (_16161_, _16160_, _16154_);
  or (_16162_, _16161_, _02202_);
  or (_16163_, _16162_, _16159_);
  nor (_16164_, _11503_, _07625_);
  or (_16165_, _16091_, _04953_);
  or (_16167_, _16165_, _16164_);
  and (_16168_, _16167_, _04958_);
  and (_16169_, _16168_, _16163_);
  or (_16170_, _16169_, _16094_);
  and (_16171_, _16170_, _02778_);
  and (_16172_, _16103_, _02366_);
  or (_16173_, _16172_, _02081_);
  or (_16174_, _16173_, _16171_);
  and (_16175_, _11567_, _04180_);
  or (_16176_, _16091_, _02082_);
  or (_16178_, _16176_, _16175_);
  and (_16179_, _16178_, _39632_);
  and (_16180_, _16179_, _16174_);
  or (_16181_, _16180_, _16090_);
  and (_41637_, _16181_, _39026_);
  not (_16182_, \oc8051_golden_model_1.DPL [4]);
  nor (_16183_, _39632_, _16182_);
  nor (_16184_, _04180_, _16182_);
  nor (_16185_, _11587_, _07625_);
  or (_16186_, _16185_, _16184_);
  and (_16188_, _16186_, _02334_);
  or (_16189_, _16184_, _04420_);
  and (_16190_, _04831_, _03896_);
  or (_16191_, _16190_, _16184_);
  and (_16192_, _16191_, _02206_);
  and (_16193_, _16192_, _16189_);
  and (_16194_, _11588_, _04180_);
  or (_16195_, _16194_, _16184_);
  and (_16196_, _16195_, _02331_);
  nor (_16197_, _11611_, _07625_);
  or (_16199_, _16197_, _16184_);
  or (_16200_, _16199_, _03006_);
  and (_16201_, _03896_, \oc8051_golden_model_1.ACC [4]);
  or (_16202_, _16201_, _16184_);
  and (_16203_, _16202_, _02062_);
  nor (_16204_, _02062_, _16182_);
  or (_16205_, _16204_, _02158_);
  or (_16206_, _16205_, _16203_);
  and (_16207_, _16206_, _02519_);
  and (_16208_, _16207_, _16200_);
  nor (_16210_, _04372_, _07625_);
  or (_16211_, _16210_, _16184_);
  and (_16212_, _16211_, _02155_);
  or (_16213_, _16212_, _02153_);
  or (_16214_, _16213_, _16208_);
  or (_16215_, _16202_, _02549_);
  and (_16216_, _16215_, _07649_);
  and (_16217_, _16216_, _16214_);
  nor (_16218_, _07655_, \oc8051_golden_model_1.DPL [4]);
  nor (_16219_, _16218_, _07656_);
  and (_16221_, _16219_, _07648_);
  or (_16222_, _16221_, _16217_);
  and (_16223_, _16222_, _07633_);
  nor (_16224_, _04784_, _07633_);
  or (_16225_, _16224_, _06188_);
  or (_16226_, _16225_, _16223_);
  or (_16227_, _16211_, _05444_);
  and (_16228_, _16227_, _16226_);
  or (_16229_, _16228_, _02031_);
  and (_16230_, _05303_, _03896_);
  or (_16232_, _16184_, _02032_);
  or (_16233_, _16232_, _16230_);
  and (_16234_, _16233_, _02037_);
  and (_16235_, _16234_, _16229_);
  nor (_16236_, _11704_, _07625_);
  or (_16237_, _16236_, _16184_);
  and (_16238_, _16237_, _01765_);
  or (_16239_, _16238_, _07629_);
  or (_16240_, _16239_, _16235_);
  and (_16241_, _11592_, _04180_);
  or (_16243_, _16184_, _03059_);
  or (_16244_, _16243_, _16241_);
  or (_16245_, _16191_, _01995_);
  and (_16246_, _16245_, _03061_);
  and (_16247_, _16246_, _16244_);
  and (_16248_, _16247_, _16240_);
  or (_16249_, _16248_, _16196_);
  and (_16250_, _16249_, _02208_);
  or (_16251_, _16250_, _16193_);
  and (_16252_, _16251_, _03065_);
  and (_16254_, _16202_, _02342_);
  and (_16255_, _16254_, _16189_);
  or (_16256_, _16255_, _02202_);
  or (_16257_, _16256_, _16252_);
  nor (_16258_, _11590_, _07625_);
  or (_16259_, _16184_, _04953_);
  or (_16260_, _16259_, _16258_);
  and (_16261_, _16260_, _04958_);
  and (_16262_, _16261_, _16257_);
  or (_16263_, _16262_, _16188_);
  and (_16265_, _16263_, _02778_);
  and (_16266_, _16199_, _02366_);
  or (_16267_, _16266_, _02081_);
  or (_16268_, _16267_, _16265_);
  and (_16269_, _11771_, _04180_);
  or (_16270_, _16184_, _02082_);
  or (_16271_, _16270_, _16269_);
  and (_16272_, _16271_, _39632_);
  and (_16273_, _16272_, _16268_);
  or (_16274_, _16273_, _16183_);
  and (_41638_, _16274_, _39026_);
  and (_16276_, _39633_, \oc8051_golden_model_1.DPL [5]);
  and (_16277_, _07625_, \oc8051_golden_model_1.DPL [5]);
  nor (_16278_, _11785_, _07625_);
  or (_16279_, _16278_, _16277_);
  and (_16280_, _16279_, _02334_);
  nor (_16281_, _04057_, _07625_);
  or (_16282_, _16281_, _16277_);
  or (_16283_, _16282_, _05444_);
  nor (_16284_, _11804_, _07625_);
  or (_16286_, _16284_, _16277_);
  or (_16287_, _16286_, _03006_);
  and (_16288_, _03896_, \oc8051_golden_model_1.ACC [5]);
  or (_16289_, _16288_, _16277_);
  and (_16290_, _16289_, _02062_);
  and (_16291_, _02063_, \oc8051_golden_model_1.DPL [5]);
  or (_16292_, _16291_, _02158_);
  or (_16293_, _16292_, _16290_);
  and (_16294_, _16293_, _02519_);
  and (_16295_, _16294_, _16287_);
  and (_16297_, _16282_, _02155_);
  or (_16298_, _16297_, _02153_);
  or (_16299_, _16298_, _16295_);
  or (_16300_, _16289_, _02549_);
  and (_16301_, _16300_, _07649_);
  and (_16302_, _16301_, _16299_);
  nor (_16303_, _07656_, \oc8051_golden_model_1.DPL [5]);
  nor (_16304_, _16303_, _07657_);
  and (_16305_, _16304_, _07648_);
  or (_16306_, _16305_, _16302_);
  and (_16308_, _16306_, _07633_);
  nor (_16309_, _04815_, _07633_);
  or (_16310_, _16309_, _06188_);
  or (_16311_, _16310_, _16308_);
  and (_16312_, _16311_, _16283_);
  or (_16313_, _16312_, _02031_);
  or (_16314_, _16277_, _02032_);
  and (_16315_, _05258_, _03896_);
  or (_16316_, _16315_, _16314_);
  and (_16317_, _16316_, _02037_);
  and (_16319_, _16317_, _16313_);
  nor (_16320_, _11900_, _07675_);
  or (_16321_, _16320_, _16277_);
  and (_16322_, _16321_, _01765_);
  or (_16323_, _16322_, _16319_);
  or (_16324_, _16323_, _07629_);
  and (_16325_, _11915_, _04180_);
  or (_16326_, _16277_, _03059_);
  or (_16327_, _16326_, _16325_);
  and (_16328_, _04827_, _03896_);
  or (_16330_, _16328_, _16277_);
  or (_16331_, _16330_, _01995_);
  and (_16332_, _16331_, _03061_);
  and (_16333_, _16332_, _16327_);
  and (_16334_, _16333_, _16324_);
  and (_16335_, _11786_, _04180_);
  or (_16336_, _16335_, _16277_);
  and (_16337_, _16336_, _02331_);
  or (_16338_, _16337_, _16334_);
  and (_16339_, _16338_, _02208_);
  or (_16341_, _16277_, _04104_);
  and (_16342_, _16330_, _02206_);
  and (_16343_, _16342_, _16341_);
  or (_16344_, _16343_, _16339_);
  and (_16345_, _16344_, _03065_);
  and (_16346_, _16289_, _02342_);
  and (_16347_, _16346_, _16341_);
  or (_16348_, _16347_, _02202_);
  or (_16349_, _16348_, _16345_);
  nor (_16350_, _11913_, _07625_);
  or (_16352_, _16277_, _04953_);
  or (_16353_, _16352_, _16350_);
  and (_16354_, _16353_, _04958_);
  and (_16355_, _16354_, _16349_);
  or (_16356_, _16355_, _16280_);
  and (_16357_, _16356_, _02778_);
  and (_16358_, _16286_, _02366_);
  or (_16359_, _16358_, _02081_);
  or (_16360_, _16359_, _16357_);
  and (_16361_, _11974_, _04180_);
  or (_16363_, _16277_, _02082_);
  or (_16364_, _16363_, _16361_);
  and (_16365_, _16364_, _39632_);
  and (_16366_, _16365_, _16360_);
  or (_16367_, _16366_, _16276_);
  and (_41639_, _16367_, _39026_);
  not (_16368_, \oc8051_golden_model_1.DPL [6]);
  nor (_16369_, _39632_, _16368_);
  nor (_16370_, _04180_, _16368_);
  nor (_16371_, _12117_, _07625_);
  or (_16373_, _16371_, _16370_);
  and (_16374_, _16373_, _02334_);
  nor (_16375_, _03964_, _07625_);
  or (_16376_, _16375_, _16370_);
  or (_16377_, _16376_, _05444_);
  nor (_16378_, _11993_, _07625_);
  or (_16379_, _16378_, _16370_);
  or (_16380_, _16379_, _03006_);
  and (_16381_, _03896_, \oc8051_golden_model_1.ACC [6]);
  or (_16382_, _16381_, _16370_);
  and (_16384_, _16382_, _02062_);
  nor (_16385_, _02062_, _16368_);
  or (_16386_, _16385_, _02158_);
  or (_16387_, _16386_, _16384_);
  and (_16388_, _16387_, _02519_);
  and (_16389_, _16388_, _16380_);
  and (_16390_, _16376_, _02155_);
  or (_16391_, _16390_, _02153_);
  or (_16392_, _16391_, _16389_);
  or (_16393_, _16382_, _02549_);
  and (_16395_, _16393_, _07649_);
  and (_16396_, _16395_, _16392_);
  nor (_16397_, _07657_, \oc8051_golden_model_1.DPL [6]);
  nor (_16398_, _16397_, _07658_);
  and (_16399_, _16398_, _07648_);
  or (_16400_, _16399_, _16396_);
  and (_16401_, _16400_, _07633_);
  nor (_16402_, _04752_, _07633_);
  or (_16403_, _16402_, _06188_);
  or (_16404_, _16403_, _16401_);
  and (_16406_, _16404_, _16377_);
  or (_16407_, _16406_, _02031_);
  or (_16408_, _16370_, _02032_);
  and (_16409_, _05029_, _03896_);
  or (_16410_, _16409_, _16408_);
  and (_16411_, _16410_, _02037_);
  and (_16412_, _16411_, _16407_);
  nor (_16413_, _12096_, _07675_);
  or (_16414_, _16413_, _16370_);
  and (_16415_, _16414_, _01765_);
  or (_16417_, _16415_, _16412_);
  or (_16418_, _16417_, _07629_);
  and (_16419_, _12112_, _04180_);
  or (_16420_, _16370_, _03059_);
  or (_16421_, _16420_, _16419_);
  and (_16422_, _12103_, _03896_);
  or (_16423_, _16422_, _16370_);
  or (_16424_, _16423_, _01995_);
  and (_16425_, _16424_, _03061_);
  and (_16426_, _16425_, _16421_);
  and (_16428_, _16426_, _16418_);
  and (_16429_, _12118_, _04180_);
  or (_16430_, _16429_, _16370_);
  and (_16431_, _16430_, _02331_);
  or (_16432_, _16431_, _16428_);
  and (_16433_, _16432_, _02208_);
  or (_16434_, _16370_, _04011_);
  and (_16435_, _16423_, _02206_);
  and (_16436_, _16435_, _16434_);
  or (_16437_, _16436_, _16433_);
  and (_16439_, _16437_, _03065_);
  and (_16440_, _16382_, _02342_);
  and (_16441_, _16440_, _16434_);
  or (_16442_, _16441_, _02202_);
  or (_16443_, _16442_, _16439_);
  nor (_16444_, _12110_, _07625_);
  or (_16445_, _16370_, _04953_);
  or (_16446_, _16445_, _16444_);
  and (_16447_, _16446_, _04958_);
  and (_16448_, _16447_, _16443_);
  or (_16450_, _16448_, _16374_);
  and (_16451_, _16450_, _02778_);
  and (_16452_, _16379_, _02366_);
  or (_16453_, _16452_, _02081_);
  or (_16454_, _16453_, _16451_);
  and (_16455_, _12178_, _04180_);
  or (_16456_, _16370_, _02082_);
  or (_16457_, _16456_, _16455_);
  and (_16458_, _16457_, _39632_);
  and (_16459_, _16458_, _16454_);
  or (_16461_, _16459_, _16369_);
  and (_41640_, _16461_, _39026_);
  not (_16462_, \oc8051_golden_model_1.DPH [0]);
  nor (_16463_, _39632_, _16462_);
  nor (_16464_, _04202_, _16462_);
  and (_16465_, _10792_, _04202_);
  or (_16466_, _16465_, _16464_);
  and (_16467_, _16466_, _02331_);
  and (_16468_, _04202_, _03002_);
  or (_16469_, _16468_, _16464_);
  or (_16471_, _16469_, _05444_);
  nor (_16472_, _07660_, \oc8051_golden_model_1.DPH [0]);
  nor (_16473_, _16472_, _07748_);
  and (_16474_, _16473_, _07648_);
  or (_16475_, _16469_, _02519_);
  nor (_16476_, _04257_, _07723_);
  or (_16477_, _16476_, _16464_);
  and (_16478_, _16477_, _02158_);
  nor (_16479_, _02062_, _16462_);
  and (_16480_, _03889_, \oc8051_golden_model_1.ACC [0]);
  or (_16482_, _16480_, _16464_);
  and (_16483_, _16482_, _02062_);
  or (_16484_, _16483_, _16479_);
  and (_16485_, _16484_, _03006_);
  or (_16486_, _16485_, _02155_);
  or (_16487_, _16486_, _16478_);
  and (_16488_, _16487_, _16475_);
  or (_16489_, _16488_, _02153_);
  or (_16490_, _16482_, _02549_);
  and (_16491_, _16490_, _07649_);
  and (_16493_, _16491_, _16489_);
  or (_16494_, _16493_, _16474_);
  and (_16495_, _16494_, _07633_);
  nor (_16496_, _07633_, _02027_);
  or (_16497_, _16496_, _06188_);
  or (_16498_, _16497_, _16495_);
  and (_16499_, _16498_, _16471_);
  or (_16500_, _16499_, _02031_);
  or (_16501_, _16464_, _02032_);
  and (_16502_, _05120_, _03889_);
  or (_16504_, _16502_, _16501_);
  and (_16505_, _16504_, _02037_);
  and (_16506_, _16505_, _16500_);
  nor (_16507_, _10898_, _07771_);
  or (_16508_, _16507_, _16464_);
  and (_16509_, _16508_, _01765_);
  or (_16510_, _16509_, _16506_);
  or (_16511_, _16510_, _07629_);
  and (_16512_, _10914_, _04202_);
  or (_16513_, _16464_, _03059_);
  or (_16515_, _16513_, _16512_);
  and (_16516_, _03889_, _04837_);
  or (_16517_, _16516_, _16464_);
  or (_16518_, _16517_, _01995_);
  and (_16519_, _16518_, _03061_);
  and (_16520_, _16519_, _16515_);
  and (_16521_, _16520_, _16511_);
  or (_16522_, _16521_, _16467_);
  and (_16523_, _16522_, _02208_);
  nand (_16524_, _16517_, _02206_);
  nor (_16526_, _16524_, _16476_);
  or (_16527_, _16526_, _16523_);
  and (_16528_, _16527_, _03065_);
  or (_16529_, _16464_, _04257_);
  and (_16530_, _16482_, _02342_);
  and (_16531_, _16530_, _16529_);
  or (_16532_, _16531_, _02202_);
  or (_16533_, _16532_, _16528_);
  nor (_16534_, _10913_, _07723_);
  or (_16535_, _16464_, _04953_);
  or (_16537_, _16535_, _16534_);
  and (_16538_, _16537_, _04958_);
  and (_16539_, _16538_, _16533_);
  nor (_16540_, _10789_, _07723_);
  or (_16541_, _16540_, _16464_);
  and (_16542_, _16541_, _02334_);
  or (_16543_, _16542_, _15890_);
  or (_16544_, _16543_, _16539_);
  or (_16545_, _16477_, _02458_);
  and (_16546_, _16545_, _39632_);
  and (_16548_, _16546_, _16544_);
  or (_16549_, _16548_, _16463_);
  and (_41642_, _16549_, _39026_);
  not (_16550_, \oc8051_golden_model_1.DPH [1]);
  nor (_16551_, _39632_, _16550_);
  or (_16552_, _10988_, _07723_);
  or (_16553_, _04202_, \oc8051_golden_model_1.DPH [1]);
  and (_16554_, _16553_, _02206_);
  and (_16555_, _16554_, _16552_);
  or (_16556_, _11113_, _07723_);
  and (_16558_, _16553_, _02331_);
  and (_16559_, _16558_, _16556_);
  nor (_16560_, _04202_, _16550_);
  nor (_16561_, _07723_, _03161_);
  or (_16562_, _16561_, _16560_);
  or (_16563_, _16562_, _05444_);
  or (_16564_, _07748_, \oc8051_golden_model_1.DPH [1]);
  and (_16565_, _16564_, _07749_);
  and (_16566_, _16565_, _07648_);
  and (_16567_, _11001_, _04202_);
  not (_16569_, _16567_);
  and (_16570_, _16569_, _16553_);
  or (_16571_, _16570_, _03006_);
  nand (_16572_, _04202_, _01804_);
  and (_16573_, _16572_, _16553_);
  and (_16574_, _16573_, _02062_);
  nor (_16575_, _02062_, _16550_);
  or (_16576_, _16575_, _02158_);
  or (_16577_, _16576_, _16574_);
  and (_16578_, _16577_, _02519_);
  and (_16580_, _16578_, _16571_);
  and (_16581_, _16562_, _02155_);
  or (_16582_, _16581_, _02153_);
  or (_16583_, _16582_, _16580_);
  or (_16584_, _16573_, _02549_);
  and (_16585_, _16584_, _07649_);
  and (_16586_, _16585_, _16583_);
  or (_16587_, _16586_, _16566_);
  and (_16588_, _16587_, _07633_);
  nor (_16589_, _02859_, _07633_);
  or (_16591_, _16589_, _06188_);
  or (_16592_, _16591_, _16588_);
  and (_16593_, _16592_, _16563_);
  or (_16594_, _16593_, _02031_);
  or (_16595_, _16560_, _02032_);
  and (_16596_, _05075_, _03889_);
  or (_16597_, _16596_, _16595_);
  and (_16598_, _16597_, _02037_);
  and (_16599_, _16598_, _16594_);
  and (_16600_, _16553_, _01765_);
  nand (_16602_, _11096_, _04202_);
  and (_16603_, _16602_, _16600_);
  or (_16604_, _16603_, _16599_);
  and (_16605_, _16604_, _02212_);
  or (_16606_, _10989_, _07723_);
  and (_16607_, _16606_, _02210_);
  nand (_16608_, _04202_, _02893_);
  and (_16609_, _16608_, _01994_);
  or (_16610_, _16609_, _16607_);
  and (_16611_, _16610_, _16553_);
  or (_16613_, _16611_, _16605_);
  and (_16614_, _16613_, _03061_);
  or (_16615_, _16614_, _16559_);
  and (_16616_, _16615_, _02208_);
  or (_16617_, _16616_, _16555_);
  and (_16618_, _16617_, _03065_);
  or (_16619_, _16560_, _04209_);
  and (_16620_, _16573_, _02342_);
  and (_16621_, _16620_, _16619_);
  or (_16622_, _16621_, _16618_);
  and (_16624_, _16622_, _02335_);
  or (_16625_, _16572_, _04209_);
  and (_16626_, _16553_, _02334_);
  and (_16627_, _16626_, _16625_);
  or (_16628_, _16627_, _02366_);
  or (_16629_, _16608_, _04209_);
  and (_16630_, _16553_, _02202_);
  and (_16631_, _16630_, _16629_);
  or (_16632_, _16631_, _16628_);
  or (_16633_, _16632_, _16624_);
  or (_16635_, _16570_, _02778_);
  and (_16636_, _16635_, _16633_);
  or (_16637_, _16636_, _02081_);
  or (_16638_, _16560_, _02082_);
  or (_16639_, _16638_, _16567_);
  and (_16640_, _16639_, _39632_);
  and (_16641_, _16640_, _16637_);
  or (_16642_, _16641_, _16551_);
  and (_41643_, _16642_, _39026_);
  nor (_16643_, _39632_, _07747_);
  nor (_16645_, _04202_, _07747_);
  nor (_16646_, _11314_, _07723_);
  or (_16647_, _16646_, _16645_);
  and (_16648_, _16647_, _02334_);
  or (_16649_, _16645_, _04309_);
  and (_16650_, _03889_, _04866_);
  or (_16651_, _16650_, _16645_);
  and (_16652_, _16651_, _02206_);
  and (_16653_, _16652_, _16649_);
  and (_16654_, _11315_, _04202_);
  or (_16655_, _16654_, _16645_);
  and (_16656_, _16655_, _02331_);
  nor (_16657_, _11298_, _07723_);
  or (_16658_, _16645_, _02037_);
  or (_16659_, _16658_, _16657_);
  nand (_16660_, _07749_, _07747_);
  nor (_16661_, _07750_, _07649_);
  and (_16662_, _16661_, _16660_);
  nor (_16663_, _11199_, _07723_);
  or (_16664_, _16663_, _16645_);
  or (_16667_, _16664_, _03006_);
  and (_16668_, _03889_, \oc8051_golden_model_1.ACC [2]);
  or (_16669_, _16668_, _16645_);
  and (_16670_, _16669_, _02062_);
  nor (_16671_, _02062_, _07747_);
  or (_16672_, _16671_, _02158_);
  or (_16673_, _16672_, _16670_);
  and (_16674_, _16673_, _02519_);
  and (_16675_, _16674_, _16667_);
  nor (_16676_, _07723_, _03624_);
  or (_16678_, _16676_, _16645_);
  and (_16679_, _16678_, _02155_);
  or (_16680_, _16679_, _02153_);
  or (_16681_, _16680_, _16675_);
  or (_16682_, _16669_, _02549_);
  and (_16683_, _16682_, _07649_);
  and (_16684_, _16683_, _16681_);
  or (_16685_, _16684_, _16662_);
  and (_16686_, _16685_, _07633_);
  nor (_16687_, _02452_, _07633_);
  or (_16689_, _16687_, _06188_);
  or (_16690_, _16689_, _16686_);
  or (_16691_, _16678_, _05444_);
  and (_16692_, _16691_, _02032_);
  and (_16693_, _16692_, _16690_);
  and (_16694_, _05211_, _03889_);
  or (_16695_, _16694_, _16645_);
  and (_16696_, _16695_, _02031_);
  or (_16697_, _16696_, _01765_);
  or (_16698_, _16697_, _16693_);
  and (_16700_, _16698_, _16659_);
  or (_16701_, _16700_, _07629_);
  and (_16702_, _11189_, _04202_);
  or (_16703_, _16645_, _03059_);
  or (_16704_, _16703_, _16702_);
  or (_16705_, _16651_, _01995_);
  and (_16706_, _16705_, _03061_);
  and (_16707_, _16706_, _16704_);
  and (_16708_, _16707_, _16701_);
  or (_16709_, _16708_, _16656_);
  and (_16711_, _16709_, _02208_);
  or (_16712_, _16711_, _16653_);
  and (_16713_, _16712_, _03065_);
  and (_16714_, _16669_, _02342_);
  and (_16715_, _16714_, _16649_);
  or (_16716_, _16715_, _02202_);
  or (_16717_, _16716_, _16713_);
  nor (_16718_, _11187_, _07723_);
  or (_16719_, _16645_, _04953_);
  or (_16720_, _16719_, _16718_);
  and (_16722_, _16720_, _04958_);
  and (_16723_, _16722_, _16717_);
  or (_16724_, _16723_, _16648_);
  and (_16725_, _16724_, _02778_);
  and (_16726_, _16664_, _02366_);
  or (_16727_, _16726_, _02081_);
  or (_16728_, _16727_, _16725_);
  and (_16729_, _11367_, _04202_);
  or (_16730_, _16645_, _02082_);
  or (_16731_, _16730_, _16729_);
  and (_16733_, _16731_, _39632_);
  and (_16734_, _16733_, _16728_);
  or (_16735_, _16734_, _16643_);
  and (_41644_, _16735_, _39026_);
  not (_16736_, \oc8051_golden_model_1.DPH [3]);
  nor (_16737_, _39632_, _16736_);
  nor (_16738_, _04202_, _16736_);
  nor (_16739_, _11510_, _07723_);
  or (_16740_, _16739_, _16738_);
  and (_16741_, _16740_, _02334_);
  and (_16743_, _11511_, _04202_);
  or (_16744_, _16743_, _16738_);
  and (_16745_, _16744_, _02331_);
  nor (_16746_, _07723_, _03434_);
  or (_16747_, _16746_, _16738_);
  or (_16748_, _16747_, _05444_);
  or (_16749_, _07750_, \oc8051_golden_model_1.DPH [3]);
  nor (_16750_, _07751_, _07649_);
  and (_16751_, _16750_, _16749_);
  nor (_16752_, _11394_, _07723_);
  or (_16754_, _16752_, _16738_);
  or (_16755_, _16754_, _03006_);
  and (_16756_, _03889_, \oc8051_golden_model_1.ACC [3]);
  or (_16757_, _16756_, _16738_);
  and (_16758_, _16757_, _02062_);
  nor (_16759_, _02062_, _16736_);
  or (_16760_, _16759_, _02158_);
  or (_16761_, _16760_, _16758_);
  and (_16762_, _16761_, _02519_);
  and (_16763_, _16762_, _16755_);
  and (_16765_, _16747_, _02155_);
  or (_16766_, _16765_, _02153_);
  or (_16767_, _16766_, _16763_);
  or (_16768_, _16757_, _02549_);
  and (_16769_, _16768_, _07649_);
  and (_16770_, _16769_, _16767_);
  or (_16771_, _16770_, _16751_);
  and (_16772_, _16771_, _07633_);
  nor (_16773_, _07633_, _01983_);
  or (_16774_, _16773_, _06188_);
  or (_16776_, _16774_, _16772_);
  and (_16777_, _16776_, _16748_);
  or (_16778_, _16777_, _02031_);
  or (_16779_, _16738_, _02032_);
  and (_16780_, _05166_, _03889_);
  or (_16781_, _16780_, _16779_);
  and (_16782_, _16781_, _02037_);
  and (_16783_, _16782_, _16778_);
  nor (_16784_, _11490_, _07771_);
  or (_16785_, _16784_, _16738_);
  and (_16787_, _16785_, _01765_);
  or (_16788_, _16787_, _16783_);
  or (_16789_, _16788_, _07629_);
  and (_16790_, _11505_, _04202_);
  or (_16791_, _16738_, _03059_);
  or (_16792_, _16791_, _16790_);
  and (_16793_, _03889_, _04719_);
  or (_16794_, _16793_, _16738_);
  or (_16795_, _16794_, _01995_);
  and (_16796_, _16795_, _03061_);
  and (_16798_, _16796_, _16792_);
  and (_16799_, _16798_, _16789_);
  or (_16800_, _16799_, _16745_);
  and (_16801_, _16800_, _02208_);
  or (_16802_, _16738_, _04153_);
  and (_16803_, _16794_, _02206_);
  and (_16804_, _16803_, _16802_);
  or (_16805_, _16804_, _16801_);
  and (_16806_, _16805_, _03065_);
  and (_16807_, _16757_, _02342_);
  and (_16809_, _16807_, _16802_);
  or (_16810_, _16809_, _02202_);
  or (_16811_, _16810_, _16806_);
  nor (_16812_, _11503_, _07723_);
  or (_16813_, _16738_, _04953_);
  or (_16814_, _16813_, _16812_);
  and (_16815_, _16814_, _04958_);
  and (_16816_, _16815_, _16811_);
  or (_16817_, _16816_, _16741_);
  and (_16818_, _16817_, _02778_);
  and (_16820_, _16754_, _02366_);
  or (_16821_, _16820_, _02081_);
  or (_16822_, _16821_, _16818_);
  and (_16823_, _11567_, _04202_);
  or (_16824_, _16738_, _02082_);
  or (_16825_, _16824_, _16823_);
  and (_16826_, _16825_, _39632_);
  and (_16827_, _16826_, _16822_);
  or (_16828_, _16827_, _16737_);
  and (_41645_, _16828_, _39026_);
  not (_16830_, \oc8051_golden_model_1.DPH [4]);
  nor (_16831_, _39632_, _16830_);
  nor (_16832_, _04202_, _16830_);
  nor (_16833_, _11587_, _07723_);
  or (_16834_, _16833_, _16832_);
  and (_16835_, _16834_, _02334_);
  and (_16836_, _11588_, _04202_);
  or (_16837_, _16836_, _16832_);
  and (_16838_, _16837_, _02331_);
  nor (_16839_, _11611_, _07723_);
  or (_16841_, _16839_, _16832_);
  or (_16842_, _16841_, _03006_);
  and (_16843_, _03889_, \oc8051_golden_model_1.ACC [4]);
  or (_16844_, _16843_, _16832_);
  and (_16845_, _16844_, _02062_);
  nor (_16846_, _02062_, _16830_);
  or (_16847_, _16846_, _02158_);
  or (_16848_, _16847_, _16845_);
  and (_16849_, _16848_, _02519_);
  and (_16850_, _16849_, _16842_);
  nor (_16852_, _04372_, _07723_);
  or (_16853_, _16852_, _16832_);
  and (_16854_, _16853_, _02155_);
  or (_16855_, _16854_, _02153_);
  or (_16856_, _16855_, _16850_);
  or (_16857_, _16844_, _02549_);
  and (_16858_, _16857_, _07649_);
  and (_16859_, _16858_, _16856_);
  or (_16860_, _07751_, \oc8051_golden_model_1.DPH [4]);
  nor (_16861_, _07752_, _07649_);
  and (_16863_, _16861_, _16860_);
  or (_16864_, _16863_, _16859_);
  and (_16865_, _16864_, _07633_);
  nor (_16866_, _02825_, _07633_);
  or (_16867_, _16866_, _06188_);
  or (_16868_, _16867_, _16865_);
  or (_16869_, _16853_, _05444_);
  and (_16870_, _16869_, _16868_);
  or (_16871_, _16870_, _02031_);
  and (_16872_, _05303_, _03889_);
  or (_16874_, _16832_, _02032_);
  or (_16875_, _16874_, _16872_);
  and (_16876_, _16875_, _02037_);
  and (_16877_, _16876_, _16871_);
  nor (_16878_, _11704_, _07723_);
  or (_16879_, _16878_, _16832_);
  and (_16880_, _16879_, _01765_);
  or (_16881_, _16880_, _07629_);
  or (_16882_, _16881_, _16877_);
  and (_16883_, _11592_, _04202_);
  or (_16885_, _16832_, _03059_);
  or (_16886_, _16885_, _16883_);
  and (_16887_, _04831_, _03889_);
  or (_16888_, _16887_, _16832_);
  or (_16889_, _16888_, _01995_);
  and (_16890_, _16889_, _03061_);
  and (_16891_, _16890_, _16886_);
  and (_16892_, _16891_, _16882_);
  or (_16893_, _16892_, _16838_);
  and (_16894_, _16893_, _02208_);
  or (_16896_, _16832_, _04420_);
  and (_16897_, _16888_, _02206_);
  and (_16898_, _16897_, _16896_);
  or (_16899_, _16898_, _16894_);
  and (_16900_, _16899_, _03065_);
  and (_16901_, _16844_, _02342_);
  and (_16902_, _16901_, _16896_);
  or (_16903_, _16902_, _02202_);
  or (_16904_, _16903_, _16900_);
  nor (_16905_, _11590_, _07723_);
  or (_16907_, _16832_, _04953_);
  or (_16908_, _16907_, _16905_);
  and (_16909_, _16908_, _04958_);
  and (_16910_, _16909_, _16904_);
  or (_16911_, _16910_, _16835_);
  and (_16912_, _16911_, _02778_);
  and (_16913_, _16841_, _02366_);
  or (_16914_, _16913_, _02081_);
  or (_16915_, _16914_, _16912_);
  and (_16916_, _11771_, _04202_);
  or (_16918_, _16832_, _02082_);
  or (_16919_, _16918_, _16916_);
  and (_16920_, _16919_, _39632_);
  and (_16921_, _16920_, _16915_);
  or (_16922_, _16921_, _16831_);
  and (_41646_, _16922_, _39026_);
  and (_16923_, _39633_, \oc8051_golden_model_1.DPH [5]);
  and (_16924_, _07723_, \oc8051_golden_model_1.DPH [5]);
  nor (_16925_, _11785_, _07723_);
  or (_16926_, _16925_, _16924_);
  and (_16928_, _16926_, _02334_);
  nor (_16929_, _04057_, _07723_);
  or (_16930_, _16929_, _16924_);
  or (_16931_, _16930_, _05444_);
  nor (_16932_, _11804_, _07723_);
  or (_16933_, _16932_, _16924_);
  or (_16934_, _16933_, _03006_);
  and (_16935_, _03889_, \oc8051_golden_model_1.ACC [5]);
  or (_16936_, _16935_, _16924_);
  and (_16937_, _16936_, _02062_);
  and (_16939_, _02063_, \oc8051_golden_model_1.DPH [5]);
  or (_16940_, _16939_, _02158_);
  or (_16941_, _16940_, _16937_);
  and (_16942_, _16941_, _02519_);
  and (_16943_, _16942_, _16934_);
  and (_16944_, _16930_, _02155_);
  or (_16945_, _16944_, _02153_);
  or (_16946_, _16945_, _16943_);
  or (_16947_, _16936_, _02549_);
  and (_16948_, _16947_, _07649_);
  and (_16950_, _16948_, _16946_);
  or (_16951_, _07752_, \oc8051_golden_model_1.DPH [5]);
  nor (_16952_, _07753_, _07649_);
  and (_16953_, _16952_, _16951_);
  or (_16954_, _16953_, _16950_);
  and (_16955_, _16954_, _07633_);
  nor (_16956_, _02410_, _07633_);
  or (_16957_, _16956_, _06188_);
  or (_16958_, _16957_, _16955_);
  and (_16959_, _16958_, _16931_);
  or (_16961_, _16959_, _02031_);
  or (_16962_, _16924_, _02032_);
  and (_16963_, _05258_, _03889_);
  or (_16964_, _16963_, _16962_);
  and (_16965_, _16964_, _02037_);
  and (_16966_, _16965_, _16961_);
  nor (_16967_, _11900_, _07771_);
  or (_16968_, _16967_, _16924_);
  and (_16969_, _16968_, _01765_);
  or (_16970_, _16969_, _16966_);
  or (_16972_, _16970_, _07629_);
  and (_16973_, _11915_, _04202_);
  or (_16974_, _16924_, _03059_);
  or (_16975_, _16974_, _16973_);
  and (_16976_, _04827_, _03889_);
  or (_16977_, _16976_, _16924_);
  or (_16978_, _16977_, _01995_);
  and (_16979_, _16978_, _03061_);
  and (_16980_, _16979_, _16975_);
  and (_16981_, _16980_, _16972_);
  and (_16983_, _11786_, _04202_);
  or (_16984_, _16983_, _16924_);
  and (_16985_, _16984_, _02331_);
  or (_16986_, _16985_, _16981_);
  and (_16987_, _16986_, _02208_);
  or (_16988_, _16924_, _04104_);
  and (_16989_, _16977_, _02206_);
  and (_16990_, _16989_, _16988_);
  or (_16991_, _16990_, _16987_);
  and (_16992_, _16991_, _03065_);
  and (_16994_, _16936_, _02342_);
  and (_16995_, _16994_, _16988_);
  or (_16996_, _16995_, _02202_);
  or (_16997_, _16996_, _16992_);
  nor (_16998_, _11913_, _07723_);
  or (_16999_, _16924_, _04953_);
  or (_17000_, _16999_, _16998_);
  and (_17001_, _17000_, _04958_);
  and (_17002_, _17001_, _16997_);
  or (_17003_, _17002_, _16928_);
  and (_17005_, _17003_, _02778_);
  and (_17006_, _16933_, _02366_);
  or (_17007_, _17006_, _02081_);
  or (_17008_, _17007_, _17005_);
  and (_17009_, _11974_, _04202_);
  or (_17010_, _16924_, _02082_);
  or (_17011_, _17010_, _17009_);
  and (_17012_, _17011_, _39632_);
  and (_17013_, _17012_, _17008_);
  or (_17014_, _17013_, _16923_);
  and (_41647_, _17014_, _39026_);
  not (_17016_, \oc8051_golden_model_1.DPH [6]);
  nor (_17017_, _39632_, _17016_);
  nor (_17018_, _04202_, _17016_);
  nor (_17019_, _12117_, _07723_);
  or (_17020_, _17019_, _17018_);
  and (_17021_, _17020_, _02334_);
  nor (_17022_, _03964_, _07723_);
  or (_17023_, _17022_, _17018_);
  or (_17024_, _17023_, _05444_);
  nor (_17026_, _11993_, _07723_);
  or (_17027_, _17026_, _17018_);
  or (_17028_, _17027_, _03006_);
  and (_17029_, _03889_, \oc8051_golden_model_1.ACC [6]);
  or (_17030_, _17029_, _17018_);
  and (_17031_, _17030_, _02062_);
  nor (_17032_, _02062_, _17016_);
  or (_17033_, _17032_, _02158_);
  or (_17034_, _17033_, _17031_);
  and (_17035_, _17034_, _02519_);
  and (_17036_, _17035_, _17028_);
  and (_17037_, _17023_, _02155_);
  or (_17038_, _17037_, _02153_);
  or (_17039_, _17038_, _17036_);
  or (_17040_, _17030_, _02549_);
  and (_17041_, _17040_, _07649_);
  and (_17042_, _17041_, _17039_);
  or (_17043_, _07753_, \oc8051_golden_model_1.DPH [6]);
  nor (_17044_, _07754_, _07649_);
  and (_17045_, _17044_, _17043_);
  or (_17048_, _17045_, _17042_);
  and (_17049_, _17048_, _07633_);
  nor (_17050_, _07633_, _02118_);
  or (_17051_, _17050_, _06188_);
  or (_17052_, _17051_, _17049_);
  and (_17053_, _17052_, _17024_);
  or (_17054_, _17053_, _02031_);
  or (_17055_, _17018_, _02032_);
  and (_17056_, _05029_, _03889_);
  or (_17057_, _17056_, _17055_);
  and (_17059_, _17057_, _02037_);
  and (_17060_, _17059_, _17054_);
  nor (_17061_, _12096_, _07771_);
  or (_17062_, _17061_, _17018_);
  and (_17063_, _17062_, _01765_);
  or (_17064_, _17063_, _17060_);
  or (_17065_, _17064_, _07629_);
  and (_17066_, _12112_, _04202_);
  or (_17067_, _17018_, _03059_);
  or (_17068_, _17067_, _17066_);
  and (_17070_, _12103_, _03889_);
  or (_17071_, _17070_, _17018_);
  or (_17072_, _17071_, _01995_);
  and (_17073_, _17072_, _03061_);
  and (_17074_, _17073_, _17068_);
  and (_17075_, _17074_, _17065_);
  and (_17076_, _12118_, _04202_);
  or (_17077_, _17076_, _17018_);
  and (_17078_, _17077_, _02331_);
  or (_17079_, _17078_, _17075_);
  and (_17081_, _17079_, _02208_);
  or (_17082_, _17018_, _04011_);
  and (_17083_, _17071_, _02206_);
  and (_17084_, _17083_, _17082_);
  or (_17085_, _17084_, _17081_);
  and (_17086_, _17085_, _03065_);
  and (_17087_, _17030_, _02342_);
  and (_17088_, _17087_, _17082_);
  or (_17089_, _17088_, _02202_);
  or (_17090_, _17089_, _17086_);
  nor (_17092_, _12110_, _07723_);
  or (_17093_, _17018_, _04953_);
  or (_17094_, _17093_, _17092_);
  and (_17095_, _17094_, _04958_);
  and (_17096_, _17095_, _17090_);
  or (_17097_, _17096_, _17021_);
  and (_17098_, _17097_, _02778_);
  and (_17099_, _17027_, _02366_);
  or (_17100_, _17099_, _02081_);
  or (_17101_, _17100_, _17098_);
  and (_17103_, _12178_, _04202_);
  or (_17104_, _17018_, _02082_);
  or (_17105_, _17104_, _17103_);
  and (_17106_, _17105_, _39632_);
  and (_17107_, _17106_, _17101_);
  or (_17108_, _17107_, _17017_);
  and (_41648_, _17108_, _39026_);
  not (_17109_, \oc8051_golden_model_1.IE [0]);
  nor (_17110_, _03813_, _17109_);
  and (_17111_, _10792_, _03813_);
  nor (_17113_, _17111_, _17110_);
  nor (_17114_, _17113_, _03061_);
  and (_17115_, _03813_, _04837_);
  nor (_17116_, _17115_, _17110_);
  and (_17117_, _17116_, _01994_);
  and (_17118_, _03813_, _03002_);
  nor (_17119_, _17118_, _17110_);
  and (_17120_, _17119_, _06188_);
  and (_17121_, _03813_, \oc8051_golden_model_1.ACC [0]);
  nor (_17122_, _17121_, _17110_);
  nor (_17124_, _17122_, _02063_);
  nor (_17125_, _02062_, _17109_);
  or (_17126_, _17125_, _17124_);
  and (_17127_, _17126_, _03006_);
  nor (_17128_, _04257_, _07818_);
  nor (_17129_, _17128_, _17110_);
  nor (_17130_, _17129_, _03006_);
  or (_17131_, _17130_, _17127_);
  and (_17132_, _17131_, _02058_);
  nor (_17133_, _04473_, _17109_);
  and (_17135_, _10814_, _04473_);
  nor (_17136_, _17135_, _17133_);
  nor (_17137_, _17136_, _02058_);
  nor (_17138_, _17137_, _17132_);
  nor (_17139_, _17138_, _02155_);
  nor (_17140_, _17119_, _02519_);
  or (_17141_, _17140_, _17139_);
  and (_17142_, _17141_, _02549_);
  nor (_17143_, _17122_, _02549_);
  or (_17144_, _17143_, _17142_);
  and (_17146_, _17144_, _02054_);
  and (_17147_, _17110_, _02053_);
  or (_17148_, _17147_, _17146_);
  and (_17149_, _17148_, _02047_);
  nor (_17150_, _17129_, _02047_);
  or (_17151_, _17150_, _17149_);
  and (_17152_, _17151_, _02043_);
  nor (_17153_, _10798_, _07855_);
  nor (_17154_, _17153_, _17133_);
  nor (_17155_, _17154_, _02043_);
  or (_17157_, _17155_, _06188_);
  nor (_17158_, _17157_, _17152_);
  nor (_17159_, _17158_, _17120_);
  nor (_17160_, _17159_, _02031_);
  and (_17161_, _05120_, _03813_);
  nor (_17162_, _17110_, _02032_);
  not (_17163_, _17162_);
  nor (_17164_, _17163_, _17161_);
  or (_17165_, _17164_, _01765_);
  nor (_17166_, _17165_, _17160_);
  nor (_17168_, _10898_, _07818_);
  nor (_17169_, _17168_, _17110_);
  nor (_17170_, _17169_, _02037_);
  or (_17171_, _17170_, _01994_);
  nor (_17172_, _17171_, _17166_);
  nor (_17173_, _17172_, _17117_);
  or (_17174_, _17173_, _02210_);
  and (_17175_, _10914_, _03813_);
  or (_17176_, _17175_, _17110_);
  or (_17177_, _17176_, _03059_);
  and (_17179_, _17177_, _03061_);
  and (_17180_, _17179_, _17174_);
  nor (_17181_, _17180_, _17114_);
  nor (_17182_, _17181_, _02206_);
  or (_17183_, _17116_, _02208_);
  nor (_17184_, _17183_, _17128_);
  nor (_17185_, _17184_, _17182_);
  nor (_17186_, _17185_, _02342_);
  nor (_17187_, _17110_, _04257_);
  or (_17188_, _17187_, _03065_);
  nor (_17190_, _17188_, _17122_);
  or (_17191_, _17190_, _02202_);
  nor (_17192_, _17191_, _17186_);
  nor (_17193_, _10913_, _07818_);
  or (_17194_, _17110_, _04953_);
  nor (_17195_, _17194_, _17193_);
  or (_17196_, _17195_, _02334_);
  nor (_17197_, _17196_, _17192_);
  nor (_17198_, _10789_, _07818_);
  nor (_17199_, _17198_, _17110_);
  nor (_17201_, _17199_, _04958_);
  or (_17202_, _17201_, _17197_);
  and (_17203_, _17202_, _02778_);
  nor (_17204_, _17129_, _02778_);
  or (_17205_, _17204_, _17203_);
  and (_17206_, _17205_, _01698_);
  and (_17207_, _17110_, _01697_);
  or (_17208_, _17207_, _17206_);
  and (_17209_, _17208_, _02082_);
  nor (_17210_, _17129_, _02082_);
  or (_17212_, _17210_, _17209_);
  or (_17213_, _17212_, _39633_);
  or (_17214_, _39632_, \oc8051_golden_model_1.IE [0]);
  and (_17215_, _17214_, _39026_);
  and (_41650_, _17215_, _17213_);
  not (_17216_, _02335_);
  not (_17217_, \oc8051_golden_model_1.IE [1]);
  nor (_17218_, _03813_, _17217_);
  and (_17219_, _05075_, _03813_);
  or (_17220_, _17219_, _17218_);
  and (_17222_, _17220_, _02031_);
  nor (_17223_, _03813_, \oc8051_golden_model_1.IE [1]);
  and (_17224_, _03813_, _01804_);
  nor (_17225_, _17224_, _17223_);
  and (_17226_, _17225_, _02062_);
  nor (_17227_, _02062_, _17217_);
  or (_17228_, _17227_, _17226_);
  and (_17229_, _17228_, _03006_);
  and (_17230_, _11001_, _03813_);
  nor (_17231_, _17230_, _17223_);
  and (_17233_, _17231_, _02158_);
  or (_17234_, _17233_, _17229_);
  and (_17235_, _17234_, _02058_);
  nor (_17236_, _04473_, _17217_);
  and (_17237_, _11005_, _04473_);
  nor (_17238_, _17237_, _17236_);
  nor (_17239_, _17238_, _02058_);
  or (_17240_, _17239_, _17235_);
  and (_17241_, _17240_, _02519_);
  nor (_17242_, _07818_, _03161_);
  nor (_17244_, _17242_, _17218_);
  nor (_17245_, _17244_, _02519_);
  or (_17246_, _17245_, _17241_);
  nor (_17247_, _17246_, _02153_);
  nor (_17248_, _17225_, _02549_);
  or (_17249_, _17248_, _02053_);
  nor (_17250_, _17249_, _17247_);
  and (_17251_, _10992_, _04473_);
  nor (_17252_, _17251_, _17236_);
  nor (_17253_, _17252_, _02054_);
  or (_17255_, _17253_, _17250_);
  and (_17256_, _17255_, _02047_);
  nor (_17257_, _17236_, _11020_);
  nor (_17258_, _17257_, _17238_);
  and (_17259_, _17258_, _02046_);
  or (_17260_, _17259_, _17256_);
  and (_17261_, _17260_, _02043_);
  nor (_17262_, _11038_, _07855_);
  nor (_17263_, _17262_, _17236_);
  nor (_17264_, _17263_, _02043_);
  nor (_17266_, _17264_, _06188_);
  not (_17267_, _17266_);
  nor (_17268_, _17267_, _17261_);
  and (_17269_, _17244_, _06188_);
  or (_17270_, _17269_, _02031_);
  nor (_17271_, _17270_, _17268_);
  or (_17272_, _17271_, _17222_);
  and (_17273_, _17272_, _02037_);
  nor (_17274_, _11096_, _07818_);
  nor (_17275_, _17274_, _17218_);
  nor (_17277_, _17275_, _02037_);
  nor (_17278_, _17277_, _17273_);
  nor (_17279_, _17278_, _07629_);
  not (_17280_, _17223_);
  nor (_17281_, _10989_, _07818_);
  nor (_17282_, _17281_, _03059_);
  and (_17283_, _03813_, _02893_);
  nor (_17284_, _17283_, _01995_);
  or (_17285_, _17284_, _17282_);
  and (_17286_, _17285_, _17280_);
  nor (_17288_, _17286_, _17279_);
  nor (_17289_, _17288_, _02331_);
  nor (_17290_, _11113_, _07818_);
  nor (_17291_, _17290_, _03061_);
  and (_17292_, _17291_, _17280_);
  nor (_17293_, _17292_, _17289_);
  nor (_17294_, _17293_, _02206_);
  nor (_17295_, _10988_, _07818_);
  nor (_17296_, _17295_, _02208_);
  and (_17297_, _17296_, _17280_);
  nor (_17299_, _17297_, _17294_);
  nor (_17300_, _17299_, _02342_);
  nor (_17301_, _17218_, _04209_);
  nor (_17302_, _17301_, _03065_);
  and (_17303_, _17302_, _17225_);
  nor (_17304_, _17303_, _17300_);
  or (_17305_, _17304_, _17216_);
  nand (_17306_, _17224_, _04208_);
  nor (_17307_, _17223_, _04958_);
  and (_17308_, _17307_, _17306_);
  nor (_17310_, _17308_, _02366_);
  and (_17311_, _17283_, _04208_);
  or (_17312_, _17223_, _04953_);
  or (_17313_, _17312_, _17311_);
  and (_17314_, _17313_, _17310_);
  and (_17315_, _17314_, _17305_);
  nor (_17316_, _17231_, _02778_);
  or (_17317_, _17316_, _01697_);
  nor (_17318_, _17317_, _17315_);
  nor (_17319_, _17252_, _01698_);
  or (_17321_, _17319_, _02081_);
  nor (_17322_, _17321_, _17318_);
  nor (_17323_, _17230_, _17218_);
  and (_17324_, _17323_, _02081_);
  nor (_17325_, _17324_, _17322_);
  or (_17326_, _17325_, _39633_);
  or (_17327_, _39632_, \oc8051_golden_model_1.IE [1]);
  and (_17328_, _17327_, _39026_);
  and (_41651_, _17328_, _17326_);
  not (_17329_, \oc8051_golden_model_1.IE [2]);
  nor (_17331_, _03813_, _17329_);
  and (_17332_, _03813_, _04866_);
  nor (_17333_, _17332_, _17331_);
  and (_17334_, _17333_, _01994_);
  nor (_17335_, _07818_, _03624_);
  nor (_17336_, _17335_, _17331_);
  and (_17337_, _17336_, _06188_);
  and (_17338_, _03813_, \oc8051_golden_model_1.ACC [2]);
  nor (_17339_, _17338_, _17331_);
  nor (_17340_, _17339_, _02063_);
  nor (_17342_, _02062_, _17329_);
  or (_17343_, _17342_, _17340_);
  and (_17344_, _17343_, _03006_);
  nor (_17345_, _11199_, _07818_);
  nor (_17346_, _17345_, _17331_);
  nor (_17347_, _17346_, _03006_);
  or (_17348_, _17347_, _17344_);
  and (_17349_, _17348_, _02058_);
  nor (_17350_, _04473_, _17329_);
  and (_17351_, _11194_, _04473_);
  nor (_17353_, _17351_, _17350_);
  nor (_17354_, _17353_, _02058_);
  or (_17355_, _17354_, _02155_);
  or (_17356_, _17355_, _17349_);
  nand (_17357_, _17336_, _02155_);
  and (_17358_, _17357_, _17356_);
  and (_17359_, _17358_, _02549_);
  nor (_17360_, _17339_, _02549_);
  or (_17361_, _17360_, _17359_);
  and (_17362_, _17361_, _02054_);
  and (_17363_, _11192_, _04473_);
  nor (_17364_, _17363_, _17350_);
  nor (_17365_, _17364_, _02054_);
  or (_17366_, _17365_, _17362_);
  and (_17367_, _17366_, _02047_);
  nor (_17368_, _17350_, _11223_);
  nor (_17369_, _17368_, _17353_);
  and (_17370_, _17369_, _02046_);
  or (_17371_, _17370_, _17367_);
  and (_17372_, _17371_, _02043_);
  nor (_17374_, _11241_, _07855_);
  nor (_17375_, _17374_, _17350_);
  nor (_17376_, _17375_, _02043_);
  nor (_17377_, _17376_, _06188_);
  not (_17378_, _17377_);
  nor (_17379_, _17378_, _17372_);
  nor (_17380_, _17379_, _17337_);
  nor (_17381_, _17380_, _02031_);
  and (_17382_, _05211_, _03813_);
  nor (_17383_, _17331_, _02032_);
  not (_17385_, _17383_);
  nor (_17386_, _17385_, _17382_);
  or (_17387_, _17386_, _01765_);
  nor (_17388_, _17387_, _17381_);
  nor (_17389_, _11298_, _07818_);
  nor (_17390_, _17331_, _17389_);
  nor (_17391_, _17390_, _02037_);
  or (_17392_, _17391_, _01994_);
  nor (_17393_, _17392_, _17388_);
  nor (_17394_, _17393_, _17334_);
  or (_17396_, _17394_, _02210_);
  and (_17397_, _11189_, _03813_);
  or (_17398_, _17397_, _17331_);
  or (_17399_, _17398_, _03059_);
  and (_17400_, _17399_, _03061_);
  and (_17401_, _17400_, _17396_);
  and (_17402_, _11315_, _03813_);
  nor (_17403_, _17402_, _17331_);
  nor (_17404_, _17403_, _03061_);
  nor (_17405_, _17404_, _17401_);
  nor (_17407_, _17405_, _02206_);
  nor (_17408_, _17331_, _04309_);
  not (_17409_, _17408_);
  nor (_17410_, _17333_, _02208_);
  and (_17411_, _17410_, _17409_);
  nor (_17412_, _17411_, _17407_);
  nor (_17413_, _17412_, _02342_);
  or (_17414_, _17408_, _03065_);
  nor (_17415_, _17414_, _17339_);
  or (_17416_, _17415_, _02202_);
  nor (_17418_, _17416_, _17413_);
  nor (_17419_, _11187_, _07818_);
  or (_17420_, _17331_, _04953_);
  nor (_17421_, _17420_, _17419_);
  or (_17422_, _17421_, _02334_);
  nor (_17423_, _17422_, _17418_);
  nor (_17424_, _11314_, _07818_);
  nor (_17425_, _17424_, _17331_);
  nor (_17426_, _17425_, _04958_);
  or (_17427_, _17426_, _17423_);
  and (_17429_, _17427_, _02778_);
  nor (_17430_, _17346_, _02778_);
  or (_17431_, _17430_, _17429_);
  and (_17432_, _17431_, _01698_);
  nor (_17433_, _17364_, _01698_);
  or (_17434_, _17433_, _17432_);
  and (_17435_, _17434_, _02082_);
  and (_17436_, _11367_, _03813_);
  nor (_17437_, _17436_, _17331_);
  nor (_17438_, _17437_, _02082_);
  or (_17440_, _17438_, _17435_);
  or (_17441_, _17440_, _39633_);
  or (_17442_, _39632_, \oc8051_golden_model_1.IE [2]);
  and (_17443_, _17442_, _39026_);
  and (_41652_, _17443_, _17441_);
  not (_17444_, \oc8051_golden_model_1.IE [3]);
  nor (_17445_, _03813_, _17444_);
  and (_17446_, _03813_, _04719_);
  nor (_17447_, _17446_, _17445_);
  and (_17448_, _17447_, _01994_);
  nor (_17449_, _07818_, _03434_);
  nor (_17450_, _17449_, _17445_);
  and (_17451_, _17450_, _06188_);
  and (_17452_, _03813_, \oc8051_golden_model_1.ACC [3]);
  nor (_17453_, _17452_, _17445_);
  nor (_17454_, _17453_, _02063_);
  nor (_17455_, _02062_, _17444_);
  or (_17456_, _17455_, _17454_);
  and (_17457_, _17456_, _03006_);
  nor (_17458_, _11394_, _07818_);
  nor (_17461_, _17458_, _17445_);
  nor (_17462_, _17461_, _03006_);
  or (_17463_, _17462_, _17457_);
  and (_17464_, _17463_, _02058_);
  nor (_17465_, _04473_, _17444_);
  and (_17466_, _11398_, _04473_);
  nor (_17467_, _17466_, _17465_);
  nor (_17468_, _17467_, _02058_);
  or (_17469_, _17468_, _17464_);
  and (_17470_, _17469_, _02519_);
  nor (_17472_, _17450_, _02519_);
  or (_17473_, _17472_, _17470_);
  and (_17474_, _17473_, _02549_);
  nor (_17475_, _17453_, _02549_);
  or (_17476_, _17475_, _17474_);
  and (_17477_, _17476_, _02054_);
  and (_17478_, _11408_, _04473_);
  nor (_17479_, _17478_, _17465_);
  nor (_17480_, _17479_, _02054_);
  or (_17481_, _17480_, _02046_);
  or (_17483_, _17481_, _17477_);
  nor (_17484_, _17465_, _11415_);
  nor (_17485_, _17484_, _17467_);
  or (_17486_, _17485_, _02047_);
  and (_17487_, _17486_, _02043_);
  and (_17488_, _17487_, _17483_);
  nor (_17489_, _11433_, _07855_);
  nor (_17490_, _17489_, _17465_);
  nor (_17491_, _17490_, _02043_);
  nor (_17492_, _17491_, _06188_);
  not (_17494_, _17492_);
  nor (_17495_, _17494_, _17488_);
  nor (_17496_, _17495_, _17451_);
  nor (_17497_, _17496_, _02031_);
  and (_17498_, _05166_, _03813_);
  nor (_17499_, _17445_, _02032_);
  not (_17500_, _17499_);
  nor (_17501_, _17500_, _17498_);
  or (_17502_, _17501_, _01765_);
  nor (_17503_, _17502_, _17497_);
  nor (_17504_, _11490_, _07818_);
  nor (_17505_, _17445_, _17504_);
  nor (_17506_, _17505_, _02037_);
  or (_17507_, _17506_, _01994_);
  nor (_17508_, _17507_, _17503_);
  nor (_17509_, _17508_, _17448_);
  or (_17510_, _17509_, _02210_);
  and (_17511_, _11505_, _03813_);
  or (_17512_, _17511_, _17445_);
  or (_17513_, _17512_, _03059_);
  and (_17515_, _17513_, _03061_);
  and (_17516_, _17515_, _17510_);
  and (_17517_, _11511_, _03813_);
  nor (_17518_, _17517_, _17445_);
  nor (_17519_, _17518_, _03061_);
  nor (_17520_, _17519_, _17516_);
  nor (_17521_, _17520_, _02206_);
  nor (_17522_, _17445_, _04153_);
  not (_17523_, _17522_);
  nor (_17524_, _17447_, _02208_);
  and (_17526_, _17524_, _17523_);
  nor (_17527_, _17526_, _17521_);
  nor (_17528_, _17527_, _02342_);
  or (_17529_, _17522_, _03065_);
  nor (_17530_, _17529_, _17453_);
  or (_17531_, _17530_, _02202_);
  nor (_17532_, _17531_, _17528_);
  nor (_17533_, _11503_, _07818_);
  or (_17534_, _17445_, _04953_);
  nor (_17535_, _17534_, _17533_);
  or (_17537_, _17535_, _02334_);
  nor (_17538_, _17537_, _17532_);
  nor (_17539_, _11510_, _07818_);
  nor (_17540_, _17539_, _17445_);
  nor (_17541_, _17540_, _04958_);
  or (_17542_, _17541_, _17538_);
  and (_17543_, _17542_, _02778_);
  nor (_17544_, _17461_, _02778_);
  or (_17545_, _17544_, _17543_);
  and (_17546_, _17545_, _01698_);
  nor (_17548_, _17479_, _01698_);
  or (_17549_, _17548_, _17546_);
  and (_17550_, _17549_, _02082_);
  and (_17551_, _11567_, _03813_);
  nor (_17552_, _17551_, _17445_);
  nor (_17553_, _17552_, _02082_);
  or (_17554_, _17553_, _17550_);
  or (_17555_, _17554_, _39633_);
  or (_17556_, _39632_, \oc8051_golden_model_1.IE [3]);
  and (_17557_, _17556_, _39026_);
  and (_41653_, _17557_, _17555_);
  not (_17559_, \oc8051_golden_model_1.IE [4]);
  nor (_17560_, _03813_, _17559_);
  and (_17561_, _04831_, _03813_);
  nor (_17562_, _17561_, _17560_);
  and (_17563_, _17562_, _01994_);
  nor (_17564_, _04372_, _07818_);
  nor (_17565_, _17564_, _17560_);
  and (_17566_, _17565_, _06188_);
  and (_17567_, _03813_, \oc8051_golden_model_1.ACC [4]);
  nor (_17569_, _17567_, _17560_);
  nor (_17570_, _17569_, _02063_);
  nor (_17571_, _02062_, _17559_);
  or (_17572_, _17571_, _17570_);
  and (_17573_, _17572_, _03006_);
  nor (_17574_, _11611_, _07818_);
  nor (_17575_, _17574_, _17560_);
  nor (_17576_, _17575_, _03006_);
  or (_17577_, _17576_, _17573_);
  and (_17578_, _17577_, _02058_);
  nor (_17580_, _04473_, _17559_);
  and (_17581_, _11597_, _04473_);
  nor (_17582_, _17581_, _17580_);
  nor (_17583_, _17582_, _02058_);
  or (_17584_, _17583_, _17578_);
  and (_17585_, _17584_, _02519_);
  nor (_17586_, _17565_, _02519_);
  or (_17587_, _17586_, _17585_);
  and (_17588_, _17587_, _02549_);
  nor (_17589_, _17569_, _02549_);
  or (_17591_, _17589_, _17588_);
  and (_17592_, _17591_, _02054_);
  and (_17593_, _11595_, _04473_);
  nor (_17594_, _17593_, _17580_);
  nor (_17595_, _17594_, _02054_);
  or (_17596_, _17595_, _17592_);
  and (_17597_, _17596_, _02047_);
  nor (_17598_, _17580_, _11628_);
  nor (_17599_, _17598_, _17582_);
  and (_17600_, _17599_, _02046_);
  or (_17602_, _17600_, _17597_);
  and (_17603_, _17602_, _02043_);
  nor (_17604_, _11646_, _07855_);
  nor (_17605_, _17604_, _17580_);
  nor (_17606_, _17605_, _02043_);
  nor (_17607_, _17606_, _06188_);
  not (_17608_, _17607_);
  nor (_17609_, _17608_, _17603_);
  nor (_17610_, _17609_, _17566_);
  nor (_17611_, _17610_, _02031_);
  and (_17613_, _05303_, _03813_);
  nor (_17614_, _17560_, _02032_);
  not (_17615_, _17614_);
  nor (_17616_, _17615_, _17613_);
  or (_17617_, _17616_, _01765_);
  nor (_17618_, _17617_, _17611_);
  nor (_17619_, _11704_, _07818_);
  nor (_17620_, _17560_, _17619_);
  nor (_17621_, _17620_, _02037_);
  or (_17622_, _17621_, _01994_);
  nor (_17624_, _17622_, _17618_);
  nor (_17625_, _17624_, _17563_);
  or (_17626_, _17625_, _02210_);
  and (_17627_, _11592_, _03813_);
  or (_17628_, _17627_, _17560_);
  or (_17629_, _17628_, _03059_);
  and (_17630_, _17629_, _03061_);
  and (_17631_, _17630_, _17626_);
  and (_17632_, _11588_, _03813_);
  nor (_17633_, _17632_, _17560_);
  nor (_17635_, _17633_, _03061_);
  nor (_17636_, _17635_, _17631_);
  nor (_17637_, _17636_, _02206_);
  nor (_17638_, _17560_, _04420_);
  not (_17639_, _17638_);
  nor (_17640_, _17562_, _02208_);
  and (_17641_, _17640_, _17639_);
  nor (_17642_, _17641_, _17637_);
  nor (_17643_, _17642_, _02342_);
  or (_17644_, _17638_, _03065_);
  nor (_17646_, _17644_, _17569_);
  or (_17647_, _17646_, _02202_);
  nor (_17648_, _17647_, _17643_);
  nor (_17649_, _11590_, _07818_);
  or (_17650_, _17560_, _04953_);
  nor (_17651_, _17650_, _17649_);
  or (_17652_, _17651_, _02334_);
  nor (_17653_, _17652_, _17648_);
  nor (_17654_, _11587_, _07818_);
  nor (_17655_, _17654_, _17560_);
  nor (_17657_, _17655_, _04958_);
  or (_17658_, _17657_, _17653_);
  and (_17659_, _17658_, _02778_);
  nor (_17660_, _17575_, _02778_);
  or (_17661_, _17660_, _17659_);
  and (_17662_, _17661_, _01698_);
  nor (_17663_, _17594_, _01698_);
  or (_17664_, _17663_, _17662_);
  and (_17665_, _17664_, _02082_);
  and (_17666_, _11771_, _03813_);
  nor (_17668_, _17666_, _17560_);
  nor (_17669_, _17668_, _02082_);
  or (_17670_, _17669_, _17665_);
  or (_17671_, _17670_, _39633_);
  or (_17672_, _39632_, \oc8051_golden_model_1.IE [4]);
  and (_17673_, _17672_, _39026_);
  and (_41655_, _17673_, _17671_);
  not (_17674_, \oc8051_golden_model_1.IE [5]);
  nor (_17675_, _03813_, _17674_);
  and (_17676_, _04827_, _03813_);
  nor (_17678_, _17676_, _17675_);
  and (_17679_, _17678_, _01994_);
  nor (_17680_, _04057_, _07818_);
  nor (_17681_, _17680_, _17675_);
  and (_17682_, _17681_, _06188_);
  and (_17683_, _03813_, \oc8051_golden_model_1.ACC [5]);
  nor (_17684_, _17683_, _17675_);
  nor (_17685_, _17684_, _02063_);
  nor (_17686_, _02062_, _17674_);
  or (_17687_, _17686_, _17685_);
  and (_17689_, _17687_, _03006_);
  nor (_17690_, _11804_, _07818_);
  nor (_17691_, _17690_, _17675_);
  nor (_17692_, _17691_, _03006_);
  or (_17693_, _17692_, _17689_);
  and (_17694_, _17693_, _02058_);
  nor (_17695_, _04473_, _17674_);
  and (_17696_, _11789_, _04473_);
  nor (_17697_, _17696_, _17695_);
  nor (_17698_, _17697_, _02058_);
  or (_17699_, _17698_, _17694_);
  and (_17700_, _17699_, _02519_);
  nor (_17701_, _17681_, _02519_);
  or (_17702_, _17701_, _17700_);
  and (_17703_, _17702_, _02549_);
  nor (_17704_, _17684_, _02549_);
  or (_17705_, _17704_, _17703_);
  and (_17706_, _17705_, _02054_);
  and (_17707_, _11816_, _04473_);
  nor (_17708_, _17707_, _17695_);
  nor (_17710_, _17708_, _02054_);
  or (_17711_, _17710_, _17706_);
  and (_17712_, _17711_, _02047_);
  nor (_17713_, _17695_, _11823_);
  nor (_17714_, _17713_, _17697_);
  and (_17715_, _17714_, _02046_);
  or (_17716_, _17715_, _17712_);
  and (_17717_, _17716_, _02043_);
  nor (_17718_, _11841_, _07855_);
  nor (_17719_, _17718_, _17695_);
  nor (_17721_, _17719_, _02043_);
  nor (_17722_, _17721_, _06188_);
  not (_17723_, _17722_);
  nor (_17724_, _17723_, _17717_);
  nor (_17725_, _17724_, _17682_);
  nor (_17726_, _17725_, _02031_);
  and (_17727_, _05258_, _03813_);
  nor (_17728_, _17675_, _02032_);
  not (_17729_, _17728_);
  nor (_17730_, _17729_, _17727_);
  or (_17732_, _17730_, _01765_);
  nor (_17733_, _17732_, _17726_);
  nor (_17734_, _11900_, _07818_);
  nor (_17735_, _17734_, _17675_);
  nor (_17736_, _17735_, _02037_);
  or (_17737_, _17736_, _01994_);
  nor (_17738_, _17737_, _17733_);
  nor (_17739_, _17738_, _17679_);
  or (_17740_, _17739_, _02210_);
  and (_17741_, _11915_, _03813_);
  or (_17743_, _17741_, _17675_);
  or (_17744_, _17743_, _03059_);
  and (_17745_, _17744_, _03061_);
  and (_17746_, _17745_, _17740_);
  and (_17747_, _11786_, _03813_);
  nor (_17748_, _17747_, _17675_);
  nor (_17749_, _17748_, _03061_);
  nor (_17750_, _17749_, _17746_);
  nor (_17751_, _17750_, _02206_);
  nor (_17752_, _17675_, _04104_);
  not (_17754_, _17752_);
  nor (_17755_, _17678_, _02208_);
  and (_17756_, _17755_, _17754_);
  nor (_17757_, _17756_, _17751_);
  nor (_17758_, _17757_, _02342_);
  or (_17759_, _17752_, _03065_);
  nor (_17760_, _17759_, _17684_);
  or (_17761_, _17760_, _02202_);
  nor (_17762_, _17761_, _17758_);
  nor (_17763_, _11913_, _07818_);
  or (_17765_, _17675_, _04953_);
  nor (_17766_, _17765_, _17763_);
  or (_17767_, _17766_, _02334_);
  nor (_17768_, _17767_, _17762_);
  nor (_17769_, _11785_, _07818_);
  nor (_17770_, _17769_, _17675_);
  nor (_17771_, _17770_, _04958_);
  or (_17772_, _17771_, _17768_);
  and (_17773_, _17772_, _02778_);
  nor (_17774_, _17691_, _02778_);
  or (_17776_, _17774_, _17773_);
  and (_17777_, _17776_, _01698_);
  nor (_17778_, _17708_, _01698_);
  nor (_17779_, _17778_, _02081_);
  not (_17780_, _17779_);
  nor (_17781_, _17780_, _17777_);
  and (_17782_, _11974_, _03813_);
  nor (_17783_, _17782_, _17675_);
  and (_17784_, _17783_, _02081_);
  nor (_17785_, _17784_, _17781_);
  or (_17787_, _17785_, _39633_);
  or (_17788_, _39632_, \oc8051_golden_model_1.IE [5]);
  and (_17789_, _17788_, _39026_);
  and (_41656_, _17789_, _17787_);
  not (_17790_, \oc8051_golden_model_1.IE [6]);
  nor (_17791_, _03813_, _17790_);
  and (_17792_, _12103_, _03813_);
  nor (_17793_, _17792_, _17791_);
  and (_17794_, _17793_, _01994_);
  nor (_17795_, _03964_, _07818_);
  nor (_17797_, _17795_, _17791_);
  and (_17798_, _17797_, _06188_);
  and (_17799_, _03813_, \oc8051_golden_model_1.ACC [6]);
  nor (_17800_, _17799_, _17791_);
  nor (_17801_, _17800_, _02063_);
  nor (_17802_, _02062_, _17790_);
  or (_17803_, _17802_, _17801_);
  and (_17804_, _17803_, _03006_);
  nor (_17805_, _11993_, _07818_);
  nor (_17806_, _17805_, _17791_);
  nor (_17808_, _17806_, _03006_);
  or (_17809_, _17808_, _17804_);
  and (_17810_, _17809_, _02058_);
  nor (_17811_, _04473_, _17790_);
  and (_17812_, _11990_, _04473_);
  nor (_17813_, _17812_, _17811_);
  nor (_17814_, _17813_, _02058_);
  or (_17815_, _17814_, _17810_);
  and (_17816_, _17815_, _02519_);
  nor (_17817_, _17797_, _02519_);
  or (_17819_, _17817_, _17816_);
  and (_17820_, _17819_, _02549_);
  nor (_17821_, _17800_, _02549_);
  or (_17822_, _17821_, _17820_);
  and (_17823_, _17822_, _02054_);
  and (_17824_, _12017_, _04473_);
  nor (_17825_, _17824_, _17811_);
  nor (_17826_, _17825_, _02054_);
  or (_17827_, _17826_, _17823_);
  and (_17828_, _17827_, _02047_);
  nor (_17830_, _17811_, _12024_);
  nor (_17831_, _17830_, _17813_);
  and (_17832_, _17831_, _02046_);
  or (_17833_, _17832_, _17828_);
  and (_17834_, _17833_, _02043_);
  nor (_17835_, _12042_, _07855_);
  nor (_17836_, _17835_, _17811_);
  nor (_17837_, _17836_, _02043_);
  nor (_17838_, _17837_, _06188_);
  not (_17839_, _17838_);
  nor (_17841_, _17839_, _17834_);
  nor (_17842_, _17841_, _17798_);
  nor (_17843_, _17842_, _02031_);
  and (_17844_, _05029_, _03813_);
  nor (_17845_, _17791_, _02032_);
  not (_17846_, _17845_);
  nor (_17847_, _17846_, _17844_);
  or (_17848_, _17847_, _01765_);
  nor (_17849_, _17848_, _17843_);
  nor (_17850_, _12096_, _07818_);
  nor (_17852_, _17850_, _17791_);
  nor (_17853_, _17852_, _02037_);
  or (_17854_, _17853_, _01994_);
  nor (_17855_, _17854_, _17849_);
  nor (_17856_, _17855_, _17794_);
  or (_17857_, _17856_, _02210_);
  and (_17858_, _12112_, _03813_);
  or (_17859_, _17858_, _17791_);
  or (_17860_, _17859_, _03059_);
  and (_17861_, _17860_, _03061_);
  and (_17863_, _17861_, _17857_);
  and (_17864_, _12118_, _03813_);
  nor (_17865_, _17864_, _17791_);
  nor (_17866_, _17865_, _03061_);
  nor (_17867_, _17866_, _17863_);
  nor (_17868_, _17867_, _02206_);
  nor (_17869_, _17791_, _04011_);
  not (_17870_, _17869_);
  nor (_17871_, _17793_, _02208_);
  and (_17872_, _17871_, _17870_);
  nor (_17873_, _17872_, _17868_);
  nor (_17874_, _17873_, _02342_);
  or (_17875_, _17869_, _03065_);
  nor (_17876_, _17875_, _17800_);
  or (_17877_, _17876_, _02202_);
  nor (_17878_, _17877_, _17874_);
  nor (_17879_, _12110_, _07818_);
  or (_17880_, _17791_, _04953_);
  nor (_17881_, _17880_, _17879_);
  or (_17882_, _17881_, _02334_);
  nor (_17884_, _17882_, _17878_);
  nor (_17885_, _12117_, _07818_);
  nor (_17886_, _17885_, _17791_);
  nor (_17887_, _17886_, _04958_);
  or (_17888_, _17887_, _17884_);
  and (_17889_, _17888_, _02778_);
  nor (_17890_, _17806_, _02778_);
  or (_17891_, _17890_, _17889_);
  and (_17892_, _17891_, _01698_);
  nor (_17893_, _17825_, _01698_);
  or (_17895_, _17893_, _17892_);
  and (_17896_, _17895_, _02082_);
  and (_17897_, _12178_, _03813_);
  nor (_17898_, _17897_, _17791_);
  nor (_17899_, _17898_, _02082_);
  or (_17900_, _17899_, _17896_);
  or (_17901_, _17900_, _39633_);
  or (_17902_, _39632_, \oc8051_golden_model_1.IE [6]);
  and (_17903_, _17902_, _39026_);
  and (_41657_, _17903_, _17901_);
  nor (_17905_, _04257_, _07925_);
  not (_17906_, \oc8051_golden_model_1.IP [0]);
  nor (_17907_, _03844_, _17906_);
  and (_17908_, _03844_, _04837_);
  nor (_17909_, _17908_, _17907_);
  nor (_17910_, _17909_, _02208_);
  not (_17911_, _17910_);
  nor (_17912_, _17911_, _17905_);
  and (_17913_, _10792_, _03844_);
  nor (_17914_, _17913_, _17907_);
  nor (_17916_, _17914_, _03061_);
  and (_17917_, _17909_, _01994_);
  and (_17918_, _03844_, _03002_);
  nor (_17919_, _17918_, _17907_);
  and (_17920_, _17919_, _06188_);
  and (_17921_, _03844_, \oc8051_golden_model_1.ACC [0]);
  nor (_17922_, _17921_, _17907_);
  nor (_17923_, _17922_, _02063_);
  nor (_17924_, _02062_, _17906_);
  or (_17925_, _17924_, _17923_);
  and (_17927_, _17925_, _03006_);
  nor (_17928_, _17905_, _17907_);
  nor (_17929_, _17928_, _03006_);
  or (_17930_, _17929_, _17927_);
  and (_17931_, _17930_, _02058_);
  nor (_17932_, _04481_, _17906_);
  and (_17933_, _10814_, _04481_);
  nor (_17934_, _17933_, _17932_);
  nor (_17935_, _17934_, _02058_);
  nor (_17936_, _17935_, _17931_);
  nor (_17938_, _17936_, _02155_);
  nor (_17939_, _17919_, _02519_);
  or (_17940_, _17939_, _17938_);
  and (_17941_, _17940_, _02549_);
  nor (_17942_, _17922_, _02549_);
  or (_17943_, _17942_, _17941_);
  and (_17944_, _17943_, _02054_);
  and (_17945_, _17907_, _02053_);
  or (_17946_, _17945_, _17944_);
  and (_17947_, _17946_, _02047_);
  nor (_17949_, _17928_, _02047_);
  or (_17950_, _17949_, _17947_);
  and (_17951_, _17950_, _02043_);
  nor (_17952_, _10798_, _07962_);
  nor (_17953_, _17952_, _17932_);
  nor (_17954_, _17953_, _02043_);
  or (_17955_, _17954_, _06188_);
  nor (_17956_, _17955_, _17951_);
  nor (_17957_, _17956_, _17920_);
  nor (_17958_, _17957_, _02031_);
  and (_17960_, _05120_, _03844_);
  nor (_17961_, _17907_, _02032_);
  not (_17962_, _17961_);
  nor (_17963_, _17962_, _17960_);
  or (_17964_, _17963_, _01765_);
  nor (_17965_, _17964_, _17958_);
  nor (_17966_, _10898_, _07925_);
  nor (_17967_, _17966_, _17907_);
  nor (_17968_, _17967_, _02037_);
  or (_17969_, _17968_, _01994_);
  nor (_17971_, _17969_, _17965_);
  nor (_17972_, _17971_, _17917_);
  or (_17973_, _17972_, _02210_);
  and (_17974_, _10914_, _03844_);
  or (_17975_, _17974_, _17907_);
  or (_17976_, _17975_, _03059_);
  and (_17977_, _17976_, _03061_);
  and (_17978_, _17977_, _17973_);
  nor (_17979_, _17978_, _17916_);
  nor (_17980_, _17979_, _02206_);
  nor (_17982_, _17980_, _17912_);
  nor (_17983_, _17982_, _02342_);
  nor (_17984_, _17907_, _04257_);
  or (_17985_, _17984_, _03065_);
  nor (_17986_, _17985_, _17922_);
  or (_17987_, _17986_, _02202_);
  nor (_17988_, _17987_, _17983_);
  nor (_17989_, _10913_, _07925_);
  or (_17990_, _17907_, _04953_);
  nor (_17991_, _17990_, _17989_);
  or (_17993_, _17991_, _02334_);
  nor (_17994_, _17993_, _17988_);
  nor (_17995_, _10789_, _07925_);
  nor (_17996_, _17995_, _17907_);
  nor (_17997_, _17996_, _04958_);
  or (_17998_, _17997_, _17994_);
  and (_17999_, _17998_, _02778_);
  nor (_18000_, _17928_, _02778_);
  or (_18001_, _18000_, _17999_);
  and (_18002_, _18001_, _01698_);
  and (_18004_, _17907_, _01697_);
  or (_18005_, _18004_, _18002_);
  and (_18006_, _18005_, _02082_);
  nor (_18007_, _17928_, _02082_);
  or (_18008_, _18007_, _18006_);
  or (_18009_, _18008_, _39633_);
  or (_18010_, _39632_, \oc8051_golden_model_1.IP [0]);
  and (_18011_, _18010_, _39026_);
  and (_41659_, _18011_, _18009_);
  not (_18012_, \oc8051_golden_model_1.IP [1]);
  nor (_18014_, _03844_, _18012_);
  and (_18015_, _05075_, _03844_);
  or (_18016_, _18015_, _18014_);
  and (_18017_, _18016_, _02031_);
  nor (_18018_, _03844_, \oc8051_golden_model_1.IP [1]);
  and (_18019_, _03844_, _01804_);
  nor (_18020_, _18019_, _18018_);
  and (_18021_, _18020_, _02062_);
  nor (_18022_, _02062_, _18012_);
  or (_18023_, _18022_, _18021_);
  and (_18025_, _18023_, _03006_);
  and (_18026_, _11001_, _03844_);
  nor (_18027_, _18026_, _18018_);
  and (_18028_, _18027_, _02158_);
  or (_18029_, _18028_, _18025_);
  and (_18030_, _18029_, _02058_);
  nor (_18031_, _04481_, _18012_);
  and (_18032_, _11005_, _04481_);
  nor (_18033_, _18032_, _18031_);
  nor (_18034_, _18033_, _02058_);
  or (_18036_, _18034_, _18030_);
  and (_18037_, _18036_, _02519_);
  nor (_18038_, _07925_, _03161_);
  nor (_18039_, _18038_, _18014_);
  nor (_18040_, _18039_, _02519_);
  or (_18041_, _18040_, _18037_);
  nor (_18042_, _18041_, _02153_);
  nor (_18043_, _18020_, _02549_);
  or (_18044_, _18043_, _02053_);
  nor (_18045_, _18044_, _18042_);
  and (_18047_, _10992_, _04481_);
  nor (_18048_, _18047_, _18031_);
  nor (_18049_, _18048_, _02054_);
  or (_18050_, _18049_, _18045_);
  and (_18051_, _18050_, _02047_);
  nor (_18052_, _18031_, _11020_);
  nor (_18053_, _18052_, _18033_);
  and (_18054_, _18053_, _02046_);
  or (_18055_, _18054_, _18051_);
  and (_18056_, _18055_, _02043_);
  nor (_18057_, _11038_, _07962_);
  nor (_18058_, _18057_, _18031_);
  nor (_18059_, _18058_, _02043_);
  nor (_18060_, _18059_, _06188_);
  not (_18061_, _18060_);
  nor (_18062_, _18061_, _18056_);
  and (_18063_, _18039_, _06188_);
  or (_18064_, _18063_, _02031_);
  nor (_18065_, _18064_, _18062_);
  or (_18066_, _18065_, _18017_);
  and (_18068_, _18066_, _02037_);
  nor (_18069_, _11096_, _07925_);
  nor (_18070_, _18069_, _18014_);
  nor (_18071_, _18070_, _02037_);
  nor (_18072_, _18071_, _18068_);
  nor (_18073_, _18072_, _07629_);
  not (_18074_, _18018_);
  nor (_18075_, _10989_, _07925_);
  nor (_18076_, _18075_, _03059_);
  and (_18077_, _03844_, _02893_);
  nor (_18079_, _18077_, _01995_);
  or (_18080_, _18079_, _18076_);
  and (_18081_, _18080_, _18074_);
  nor (_18082_, _18081_, _18073_);
  nor (_18083_, _18082_, _02331_);
  nor (_18084_, _11113_, _07925_);
  nor (_18085_, _18084_, _03061_);
  and (_18086_, _18085_, _18074_);
  nor (_18087_, _18086_, _18083_);
  nor (_18088_, _18087_, _02206_);
  nor (_18090_, _10988_, _07925_);
  nor (_18091_, _18090_, _02208_);
  and (_18092_, _18091_, _18074_);
  nor (_18093_, _18092_, _18088_);
  nor (_18094_, _18093_, _02342_);
  nor (_18095_, _18014_, _04209_);
  nor (_18096_, _18095_, _03065_);
  and (_18097_, _18096_, _18020_);
  nor (_18098_, _18097_, _18094_);
  or (_18099_, _18098_, _17216_);
  and (_18101_, _18019_, _04208_);
  nor (_18102_, _18101_, _04958_);
  and (_18103_, _18102_, _18074_);
  nor (_18104_, _18103_, _02366_);
  and (_18105_, _18077_, _04208_);
  or (_18106_, _18018_, _04953_);
  or (_18107_, _18106_, _18105_);
  and (_18108_, _18107_, _18104_);
  and (_18109_, _18108_, _18099_);
  nor (_18110_, _18027_, _02778_);
  or (_18112_, _18110_, _01697_);
  nor (_18113_, _18112_, _18109_);
  nor (_18114_, _18048_, _01698_);
  or (_18115_, _18114_, _02081_);
  nor (_18116_, _18115_, _18113_);
  nor (_18117_, _18026_, _18014_);
  and (_18118_, _18117_, _02081_);
  nor (_18119_, _18118_, _18116_);
  or (_18120_, _18119_, _39633_);
  or (_18121_, _39632_, \oc8051_golden_model_1.IP [1]);
  and (_18123_, _18121_, _39026_);
  and (_41660_, _18123_, _18120_);
  not (_18124_, \oc8051_golden_model_1.IP [2]);
  nor (_18125_, _03844_, _18124_);
  and (_18126_, _11315_, _03844_);
  nor (_18127_, _18126_, _18125_);
  nor (_18128_, _18127_, _03061_);
  and (_18129_, _03844_, _04866_);
  nor (_18130_, _18129_, _18125_);
  and (_18131_, _18130_, _01994_);
  nor (_18133_, _07925_, _03624_);
  nor (_18134_, _18133_, _18125_);
  and (_18135_, _18134_, _06188_);
  and (_18136_, _03844_, \oc8051_golden_model_1.ACC [2]);
  nor (_18137_, _18136_, _18125_);
  nor (_18138_, _18137_, _02063_);
  nor (_18139_, _02062_, _18124_);
  or (_18140_, _18139_, _18138_);
  and (_18141_, _18140_, _03006_);
  nor (_18142_, _11199_, _07925_);
  nor (_18144_, _18142_, _18125_);
  nor (_18145_, _18144_, _03006_);
  or (_18146_, _18145_, _18141_);
  and (_18147_, _18146_, _02058_);
  nor (_18148_, _04481_, _18124_);
  and (_18149_, _11194_, _04481_);
  nor (_18150_, _18149_, _18148_);
  nor (_18151_, _18150_, _02058_);
  or (_18152_, _18151_, _02155_);
  or (_18153_, _18152_, _18147_);
  nand (_18155_, _18134_, _02155_);
  and (_18156_, _18155_, _18153_);
  and (_18157_, _18156_, _02549_);
  nor (_18158_, _18137_, _02549_);
  or (_18159_, _18158_, _18157_);
  and (_18160_, _18159_, _02054_);
  and (_18161_, _11192_, _04481_);
  nor (_18162_, _18161_, _18148_);
  nor (_18163_, _18162_, _02054_);
  or (_18164_, _18163_, _02046_);
  or (_18166_, _18164_, _18160_);
  nor (_18167_, _18148_, _11223_);
  nor (_18168_, _18167_, _18150_);
  or (_18169_, _18168_, _02047_);
  and (_18170_, _18169_, _02043_);
  and (_18171_, _18170_, _18166_);
  nor (_18172_, _11241_, _07962_);
  nor (_18173_, _18172_, _18148_);
  nor (_18174_, _18173_, _02043_);
  nor (_18175_, _18174_, _06188_);
  not (_18177_, _18175_);
  nor (_18178_, _18177_, _18171_);
  nor (_18179_, _18178_, _18135_);
  nor (_18180_, _18179_, _02031_);
  and (_18181_, _05211_, _03844_);
  nor (_18182_, _18125_, _02032_);
  not (_18183_, _18182_);
  nor (_18184_, _18183_, _18181_);
  or (_18185_, _18184_, _01765_);
  nor (_18186_, _18185_, _18180_);
  nor (_18188_, _11298_, _07925_);
  nor (_18189_, _18188_, _18125_);
  nor (_18190_, _18189_, _02037_);
  or (_18191_, _18190_, _01994_);
  nor (_18192_, _18191_, _18186_);
  nor (_18193_, _18192_, _18131_);
  or (_18194_, _18193_, _02210_);
  and (_18195_, _11189_, _03844_);
  or (_18196_, _18195_, _18125_);
  or (_18197_, _18196_, _03059_);
  and (_18199_, _18197_, _03061_);
  and (_18200_, _18199_, _18194_);
  nor (_18201_, _18200_, _18128_);
  nor (_18202_, _18201_, _02206_);
  nor (_18203_, _18125_, _04309_);
  not (_18204_, _18203_);
  nor (_18205_, _18130_, _02208_);
  and (_18206_, _18205_, _18204_);
  nor (_18207_, _18206_, _18202_);
  nor (_18208_, _18207_, _02342_);
  or (_18210_, _18203_, _03065_);
  nor (_18211_, _18210_, _18137_);
  or (_18212_, _18211_, _02202_);
  nor (_18213_, _18212_, _18208_);
  nor (_18214_, _11187_, _07925_);
  or (_18215_, _18125_, _04953_);
  nor (_18216_, _18215_, _18214_);
  or (_18217_, _18216_, _02334_);
  nor (_18218_, _18217_, _18213_);
  nor (_18219_, _11314_, _07925_);
  nor (_18221_, _18219_, _18125_);
  nor (_18222_, _18221_, _04958_);
  or (_18223_, _18222_, _18218_);
  and (_18224_, _18223_, _02778_);
  nor (_18225_, _18144_, _02778_);
  or (_18226_, _18225_, _18224_);
  and (_18227_, _18226_, _01698_);
  nor (_18228_, _18162_, _01698_);
  or (_18229_, _18228_, _18227_);
  and (_18230_, _18229_, _02082_);
  and (_18231_, _11367_, _03844_);
  nor (_18232_, _18231_, _18125_);
  nor (_18233_, _18232_, _02082_);
  or (_18234_, _18233_, _18230_);
  or (_18235_, _18234_, _39633_);
  or (_18236_, _39632_, \oc8051_golden_model_1.IP [2]);
  and (_18237_, _18236_, _39026_);
  and (_41661_, _18237_, _18235_);
  not (_18238_, \oc8051_golden_model_1.IP [3]);
  nor (_18239_, _03844_, _18238_);
  and (_18241_, _03844_, _04719_);
  nor (_18242_, _18241_, _18239_);
  and (_18243_, _18242_, _01994_);
  nor (_18244_, _07925_, _03434_);
  nor (_18245_, _18244_, _18239_);
  and (_18246_, _18245_, _06188_);
  and (_18247_, _03844_, \oc8051_golden_model_1.ACC [3]);
  nor (_18248_, _18247_, _18239_);
  nor (_18249_, _18248_, _02063_);
  nor (_18250_, _02062_, _18238_);
  or (_18252_, _18250_, _18249_);
  and (_18253_, _18252_, _03006_);
  nor (_18254_, _11394_, _07925_);
  nor (_18255_, _18254_, _18239_);
  nor (_18256_, _18255_, _03006_);
  or (_18257_, _18256_, _18253_);
  and (_18258_, _18257_, _02058_);
  nor (_18259_, _04481_, _18238_);
  and (_18260_, _11398_, _04481_);
  nor (_18261_, _18260_, _18259_);
  nor (_18263_, _18261_, _02058_);
  or (_18264_, _18263_, _18258_);
  and (_18265_, _18264_, _02519_);
  nor (_18266_, _18245_, _02519_);
  or (_18267_, _18266_, _18265_);
  and (_18268_, _18267_, _02549_);
  nor (_18269_, _18248_, _02549_);
  or (_18270_, _18269_, _18268_);
  and (_18271_, _18270_, _02054_);
  and (_18272_, _11408_, _04481_);
  nor (_18274_, _18272_, _18259_);
  nor (_18275_, _18274_, _02054_);
  or (_18276_, _18275_, _18271_);
  and (_18277_, _18276_, _02047_);
  nor (_18278_, _18259_, _11415_);
  nor (_18279_, _18278_, _18261_);
  and (_18280_, _18279_, _02046_);
  or (_18281_, _18280_, _18277_);
  and (_18282_, _18281_, _02043_);
  nor (_18283_, _11433_, _07962_);
  nor (_18285_, _18283_, _18259_);
  nor (_18286_, _18285_, _02043_);
  nor (_18287_, _18286_, _06188_);
  not (_18288_, _18287_);
  nor (_18289_, _18288_, _18282_);
  nor (_18290_, _18289_, _18246_);
  nor (_18291_, _18290_, _02031_);
  and (_18292_, _05166_, _03844_);
  nor (_18293_, _18239_, _02032_);
  not (_18294_, _18293_);
  nor (_18296_, _18294_, _18292_);
  or (_18297_, _18296_, _01765_);
  nor (_18298_, _18297_, _18291_);
  nor (_18299_, _11490_, _07925_);
  nor (_18300_, _18239_, _18299_);
  nor (_18301_, _18300_, _02037_);
  or (_18302_, _18301_, _01994_);
  nor (_18303_, _18302_, _18298_);
  nor (_18304_, _18303_, _18243_);
  or (_18305_, _18304_, _02210_);
  and (_18307_, _11505_, _03844_);
  or (_18308_, _18307_, _18239_);
  or (_18309_, _18308_, _03059_);
  and (_18310_, _18309_, _03061_);
  and (_18311_, _18310_, _18305_);
  and (_18312_, _11511_, _03844_);
  nor (_18313_, _18312_, _18239_);
  nor (_18314_, _18313_, _03061_);
  nor (_18315_, _18314_, _18311_);
  nor (_18316_, _18315_, _02206_);
  nor (_18318_, _18239_, _04153_);
  not (_18319_, _18318_);
  nor (_18320_, _18242_, _02208_);
  and (_18321_, _18320_, _18319_);
  nor (_18322_, _18321_, _18316_);
  nor (_18323_, _18322_, _02342_);
  or (_18324_, _18318_, _03065_);
  nor (_18325_, _18324_, _18248_);
  or (_18326_, _18325_, _02202_);
  nor (_18327_, _18326_, _18323_);
  nor (_18328_, _11503_, _07925_);
  or (_18329_, _18239_, _04953_);
  nor (_18330_, _18329_, _18328_);
  or (_18331_, _18330_, _02334_);
  nor (_18332_, _18331_, _18327_);
  nor (_18333_, _11510_, _07925_);
  nor (_18334_, _18333_, _18239_);
  nor (_18335_, _18334_, _04958_);
  or (_18336_, _18335_, _18332_);
  and (_18337_, _18336_, _02778_);
  nor (_18340_, _18255_, _02778_);
  or (_18341_, _18340_, _18337_);
  and (_18342_, _18341_, _01698_);
  nor (_18343_, _18274_, _01698_);
  or (_18344_, _18343_, _18342_);
  and (_18345_, _18344_, _02082_);
  and (_18346_, _11567_, _03844_);
  nor (_18347_, _18346_, _18239_);
  nor (_18348_, _18347_, _02082_);
  or (_18349_, _18348_, _18345_);
  or (_18351_, _18349_, _39633_);
  or (_18352_, _39632_, \oc8051_golden_model_1.IP [3]);
  and (_18353_, _18352_, _39026_);
  and (_41662_, _18353_, _18351_);
  not (_18354_, \oc8051_golden_model_1.IP [4]);
  nor (_18355_, _03844_, _18354_);
  and (_18356_, _04831_, _03844_);
  nor (_18357_, _18356_, _18355_);
  and (_18358_, _18357_, _01994_);
  nor (_18359_, _04372_, _07925_);
  nor (_18361_, _18359_, _18355_);
  and (_18362_, _18361_, _06188_);
  and (_18363_, _03844_, \oc8051_golden_model_1.ACC [4]);
  nor (_18364_, _18363_, _18355_);
  nor (_18365_, _18364_, _02063_);
  nor (_18366_, _02062_, _18354_);
  or (_18367_, _18366_, _18365_);
  and (_18368_, _18367_, _03006_);
  nor (_18369_, _11611_, _07925_);
  nor (_18370_, _18369_, _18355_);
  nor (_18372_, _18370_, _03006_);
  or (_18373_, _18372_, _18368_);
  and (_18374_, _18373_, _02058_);
  nor (_18375_, _04481_, _18354_);
  and (_18376_, _11597_, _04481_);
  nor (_18377_, _18376_, _18375_);
  nor (_18378_, _18377_, _02058_);
  or (_18379_, _18378_, _18374_);
  and (_18380_, _18379_, _02519_);
  nor (_18381_, _18361_, _02519_);
  or (_18383_, _18381_, _18380_);
  and (_18384_, _18383_, _02549_);
  nor (_18385_, _18364_, _02549_);
  or (_18386_, _18385_, _18384_);
  and (_18387_, _18386_, _02054_);
  and (_18388_, _11595_, _04481_);
  nor (_18389_, _18388_, _18375_);
  nor (_18390_, _18389_, _02054_);
  or (_18391_, _18390_, _18387_);
  and (_18392_, _18391_, _02047_);
  nor (_18394_, _18375_, _11628_);
  nor (_18395_, _18394_, _18377_);
  and (_18396_, _18395_, _02046_);
  or (_18397_, _18396_, _18392_);
  and (_18398_, _18397_, _02043_);
  nor (_18399_, _11646_, _07962_);
  nor (_18400_, _18399_, _18375_);
  nor (_18401_, _18400_, _02043_);
  nor (_18402_, _18401_, _06188_);
  not (_18403_, _18402_);
  nor (_18404_, _18403_, _18398_);
  nor (_18405_, _18404_, _18362_);
  nor (_18406_, _18405_, _02031_);
  and (_18407_, _05303_, _03844_);
  nor (_18408_, _18355_, _02032_);
  not (_18409_, _18408_);
  nor (_18410_, _18409_, _18407_);
  or (_18411_, _18410_, _01765_);
  nor (_18412_, _18411_, _18406_);
  nor (_18413_, _11704_, _07925_);
  nor (_18415_, _18355_, _18413_);
  nor (_18416_, _18415_, _02037_);
  or (_18417_, _18416_, _01994_);
  nor (_18418_, _18417_, _18412_);
  nor (_18419_, _18418_, _18358_);
  or (_18420_, _18419_, _02210_);
  and (_18421_, _11592_, _03844_);
  or (_18422_, _18421_, _18355_);
  or (_18423_, _18422_, _03059_);
  and (_18424_, _18423_, _03061_);
  and (_18426_, _18424_, _18420_);
  and (_18427_, _11588_, _03844_);
  nor (_18428_, _18427_, _18355_);
  nor (_18429_, _18428_, _03061_);
  nor (_18430_, _18429_, _18426_);
  nor (_18431_, _18430_, _02206_);
  nor (_18432_, _18355_, _04420_);
  not (_18433_, _18432_);
  nor (_18434_, _18357_, _02208_);
  and (_18435_, _18434_, _18433_);
  nor (_18437_, _18435_, _18431_);
  nor (_18438_, _18437_, _02342_);
  or (_18439_, _18432_, _03065_);
  nor (_18440_, _18439_, _18364_);
  or (_18441_, _18440_, _02202_);
  nor (_18442_, _18441_, _18438_);
  nor (_18443_, _11590_, _07925_);
  or (_18444_, _18355_, _04953_);
  nor (_18445_, _18444_, _18443_);
  or (_18446_, _18445_, _02334_);
  nor (_18448_, _18446_, _18442_);
  nor (_18449_, _11587_, _07925_);
  nor (_18450_, _18449_, _18355_);
  nor (_18451_, _18450_, _04958_);
  or (_18452_, _18451_, _18448_);
  and (_18453_, _18452_, _02778_);
  nor (_18454_, _18370_, _02778_);
  or (_18455_, _18454_, _18453_);
  and (_18456_, _18455_, _01698_);
  nor (_18457_, _18389_, _01698_);
  or (_18459_, _18457_, _18456_);
  and (_18460_, _18459_, _02082_);
  and (_18461_, _11771_, _03844_);
  nor (_18462_, _18461_, _18355_);
  nor (_18463_, _18462_, _02082_);
  or (_18464_, _18463_, _18460_);
  or (_18465_, _18464_, _39633_);
  or (_18466_, _39632_, \oc8051_golden_model_1.IP [4]);
  and (_18467_, _18466_, _39026_);
  and (_41663_, _18467_, _18465_);
  not (_18469_, \oc8051_golden_model_1.IP [5]);
  nor (_18470_, _03844_, _18469_);
  and (_18471_, _04827_, _03844_);
  nor (_18472_, _18471_, _18470_);
  and (_18473_, _18472_, _01994_);
  nor (_18474_, _04057_, _07925_);
  nor (_18475_, _18474_, _18470_);
  and (_18476_, _18475_, _06188_);
  and (_18477_, _03844_, \oc8051_golden_model_1.ACC [5]);
  nor (_18478_, _18477_, _18470_);
  nor (_18480_, _18478_, _02063_);
  nor (_18481_, _02062_, _18469_);
  or (_18482_, _18481_, _18480_);
  and (_18483_, _18482_, _03006_);
  nor (_18484_, _11804_, _07925_);
  nor (_18485_, _18484_, _18470_);
  nor (_18486_, _18485_, _03006_);
  or (_18487_, _18486_, _18483_);
  and (_18488_, _18487_, _02058_);
  nor (_18489_, _04481_, _18469_);
  and (_18491_, _11789_, _04481_);
  nor (_18492_, _18491_, _18489_);
  nor (_18493_, _18492_, _02058_);
  or (_18494_, _18493_, _18488_);
  and (_18495_, _18494_, _02519_);
  nor (_18496_, _18475_, _02519_);
  or (_18497_, _18496_, _18495_);
  and (_18498_, _18497_, _02549_);
  nor (_18499_, _18478_, _02549_);
  or (_18500_, _18499_, _18498_);
  and (_18502_, _18500_, _02054_);
  and (_18503_, _11816_, _04481_);
  nor (_18504_, _18503_, _18489_);
  nor (_18505_, _18504_, _02054_);
  or (_18506_, _18505_, _18502_);
  and (_18507_, _18506_, _02047_);
  nor (_18508_, _18489_, _11823_);
  nor (_18509_, _18508_, _18492_);
  and (_18510_, _18509_, _02046_);
  or (_18511_, _18510_, _18507_);
  and (_18513_, _18511_, _02043_);
  nor (_18514_, _11841_, _07962_);
  nor (_18515_, _18514_, _18489_);
  nor (_18516_, _18515_, _02043_);
  nor (_18517_, _18516_, _06188_);
  not (_18518_, _18517_);
  nor (_18519_, _18518_, _18513_);
  nor (_18520_, _18519_, _18476_);
  nor (_18521_, _18520_, _02031_);
  and (_18522_, _05258_, _03844_);
  nor (_18524_, _18470_, _02032_);
  not (_18525_, _18524_);
  nor (_18526_, _18525_, _18522_);
  or (_18527_, _18526_, _01765_);
  nor (_18528_, _18527_, _18521_);
  nor (_18529_, _11900_, _07925_);
  nor (_18530_, _18529_, _18470_);
  nor (_18531_, _18530_, _02037_);
  or (_18532_, _18531_, _01994_);
  nor (_18533_, _18532_, _18528_);
  nor (_18535_, _18533_, _18473_);
  or (_18536_, _18535_, _02210_);
  and (_18537_, _11915_, _03844_);
  or (_18538_, _18537_, _18470_);
  or (_18539_, _18538_, _03059_);
  and (_18540_, _18539_, _03061_);
  and (_18541_, _18540_, _18536_);
  and (_18542_, _11786_, _03844_);
  nor (_18543_, _18542_, _18470_);
  nor (_18544_, _18543_, _03061_);
  nor (_18546_, _18544_, _18541_);
  nor (_18547_, _18546_, _02206_);
  nor (_18548_, _18470_, _04104_);
  not (_18549_, _18548_);
  nor (_18550_, _18472_, _02208_);
  and (_18551_, _18550_, _18549_);
  nor (_18552_, _18551_, _18547_);
  nor (_18553_, _18552_, _02342_);
  or (_18554_, _18548_, _03065_);
  nor (_18555_, _18554_, _18478_);
  or (_18557_, _18555_, _02202_);
  nor (_18558_, _18557_, _18553_);
  nor (_18559_, _11913_, _07925_);
  or (_18560_, _18470_, _04953_);
  nor (_18561_, _18560_, _18559_);
  or (_18562_, _18561_, _02334_);
  nor (_18563_, _18562_, _18558_);
  nor (_18564_, _11785_, _07925_);
  nor (_18565_, _18564_, _18470_);
  nor (_18566_, _18565_, _04958_);
  or (_18568_, _18566_, _18563_);
  and (_18569_, _18568_, _02778_);
  nor (_18570_, _18485_, _02778_);
  or (_18571_, _18570_, _18569_);
  and (_18572_, _18571_, _01698_);
  nor (_18573_, _18504_, _01698_);
  or (_18574_, _18573_, _18572_);
  and (_18575_, _18574_, _02082_);
  and (_18576_, _11974_, _03844_);
  nor (_18577_, _18576_, _18470_);
  nor (_18578_, _18577_, _02082_);
  or (_18579_, _18578_, _18575_);
  or (_18580_, _18579_, _39633_);
  or (_18581_, _39632_, \oc8051_golden_model_1.IP [5]);
  and (_18582_, _18581_, _39026_);
  and (_41664_, _18582_, _18580_);
  not (_18583_, \oc8051_golden_model_1.IP [6]);
  nor (_18584_, _03844_, _18583_);
  and (_18585_, _12103_, _03844_);
  nor (_18586_, _18585_, _18584_);
  and (_18588_, _18586_, _01994_);
  nor (_18589_, _03964_, _07925_);
  nor (_18590_, _18589_, _18584_);
  and (_18591_, _18590_, _06188_);
  and (_18592_, _03844_, \oc8051_golden_model_1.ACC [6]);
  nor (_18593_, _18592_, _18584_);
  nor (_18594_, _18593_, _02063_);
  nor (_18595_, _02062_, _18583_);
  or (_18596_, _18595_, _18594_);
  and (_18597_, _18596_, _03006_);
  nor (_18599_, _11993_, _07925_);
  nor (_18600_, _18599_, _18584_);
  nor (_18601_, _18600_, _03006_);
  or (_18602_, _18601_, _18597_);
  and (_18603_, _18602_, _02058_);
  nor (_18604_, _04481_, _18583_);
  and (_18605_, _11990_, _04481_);
  nor (_18606_, _18605_, _18604_);
  nor (_18607_, _18606_, _02058_);
  or (_18608_, _18607_, _18603_);
  and (_18610_, _18608_, _02519_);
  nor (_18611_, _18590_, _02519_);
  or (_18612_, _18611_, _18610_);
  and (_18613_, _18612_, _02549_);
  nor (_18614_, _18593_, _02549_);
  or (_18615_, _18614_, _18613_);
  and (_18616_, _18615_, _02054_);
  and (_18617_, _12017_, _04481_);
  nor (_18618_, _18617_, _18604_);
  nor (_18619_, _18618_, _02054_);
  or (_18621_, _18619_, _18616_);
  and (_18622_, _18621_, _02047_);
  nor (_18623_, _18604_, _12024_);
  nor (_18624_, _18623_, _18606_);
  and (_18625_, _18624_, _02046_);
  or (_18626_, _18625_, _18622_);
  and (_18627_, _18626_, _02043_);
  nor (_18628_, _12042_, _07962_);
  nor (_18629_, _18628_, _18604_);
  nor (_18630_, _18629_, _02043_);
  nor (_18632_, _18630_, _06188_);
  not (_18633_, _18632_);
  nor (_18634_, _18633_, _18627_);
  nor (_18635_, _18634_, _18591_);
  nor (_18636_, _18635_, _02031_);
  and (_18637_, _05029_, _03844_);
  nor (_18638_, _18584_, _02032_);
  not (_18639_, _18638_);
  nor (_18640_, _18639_, _18637_);
  or (_18641_, _18640_, _01765_);
  nor (_18643_, _18641_, _18636_);
  nor (_18644_, _12096_, _07925_);
  nor (_18645_, _18644_, _18584_);
  nor (_18646_, _18645_, _02037_);
  or (_18647_, _18646_, _01994_);
  nor (_18648_, _18647_, _18643_);
  nor (_18649_, _18648_, _18588_);
  or (_18650_, _18649_, _02210_);
  and (_18651_, _12112_, _03844_);
  or (_18652_, _18651_, _18584_);
  or (_18654_, _18652_, _03059_);
  and (_18655_, _18654_, _03061_);
  and (_18656_, _18655_, _18650_);
  and (_18657_, _12118_, _03844_);
  nor (_18658_, _18657_, _18584_);
  nor (_18659_, _18658_, _03061_);
  nor (_18660_, _18659_, _18656_);
  nor (_18661_, _18660_, _02206_);
  nor (_18662_, _18584_, _04011_);
  not (_18663_, _18662_);
  nor (_18665_, _18586_, _02208_);
  and (_18666_, _18665_, _18663_);
  nor (_18667_, _18666_, _18661_);
  nor (_18668_, _18667_, _02342_);
  or (_18669_, _18662_, _03065_);
  nor (_18670_, _18669_, _18593_);
  or (_18671_, _18670_, _02202_);
  nor (_18672_, _18671_, _18668_);
  nor (_18673_, _12110_, _07925_);
  or (_18674_, _18584_, _04953_);
  nor (_18676_, _18674_, _18673_);
  or (_18677_, _18676_, _02334_);
  nor (_18678_, _18677_, _18672_);
  nor (_18679_, _12117_, _07925_);
  nor (_18680_, _18679_, _18584_);
  nor (_18681_, _18680_, _04958_);
  or (_18682_, _18681_, _18678_);
  and (_18683_, _18682_, _02778_);
  nor (_18684_, _18600_, _02778_);
  or (_18685_, _18684_, _18683_);
  and (_18687_, _18685_, _01698_);
  nor (_18688_, _18618_, _01698_);
  or (_18689_, _18688_, _18687_);
  and (_18690_, _18689_, _02082_);
  and (_18691_, _12178_, _03844_);
  nor (_18692_, _18691_, _18584_);
  nor (_18693_, _18692_, _02082_);
  or (_18694_, _18693_, _18690_);
  or (_18695_, _18694_, _39633_);
  or (_18696_, _39632_, \oc8051_golden_model_1.IP [6]);
  and (_18698_, _18696_, _39026_);
  and (_41665_, _18698_, _18695_);
  not (_18699_, \oc8051_golden_model_1.P0 [0]);
  nor (_18700_, _03885_, _18699_);
  and (_18701_, _10792_, _04162_);
  or (_18702_, _18701_, _18700_);
  and (_18703_, _18702_, _02331_);
  and (_18704_, _04162_, _03002_);
  or (_18705_, _18704_, _18700_);
  or (_18706_, _18705_, _05444_);
  nor (_18708_, _04257_, _08034_);
  or (_18709_, _18708_, _18700_);
  or (_18710_, _18709_, _03006_);
  and (_18711_, _03885_, \oc8051_golden_model_1.ACC [0]);
  or (_18712_, _18711_, _18700_);
  and (_18713_, _18712_, _02062_);
  nor (_18714_, _02062_, _18699_);
  or (_18715_, _18714_, _02158_);
  or (_18716_, _18715_, _18713_);
  and (_18717_, _18716_, _02058_);
  and (_18719_, _18717_, _18710_);
  nor (_18720_, _03825_, _18699_);
  and (_18721_, _10814_, _03825_);
  or (_18722_, _18721_, _18720_);
  and (_18723_, _18722_, _02057_);
  or (_18724_, _18723_, _18719_);
  and (_18725_, _18724_, _02519_);
  and (_18726_, _18705_, _02155_);
  or (_18727_, _18726_, _02153_);
  or (_18728_, _18727_, _18725_);
  or (_18730_, _18712_, _02549_);
  and (_18731_, _18730_, _02054_);
  and (_18732_, _18731_, _18728_);
  and (_18733_, _18700_, _02053_);
  or (_18734_, _18733_, _02046_);
  or (_18735_, _18734_, _18732_);
  or (_18736_, _18709_, _02047_);
  and (_18737_, _18736_, _02043_);
  and (_18738_, _18737_, _18735_);
  or (_18739_, _10823_, _10797_);
  and (_18741_, _18739_, _03825_);
  or (_18742_, _18741_, _18720_);
  and (_18743_, _18742_, _02042_);
  or (_18744_, _18743_, _06188_);
  or (_18745_, _18744_, _18738_);
  and (_18746_, _18745_, _18706_);
  or (_18747_, _18746_, _02031_);
  or (_18748_, _18700_, _02032_);
  and (_18749_, _05120_, _03885_);
  or (_18750_, _18749_, _18748_);
  and (_18752_, _18750_, _02037_);
  and (_18753_, _18752_, _18747_);
  and (_18754_, _04882_, \oc8051_golden_model_1.P1 [0]);
  and (_18755_, _04875_, \oc8051_golden_model_1.P0 [0]);
  and (_18756_, _04885_, \oc8051_golden_model_1.P2 [0]);
  and (_18757_, _08088_, \oc8051_golden_model_1.P3 [0]);
  or (_18758_, _18757_, _18756_);
  or (_18759_, _18758_, _18755_);
  or (_18760_, _18759_, _18754_);
  nor (_18761_, _18760_, _10874_);
  and (_18763_, _18761_, _10893_);
  and (_18764_, _18763_, _10873_);
  nand (_18765_, _18764_, _10866_);
  or (_18766_, _18765_, _10852_);
  and (_18767_, _18766_, _03885_);
  or (_18768_, _18767_, _18700_);
  and (_18769_, _18768_, _01765_);
  or (_18770_, _18769_, _18753_);
  or (_18771_, _18770_, _07629_);
  and (_18772_, _10914_, _04162_);
  or (_18774_, _18700_, _03059_);
  or (_18775_, _18774_, _18772_);
  and (_18776_, _03885_, _04837_);
  or (_18777_, _18776_, _18700_);
  or (_18778_, _18777_, _01995_);
  and (_18779_, _18778_, _03061_);
  and (_18780_, _18779_, _18775_);
  and (_18781_, _18780_, _18771_);
  or (_18782_, _18781_, _18703_);
  and (_18783_, _18782_, _02208_);
  nand (_18785_, _18777_, _02206_);
  nor (_18786_, _18785_, _18708_);
  or (_18787_, _18786_, _18783_);
  and (_18788_, _18787_, _03065_);
  or (_18789_, _18700_, _04257_);
  and (_18790_, _18712_, _02342_);
  and (_18791_, _18790_, _18789_);
  or (_18792_, _18791_, _02202_);
  or (_18793_, _18792_, _18788_);
  nor (_18794_, _10913_, _08034_);
  or (_18796_, _18700_, _04953_);
  or (_18797_, _18796_, _18794_);
  and (_18798_, _18797_, _04958_);
  and (_18799_, _18798_, _18793_);
  nor (_18800_, _10789_, _08034_);
  or (_18801_, _18800_, _18700_);
  and (_18802_, _18801_, _02334_);
  or (_18803_, _18802_, _02366_);
  or (_18804_, _18803_, _18799_);
  or (_18805_, _18709_, _02778_);
  and (_18806_, _18805_, _01698_);
  and (_18807_, _18806_, _18804_);
  and (_18808_, _18700_, _01697_);
  or (_18809_, _18808_, _02081_);
  or (_18810_, _18809_, _18807_);
  or (_18811_, _18709_, _02082_);
  and (_18812_, _18811_, _39632_);
  and (_18813_, _18812_, _18810_);
  nor (_18814_, _39632_, _18699_);
  or (_18815_, _18814_, rst);
  or (_41667_, _18815_, _18813_);
  and (_18818_, _08032_, \oc8051_golden_model_1.P0 [1]);
  nor (_18819_, _08034_, _03161_);
  or (_18820_, _18819_, _18818_);
  or (_18821_, _18820_, _02519_);
  or (_18822_, _03885_, \oc8051_golden_model_1.P0 [1]);
  nand (_18823_, _11001_, _04162_);
  and (_18824_, _18823_, _18822_);
  or (_18825_, _18824_, _03006_);
  nand (_18826_, _04162_, _01804_);
  and (_18828_, _18826_, _18822_);
  and (_18829_, _18828_, _02062_);
  and (_18830_, _02063_, \oc8051_golden_model_1.P0 [1]);
  or (_18831_, _18830_, _02158_);
  or (_18832_, _18831_, _18829_);
  and (_18833_, _18832_, _02058_);
  and (_18834_, _18833_, _18825_);
  and (_18835_, _08050_, \oc8051_golden_model_1.P0 [1]);
  and (_18836_, _11005_, _03825_);
  or (_18837_, _18836_, _18835_);
  and (_18839_, _18837_, _02057_);
  or (_18840_, _18839_, _02155_);
  or (_18841_, _18840_, _18834_);
  and (_18842_, _18841_, _18821_);
  or (_18843_, _18842_, _02153_);
  or (_18844_, _18828_, _02549_);
  and (_18845_, _18844_, _02054_);
  and (_18846_, _18845_, _18843_);
  and (_18847_, _10992_, _03825_);
  or (_18848_, _18847_, _18835_);
  and (_18850_, _18848_, _02053_);
  or (_18851_, _18850_, _18846_);
  or (_18852_, _18851_, _02046_);
  or (_18853_, _18835_, _11020_);
  and (_18854_, _18853_, _18837_);
  or (_18855_, _18854_, _02047_);
  and (_18856_, _18855_, _02043_);
  and (_18857_, _18856_, _18852_);
  or (_18858_, _11037_, _10992_);
  and (_18859_, _18858_, _03825_);
  or (_18861_, _18859_, _18835_);
  and (_18862_, _18861_, _02042_);
  or (_18863_, _18862_, _06188_);
  or (_18864_, _18863_, _18857_);
  or (_18865_, _18820_, _05444_);
  and (_18866_, _18865_, _18864_);
  or (_18867_, _18866_, _02031_);
  and (_18868_, _05075_, _03885_);
  or (_18869_, _18818_, _02032_);
  or (_18870_, _18869_, _18868_);
  and (_18872_, _18870_, _02037_);
  and (_18873_, _18872_, _18867_);
  and (_18874_, _18822_, _01765_);
  and (_18875_, _04875_, \oc8051_golden_model_1.P0 [1]);
  and (_18876_, _04882_, \oc8051_golden_model_1.P1 [1]);
  and (_18877_, _04885_, \oc8051_golden_model_1.P2 [1]);
  and (_18878_, _08088_, \oc8051_golden_model_1.P3 [1]);
  or (_18879_, _18878_, _18877_);
  or (_18880_, _18879_, _18876_);
  or (_18881_, _18880_, _18875_);
  nor (_18883_, _18881_, _11072_);
  and (_18884_, _18883_, _11091_);
  and (_18885_, _18884_, _11071_);
  nand (_18886_, _18885_, _11064_);
  or (_18887_, _18886_, _11050_);
  or (_18888_, _18887_, _08034_);
  and (_18889_, _18888_, _18874_);
  or (_18890_, _18889_, _18873_);
  and (_18891_, _18890_, _02212_);
  or (_18892_, _10989_, _08034_);
  and (_18894_, _18892_, _02210_);
  nand (_18895_, _04162_, _02893_);
  and (_18896_, _18895_, _01994_);
  or (_18897_, _18896_, _18894_);
  and (_18898_, _18897_, _18822_);
  or (_18899_, _18898_, _18891_);
  and (_18900_, _18899_, _03061_);
  or (_18901_, _11113_, _08034_);
  and (_18902_, _18822_, _02331_);
  and (_18903_, _18902_, _18901_);
  or (_18905_, _18903_, _18900_);
  and (_18906_, _18905_, _02208_);
  and (_18907_, _10988_, _03885_);
  or (_18908_, _18907_, _18818_);
  and (_18909_, _18908_, _02206_);
  or (_18910_, _18909_, _18906_);
  and (_18911_, _18910_, _03065_);
  or (_18912_, _18818_, _04209_);
  and (_18913_, _18828_, _02342_);
  and (_18914_, _18913_, _18912_);
  or (_18916_, _18914_, _18911_);
  and (_18917_, _18916_, _02335_);
  or (_18918_, _18826_, _04209_);
  and (_18919_, _18822_, _02334_);
  and (_18920_, _18919_, _18918_);
  or (_18921_, _18920_, _02366_);
  or (_18922_, _18895_, _04209_);
  and (_18923_, _18822_, _02202_);
  and (_18924_, _18923_, _18922_);
  or (_18925_, _18924_, _18921_);
  or (_18927_, _18925_, _18917_);
  or (_18928_, _18824_, _02778_);
  and (_18929_, _18928_, _01698_);
  and (_18930_, _18929_, _18927_);
  and (_18931_, _18848_, _01697_);
  or (_18932_, _18931_, _02081_);
  or (_18933_, _18932_, _18930_);
  nor (_18934_, _18818_, _02082_);
  nand (_18935_, _18934_, _18823_);
  and (_18936_, _18935_, _39632_);
  and (_18938_, _18936_, _18933_);
  nor (_18939_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_18940_, _18939_, _00001_);
  or (_41668_, _18940_, _18938_);
  not (_18941_, \oc8051_golden_model_1.P0 [2]);
  nor (_18942_, _03885_, _18941_);
  nor (_18943_, _08034_, _03624_);
  or (_18944_, _18943_, _18942_);
  or (_18945_, _18944_, _05444_);
  nor (_18946_, _11199_, _08034_);
  or (_18948_, _18946_, _18942_);
  or (_18949_, _18948_, _03006_);
  and (_18950_, _03885_, \oc8051_golden_model_1.ACC [2]);
  or (_18951_, _18950_, _18942_);
  and (_18952_, _18951_, _02062_);
  nor (_18953_, _02062_, _18941_);
  or (_18954_, _18953_, _02158_);
  or (_18955_, _18954_, _18952_);
  and (_18956_, _18955_, _02058_);
  and (_18957_, _18956_, _18949_);
  nor (_18959_, _03825_, _18941_);
  and (_18960_, _11194_, _03825_);
  or (_18961_, _18960_, _18959_);
  and (_18962_, _18961_, _02057_);
  or (_18963_, _18962_, _02155_);
  or (_18964_, _18963_, _18957_);
  or (_18965_, _18944_, _02519_);
  and (_18966_, _18965_, _18964_);
  or (_18967_, _18966_, _02153_);
  or (_18968_, _18951_, _02549_);
  and (_18970_, _18968_, _02054_);
  and (_18971_, _18970_, _18967_);
  and (_18972_, _11192_, _03825_);
  or (_18973_, _18972_, _18959_);
  and (_18974_, _18973_, _02053_);
  or (_18975_, _18974_, _02046_);
  or (_18976_, _18975_, _18971_);
  or (_18977_, _18959_, _11223_);
  and (_18978_, _18977_, _18961_);
  or (_18979_, _18978_, _02047_);
  and (_18981_, _18979_, _02043_);
  and (_18982_, _18981_, _18976_);
  or (_18983_, _11240_, _11192_);
  and (_18984_, _18983_, _03825_);
  or (_18985_, _18984_, _18959_);
  and (_18986_, _18985_, _02042_);
  or (_18987_, _18986_, _06188_);
  or (_18988_, _18987_, _18982_);
  and (_18989_, _18988_, _18945_);
  or (_18990_, _18989_, _02031_);
  or (_18992_, _18942_, _02032_);
  and (_18993_, _05211_, _03885_);
  or (_18994_, _18993_, _18992_);
  and (_18995_, _18994_, _02037_);
  and (_18996_, _18995_, _18990_);
  and (_18997_, _04882_, \oc8051_golden_model_1.P1 [2]);
  and (_18998_, _04875_, \oc8051_golden_model_1.P0 [2]);
  and (_18999_, _04885_, \oc8051_golden_model_1.P2 [2]);
  and (_19000_, _08088_, \oc8051_golden_model_1.P3 [2]);
  or (_19001_, _19000_, _18999_);
  or (_19003_, _19001_, _18998_);
  nor (_19004_, _19003_, _18997_);
  and (_19005_, _19004_, _11265_);
  and (_19006_, _19005_, _11279_);
  nand (_19007_, _19006_, _11295_);
  or (_19008_, _19007_, _11253_);
  and (_19009_, _19008_, _03885_);
  or (_19010_, _19009_, _18942_);
  and (_19011_, _19010_, _01765_);
  or (_19012_, _19011_, _18996_);
  or (_19014_, _19012_, _07629_);
  and (_19015_, _11189_, _04162_);
  or (_19016_, _18942_, _03059_);
  or (_19017_, _19016_, _19015_);
  and (_19018_, _03885_, _04866_);
  or (_19019_, _19018_, _18942_);
  or (_19020_, _19019_, _01995_);
  and (_19021_, _19020_, _03061_);
  and (_19022_, _19021_, _19017_);
  and (_19023_, _19022_, _19014_);
  and (_19025_, _11315_, _04162_);
  or (_19026_, _19025_, _18942_);
  and (_19027_, _19026_, _02331_);
  or (_19028_, _19027_, _19023_);
  and (_19029_, _19028_, _02208_);
  or (_19030_, _18942_, _04309_);
  and (_19031_, _19019_, _02206_);
  and (_19032_, _19031_, _19030_);
  or (_19033_, _19032_, _19029_);
  and (_19034_, _19033_, _03065_);
  and (_19036_, _18951_, _02342_);
  and (_19037_, _19036_, _19030_);
  or (_19038_, _19037_, _02202_);
  or (_19039_, _19038_, _19034_);
  nor (_19040_, _11187_, _08034_);
  or (_19041_, _18942_, _04953_);
  or (_19042_, _19041_, _19040_);
  and (_19043_, _19042_, _04958_);
  and (_19044_, _19043_, _19039_);
  nor (_19045_, _11314_, _08034_);
  or (_19047_, _19045_, _18942_);
  and (_19048_, _19047_, _02334_);
  or (_19049_, _19048_, _02366_);
  or (_19050_, _19049_, _19044_);
  or (_19051_, _18948_, _02778_);
  and (_19052_, _19051_, _01698_);
  and (_19053_, _19052_, _19050_);
  and (_19054_, _18973_, _01697_);
  or (_19055_, _19054_, _02081_);
  or (_19056_, _19055_, _19053_);
  and (_19058_, _11367_, _04162_);
  or (_19059_, _18942_, _02082_);
  or (_19060_, _19059_, _19058_);
  and (_19061_, _19060_, _39632_);
  and (_19062_, _19061_, _19056_);
  nor (_19063_, _39632_, _18941_);
  or (_19064_, _19063_, rst);
  or (_41669_, _19064_, _19062_);
  and (_19065_, _08032_, \oc8051_golden_model_1.P0 [3]);
  nor (_19066_, _08034_, _03434_);
  or (_19068_, _19066_, _19065_);
  or (_19069_, _19068_, _05444_);
  or (_19070_, _19068_, _02519_);
  nor (_19071_, _11394_, _08034_);
  or (_19072_, _19071_, _19065_);
  or (_19073_, _19072_, _03006_);
  and (_19074_, _03885_, \oc8051_golden_model_1.ACC [3]);
  or (_19075_, _19074_, _19065_);
  and (_19076_, _19075_, _02062_);
  and (_19077_, _02063_, \oc8051_golden_model_1.P0 [3]);
  or (_19079_, _19077_, _02158_);
  or (_19080_, _19079_, _19076_);
  and (_19081_, _19080_, _02058_);
  and (_19082_, _19081_, _19073_);
  and (_19083_, _08050_, \oc8051_golden_model_1.P0 [3]);
  and (_19084_, _11398_, _03825_);
  or (_19085_, _19084_, _19083_);
  and (_19086_, _19085_, _02057_);
  or (_19087_, _19086_, _02155_);
  or (_19088_, _19087_, _19082_);
  and (_19090_, _19088_, _19070_);
  or (_19091_, _19090_, _02153_);
  or (_19092_, _19075_, _02549_);
  and (_19093_, _19092_, _02054_);
  and (_19094_, _19093_, _19091_);
  and (_19095_, _11408_, _03825_);
  or (_19096_, _19095_, _19083_);
  and (_19097_, _19096_, _02053_);
  or (_19098_, _19097_, _02046_);
  or (_19099_, _19098_, _19094_);
  or (_19101_, _19083_, _11415_);
  and (_19102_, _19101_, _19085_);
  or (_19103_, _19102_, _02047_);
  and (_19104_, _19103_, _02043_);
  and (_19105_, _19104_, _19099_);
  or (_19106_, _11408_, _11431_);
  and (_19107_, _19106_, _03825_);
  or (_19108_, _19107_, _19083_);
  and (_19109_, _19108_, _02042_);
  or (_19110_, _19109_, _06188_);
  or (_19112_, _19110_, _19105_);
  and (_19113_, _19112_, _19069_);
  or (_19114_, _19113_, _02031_);
  or (_19115_, _19065_, _02032_);
  and (_19116_, _05166_, _03885_);
  or (_19117_, _19116_, _19115_);
  and (_19118_, _19117_, _02037_);
  and (_19119_, _19118_, _19114_);
  and (_19120_, _04875_, \oc8051_golden_model_1.P0 [3]);
  and (_19121_, _04882_, \oc8051_golden_model_1.P1 [3]);
  and (_19123_, _04885_, \oc8051_golden_model_1.P2 [3]);
  and (_19124_, _08088_, \oc8051_golden_model_1.P3 [3]);
  or (_19125_, _19124_, _19123_);
  or (_19126_, _19125_, _19121_);
  nor (_19127_, _19126_, _19120_);
  and (_19128_, _19127_, _11457_);
  and (_19129_, _19128_, _11471_);
  nand (_19130_, _19129_, _11487_);
  or (_19131_, _19130_, _11445_);
  and (_19132_, _19131_, _03885_);
  or (_19134_, _19132_, _19065_);
  and (_19135_, _19134_, _01765_);
  or (_19136_, _19135_, _19119_);
  or (_19137_, _19136_, _07629_);
  and (_19138_, _11505_, _04162_);
  or (_19139_, _19065_, _03059_);
  or (_19140_, _19139_, _19138_);
  and (_19141_, _03885_, _04719_);
  or (_19142_, _19141_, _19065_);
  or (_19143_, _19142_, _01995_);
  and (_19145_, _19143_, _03061_);
  and (_19146_, _19145_, _19140_);
  and (_19147_, _19146_, _19137_);
  and (_19148_, _11511_, _04162_);
  or (_19149_, _19148_, _19065_);
  and (_19150_, _19149_, _02331_);
  or (_19151_, _19150_, _19147_);
  and (_19152_, _19151_, _02208_);
  or (_19153_, _19065_, _04153_);
  and (_19154_, _19142_, _02206_);
  and (_19156_, _19154_, _19153_);
  or (_19157_, _19156_, _19152_);
  and (_19158_, _19157_, _03065_);
  and (_19159_, _19075_, _02342_);
  and (_19160_, _19159_, _19153_);
  or (_19161_, _19160_, _02202_);
  or (_19162_, _19161_, _19158_);
  nor (_19163_, _11503_, _08034_);
  or (_19164_, _19065_, _04953_);
  or (_19165_, _19164_, _19163_);
  and (_19167_, _19165_, _04958_);
  and (_19168_, _19167_, _19162_);
  nor (_19169_, _11510_, _08034_);
  or (_19170_, _19169_, _19065_);
  and (_19171_, _19170_, _02334_);
  or (_19172_, _19171_, _02366_);
  or (_19173_, _19172_, _19168_);
  or (_19174_, _19072_, _02778_);
  and (_19175_, _19174_, _01698_);
  and (_19176_, _19175_, _19173_);
  and (_19178_, _19096_, _01697_);
  or (_19179_, _19178_, _02081_);
  or (_19180_, _19179_, _19176_);
  and (_19181_, _11567_, _04162_);
  or (_19182_, _19065_, _02082_);
  or (_19183_, _19182_, _19181_);
  and (_19184_, _19183_, _39632_);
  and (_19185_, _19184_, _19180_);
  nor (_19186_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_19187_, _19186_, _00001_);
  or (_41670_, _19187_, _19185_);
  not (_19189_, \oc8051_golden_model_1.P0 [4]);
  nor (_19190_, _03885_, _19189_);
  nor (_19191_, _04372_, _08034_);
  or (_19192_, _19191_, _19190_);
  or (_19193_, _19192_, _05444_);
  or (_19194_, _19192_, _02519_);
  nor (_19195_, _11611_, _08034_);
  or (_19196_, _19195_, _19190_);
  or (_19197_, _19196_, _03006_);
  and (_19199_, _03885_, \oc8051_golden_model_1.ACC [4]);
  or (_19200_, _19199_, _19190_);
  and (_19201_, _19200_, _02062_);
  nor (_19202_, _02062_, _19189_);
  or (_19203_, _19202_, _02158_);
  or (_19204_, _19203_, _19201_);
  and (_19205_, _19204_, _02058_);
  and (_19206_, _19205_, _19197_);
  nor (_19207_, _03825_, _19189_);
  and (_19208_, _11597_, _03825_);
  or (_19210_, _19208_, _19207_);
  and (_19211_, _19210_, _02057_);
  or (_19212_, _19211_, _02155_);
  or (_19213_, _19212_, _19206_);
  and (_19214_, _19213_, _19194_);
  or (_19215_, _19214_, _02153_);
  or (_19216_, _19200_, _02549_);
  and (_19217_, _19216_, _02054_);
  and (_19218_, _19217_, _19215_);
  and (_19219_, _11595_, _03825_);
  or (_19221_, _19219_, _19207_);
  and (_19222_, _19221_, _02053_);
  or (_19223_, _19222_, _02046_);
  or (_19224_, _19223_, _19218_);
  or (_19225_, _19207_, _11628_);
  and (_19226_, _19225_, _19210_);
  or (_19227_, _19226_, _02047_);
  and (_19228_, _19227_, _02043_);
  and (_19229_, _19228_, _19224_);
  or (_19230_, _11645_, _11595_);
  and (_19232_, _19230_, _03825_);
  or (_19233_, _19232_, _19207_);
  and (_19234_, _19233_, _02042_);
  or (_19235_, _19234_, _06188_);
  or (_19236_, _19235_, _19229_);
  and (_19237_, _19236_, _19193_);
  or (_19238_, _19237_, _02031_);
  or (_19239_, _19190_, _02032_);
  and (_19240_, _05303_, _03885_);
  or (_19241_, _19240_, _19239_);
  and (_19243_, _19241_, _02037_);
  and (_19244_, _19243_, _19238_);
  and (_19245_, _04882_, \oc8051_golden_model_1.P1 [4]);
  and (_19246_, _04875_, \oc8051_golden_model_1.P0 [4]);
  and (_19247_, _04885_, \oc8051_golden_model_1.P2 [4]);
  and (_19248_, _08088_, \oc8051_golden_model_1.P3 [4]);
  or (_19249_, _19248_, _19247_);
  or (_19250_, _19249_, _19246_);
  or (_19251_, _19250_, _19245_);
  nor (_19252_, _19251_, _11680_);
  and (_19254_, _19252_, _11699_);
  and (_19255_, _19254_, _11679_);
  nand (_19256_, _19255_, _11672_);
  or (_19257_, _19256_, _11658_);
  and (_19258_, _19257_, _03885_);
  or (_19259_, _19258_, _19190_);
  and (_19260_, _19259_, _01765_);
  or (_19261_, _19260_, _19244_);
  or (_19262_, _19261_, _07629_);
  and (_19263_, _11592_, _04162_);
  or (_19265_, _19190_, _03059_);
  or (_19266_, _19265_, _19263_);
  and (_19267_, _04831_, _03885_);
  or (_19268_, _19267_, _19190_);
  or (_19269_, _19268_, _01995_);
  and (_19270_, _19269_, _03061_);
  and (_19271_, _19270_, _19266_);
  and (_19272_, _19271_, _19262_);
  and (_19273_, _11588_, _04162_);
  or (_19274_, _19273_, _19190_);
  and (_19276_, _19274_, _02331_);
  or (_19277_, _19276_, _19272_);
  and (_19278_, _19277_, _02208_);
  or (_19279_, _19190_, _04420_);
  and (_19280_, _19268_, _02206_);
  and (_19281_, _19280_, _19279_);
  or (_19282_, _19281_, _19278_);
  and (_19283_, _19282_, _03065_);
  and (_19284_, _19200_, _02342_);
  and (_19285_, _19284_, _19279_);
  or (_19287_, _19285_, _02202_);
  or (_19288_, _19287_, _19283_);
  nor (_19289_, _11590_, _08034_);
  or (_19290_, _19190_, _04953_);
  or (_19291_, _19290_, _19289_);
  and (_19292_, _19291_, _04958_);
  and (_19293_, _19292_, _19288_);
  nor (_19294_, _11587_, _08034_);
  or (_19295_, _19294_, _19190_);
  and (_19296_, _19295_, _02334_);
  or (_19298_, _19296_, _02366_);
  or (_19299_, _19298_, _19293_);
  or (_19300_, _19196_, _02778_);
  and (_19301_, _19300_, _01698_);
  and (_19302_, _19301_, _19299_);
  and (_19303_, _19221_, _01697_);
  or (_19304_, _19303_, _02081_);
  or (_19305_, _19304_, _19302_);
  and (_19306_, _11771_, _04162_);
  or (_19307_, _19190_, _02082_);
  or (_19309_, _19307_, _19306_);
  and (_19310_, _19309_, _39632_);
  and (_19311_, _19310_, _19305_);
  nor (_19312_, _39632_, _19189_);
  or (_19313_, _19312_, rst);
  or (_41671_, _19313_, _19311_);
  not (_19314_, \oc8051_golden_model_1.P0 [5]);
  nor (_19315_, _03885_, _19314_);
  nor (_19316_, _04057_, _08034_);
  or (_19317_, _19316_, _19315_);
  or (_19320_, _19317_, _05444_);
  or (_19321_, _19317_, _02519_);
  nor (_19322_, _11804_, _08034_);
  or (_19323_, _19322_, _19315_);
  or (_19324_, _19323_, _03006_);
  and (_19325_, _03885_, \oc8051_golden_model_1.ACC [5]);
  or (_19326_, _19325_, _19315_);
  and (_19327_, _19326_, _02062_);
  nor (_19328_, _02062_, _19314_);
  or (_19329_, _19328_, _02158_);
  or (_19331_, _19329_, _19327_);
  and (_19332_, _19331_, _02058_);
  and (_19333_, _19332_, _19324_);
  nor (_19334_, _03825_, _19314_);
  and (_19335_, _11789_, _03825_);
  or (_19336_, _19335_, _19334_);
  and (_19337_, _19336_, _02057_);
  or (_19338_, _19337_, _02155_);
  or (_19339_, _19338_, _19333_);
  and (_19340_, _19339_, _19321_);
  or (_19343_, _19340_, _02153_);
  or (_19344_, _19326_, _02549_);
  and (_19345_, _19344_, _02054_);
  and (_19346_, _19345_, _19343_);
  and (_19347_, _11816_, _03825_);
  or (_19348_, _19347_, _19334_);
  and (_19349_, _19348_, _02053_);
  or (_19350_, _19349_, _02046_);
  or (_19351_, _19350_, _19346_);
  or (_19352_, _19334_, _11823_);
  and (_19354_, _19352_, _19336_);
  or (_19355_, _19354_, _02047_);
  and (_19356_, _19355_, _02043_);
  and (_19357_, _19356_, _19351_);
  or (_19358_, _11840_, _11816_);
  and (_19359_, _19358_, _03825_);
  or (_19360_, _19359_, _19334_);
  and (_19361_, _19360_, _02042_);
  or (_19362_, _19361_, _06188_);
  or (_19363_, _19362_, _19357_);
  and (_19366_, _19363_, _19320_);
  or (_19367_, _19366_, _02031_);
  or (_19368_, _19315_, _02032_);
  and (_19369_, _05258_, _03885_);
  or (_19370_, _19369_, _19368_);
  and (_19371_, _19370_, _02037_);
  and (_19372_, _19371_, _19367_);
  nor (_19373_, _11863_, _11861_);
  and (_19374_, _04879_, \oc8051_golden_model_1.P3 [5]);
  nor (_19375_, _19374_, _11882_);
  and (_19377_, _19375_, _19373_);
  nand (_19378_, _19377_, _11860_);
  not (_19379_, _11885_);
  and (_19380_, _11891_, _19379_);
  nand (_19381_, _19380_, _11880_);
  nor (_19382_, _11886_, _11883_);
  nand (_19383_, _19382_, _11894_);
  and (_19384_, _04885_, \oc8051_golden_model_1.P2 [5]);
  and (_19385_, _04882_, \oc8051_golden_model_1.P1 [5]);
  and (_19386_, _11864_, \oc8051_golden_model_1.P0 [5]);
  or (_19389_, _19386_, _19385_);
  or (_19390_, _19389_, _19384_);
  or (_19391_, _19390_, _19383_);
  or (_19392_, _19391_, _19381_);
  or (_19393_, _19392_, _19378_);
  or (_19394_, _19393_, _11853_);
  and (_19395_, _19394_, _03885_);
  or (_19396_, _19395_, _19315_);
  and (_19397_, _19396_, _01765_);
  or (_19398_, _19397_, _19372_);
  or (_19400_, _19398_, _07629_);
  and (_19401_, _11915_, _04162_);
  or (_19402_, _19315_, _03059_);
  or (_19403_, _19402_, _19401_);
  and (_19404_, _04827_, _03885_);
  or (_19405_, _19404_, _19315_);
  or (_19406_, _19405_, _01995_);
  and (_19407_, _19406_, _03061_);
  and (_19408_, _19407_, _19403_);
  and (_19409_, _19408_, _19400_);
  and (_19411_, _11786_, _04162_);
  or (_19412_, _19411_, _19315_);
  and (_19413_, _19412_, _02331_);
  or (_19414_, _19413_, _19409_);
  and (_19415_, _19414_, _02208_);
  or (_19416_, _19315_, _04104_);
  and (_19417_, _19405_, _02206_);
  and (_19418_, _19417_, _19416_);
  or (_19419_, _19418_, _19415_);
  and (_19420_, _19419_, _03065_);
  and (_19422_, _19326_, _02342_);
  and (_19423_, _19422_, _19416_);
  or (_19424_, _19423_, _02202_);
  or (_19425_, _19424_, _19420_);
  nor (_19426_, _11913_, _08034_);
  or (_19427_, _19315_, _04953_);
  or (_19428_, _19427_, _19426_);
  and (_19429_, _19428_, _04958_);
  and (_19430_, _19429_, _19425_);
  nor (_19431_, _11785_, _08034_);
  or (_19433_, _19431_, _19315_);
  and (_19434_, _19433_, _02334_);
  or (_19435_, _19434_, _02366_);
  or (_19436_, _19435_, _19430_);
  or (_19437_, _19323_, _02778_);
  and (_19438_, _19437_, _01698_);
  and (_19439_, _19438_, _19436_);
  and (_19440_, _19348_, _01697_);
  or (_19441_, _19440_, _02081_);
  or (_19442_, _19441_, _19439_);
  and (_19444_, _11974_, _04162_);
  or (_19445_, _19315_, _02082_);
  or (_19446_, _19445_, _19444_);
  and (_19447_, _19446_, _39632_);
  and (_19448_, _19447_, _19442_);
  nor (_19449_, _39632_, _19314_);
  or (_19450_, _19449_, rst);
  or (_41672_, _19450_, _19448_);
  not (_19451_, \oc8051_golden_model_1.P0 [6]);
  nor (_19452_, _03885_, _19451_);
  nor (_19454_, _03964_, _08034_);
  or (_19455_, _19454_, _19452_);
  or (_19456_, _19455_, _05444_);
  or (_19457_, _19455_, _02519_);
  nor (_19458_, _11993_, _08034_);
  or (_19459_, _19458_, _19452_);
  or (_19460_, _19459_, _03006_);
  and (_19461_, _03885_, \oc8051_golden_model_1.ACC [6]);
  or (_19462_, _19461_, _19452_);
  and (_19463_, _19462_, _02062_);
  nor (_19465_, _02062_, _19451_);
  or (_19466_, _19465_, _02158_);
  or (_19467_, _19466_, _19463_);
  and (_19468_, _19467_, _02058_);
  and (_19469_, _19468_, _19460_);
  nor (_19470_, _03825_, _19451_);
  and (_19471_, _11990_, _03825_);
  or (_19472_, _19471_, _19470_);
  and (_19473_, _19472_, _02057_);
  or (_19474_, _19473_, _02155_);
  or (_19476_, _19474_, _19469_);
  and (_19477_, _19476_, _19457_);
  or (_19478_, _19477_, _02153_);
  or (_19479_, _19462_, _02549_);
  and (_19480_, _19479_, _02054_);
  and (_19481_, _19480_, _19478_);
  and (_19482_, _12017_, _03825_);
  or (_19483_, _19482_, _19470_);
  and (_19484_, _19483_, _02053_);
  or (_19485_, _19484_, _02046_);
  or (_19487_, _19485_, _19481_);
  or (_19488_, _19470_, _12024_);
  and (_19489_, _19488_, _19472_);
  or (_19490_, _19489_, _02047_);
  and (_19491_, _19490_, _02043_);
  and (_19492_, _19491_, _19487_);
  or (_19493_, _12041_, _12017_);
  and (_19494_, _19493_, _03825_);
  or (_19495_, _19494_, _19470_);
  and (_19496_, _19495_, _02042_);
  or (_19498_, _19496_, _06188_);
  or (_19499_, _19498_, _19492_);
  and (_19500_, _19499_, _19456_);
  or (_19501_, _19500_, _02031_);
  or (_19502_, _19452_, _02032_);
  and (_19503_, _05029_, _03885_);
  or (_19504_, _19503_, _19502_);
  and (_19505_, _19504_, _02037_);
  and (_19506_, _19505_, _19501_);
  and (_19507_, _04882_, \oc8051_golden_model_1.P1 [6]);
  and (_19509_, _04875_, \oc8051_golden_model_1.P0 [6]);
  and (_19510_, _04885_, \oc8051_golden_model_1.P2 [6]);
  and (_19511_, _08088_, \oc8051_golden_model_1.P3 [6]);
  or (_19512_, _19511_, _19510_);
  or (_19513_, _19512_, _19509_);
  or (_19514_, _19513_, _19507_);
  or (_19515_, _19514_, _12091_);
  or (_19516_, _19515_, _12081_);
  or (_19517_, _19516_, _12076_);
  or (_19518_, _19517_, _12069_);
  or (_19520_, _19518_, _12054_);
  and (_19521_, _19520_, _03885_);
  or (_19522_, _19521_, _19452_);
  and (_19523_, _19522_, _01765_);
  or (_19524_, _19523_, _19506_);
  or (_19525_, _19524_, _07629_);
  and (_19526_, _12112_, _04162_);
  or (_19527_, _19452_, _03059_);
  or (_19528_, _19527_, _19526_);
  and (_19529_, _12103_, _03885_);
  or (_19531_, _19529_, _19452_);
  or (_19532_, _19531_, _01995_);
  and (_19533_, _19532_, _03061_);
  and (_19534_, _19533_, _19528_);
  and (_19535_, _19534_, _19525_);
  and (_19536_, _12118_, _04162_);
  or (_19537_, _19536_, _19452_);
  and (_19538_, _19537_, _02331_);
  or (_19539_, _19538_, _19535_);
  and (_19540_, _19539_, _02208_);
  or (_19542_, _19452_, _04011_);
  and (_19543_, _19531_, _02206_);
  and (_19544_, _19543_, _19542_);
  or (_19545_, _19544_, _19540_);
  and (_19546_, _19545_, _03065_);
  and (_19547_, _19462_, _02342_);
  and (_19548_, _19547_, _19542_);
  or (_19549_, _19548_, _02202_);
  or (_19550_, _19549_, _19546_);
  nor (_19551_, _12110_, _08034_);
  or (_19553_, _19452_, _04953_);
  or (_19554_, _19553_, _19551_);
  and (_19555_, _19554_, _04958_);
  and (_19556_, _19555_, _19550_);
  nor (_19557_, _12117_, _08034_);
  or (_19558_, _19557_, _19452_);
  and (_19559_, _19558_, _02334_);
  or (_19560_, _19559_, _02366_);
  or (_19561_, _19560_, _19556_);
  or (_19562_, _19459_, _02778_);
  and (_19564_, _19562_, _01698_);
  and (_19565_, _19564_, _19561_);
  and (_19566_, _19483_, _01697_);
  or (_19567_, _19566_, _02081_);
  or (_19568_, _19567_, _19565_);
  and (_19569_, _12178_, _04162_);
  or (_19570_, _19452_, _02082_);
  or (_19571_, _19570_, _19569_);
  and (_19572_, _19571_, _39632_);
  and (_19573_, _19572_, _19568_);
  nor (_19575_, _39632_, _19451_);
  or (_19576_, _19575_, rst);
  or (_41674_, _19576_, _19573_);
  not (_19577_, \oc8051_golden_model_1.P1 [0]);
  nor (_19578_, _03859_, _19577_);
  and (_19579_, _10792_, _03859_);
  or (_19580_, _19579_, _19578_);
  and (_19581_, _19580_, _02331_);
  and (_19582_, _03859_, _03002_);
  or (_19583_, _19582_, _19578_);
  or (_19585_, _19583_, _05444_);
  nor (_19586_, _04257_, _08149_);
  or (_19587_, _19586_, _19578_);
  or (_19588_, _19587_, _03006_);
  and (_19589_, _03859_, \oc8051_golden_model_1.ACC [0]);
  or (_19590_, _19589_, _19578_);
  and (_19591_, _19590_, _02062_);
  nor (_19592_, _02062_, _19577_);
  or (_19593_, _19592_, _02158_);
  or (_19594_, _19593_, _19591_);
  and (_19596_, _19594_, _02058_);
  and (_19597_, _19596_, _19588_);
  nor (_19598_, _04489_, _19577_);
  and (_19599_, _10814_, _04489_);
  or (_19600_, _19599_, _19598_);
  and (_19601_, _19600_, _02057_);
  or (_19602_, _19601_, _19597_);
  and (_19603_, _19602_, _02519_);
  and (_19604_, _19583_, _02155_);
  or (_19605_, _19604_, _02153_);
  or (_19607_, _19605_, _19603_);
  or (_19608_, _19590_, _02549_);
  and (_19609_, _19608_, _02054_);
  and (_19610_, _19609_, _19607_);
  and (_19611_, _19578_, _02053_);
  or (_19612_, _19611_, _02046_);
  or (_19613_, _19612_, _19610_);
  or (_19614_, _19587_, _02047_);
  and (_19615_, _19614_, _02043_);
  and (_19616_, _19615_, _19613_);
  and (_19618_, _18739_, _04489_);
  or (_19619_, _19618_, _19598_);
  and (_19620_, _19619_, _02042_);
  or (_19621_, _19620_, _06188_);
  or (_19622_, _19621_, _19616_);
  and (_19623_, _19622_, _19585_);
  or (_19624_, _19623_, _02031_);
  and (_19625_, _05120_, _03859_);
  or (_19626_, _19578_, _02032_);
  or (_19627_, _19626_, _19625_);
  and (_19629_, _19627_, _02037_);
  and (_19630_, _19629_, _19624_);
  and (_19631_, _18766_, _03859_);
  or (_19632_, _19631_, _19578_);
  and (_19633_, _19632_, _01765_);
  or (_19634_, _19633_, _19630_);
  or (_19635_, _19634_, _07629_);
  and (_19636_, _10914_, _03859_);
  or (_19637_, _19578_, _03059_);
  or (_19638_, _19637_, _19636_);
  and (_19640_, _03859_, _04837_);
  or (_19641_, _19640_, _19578_);
  or (_19642_, _19641_, _01995_);
  and (_19643_, _19642_, _03061_);
  and (_19644_, _19643_, _19638_);
  and (_19645_, _19644_, _19635_);
  or (_19646_, _19645_, _19581_);
  and (_19647_, _19646_, _02208_);
  nand (_19648_, _19641_, _02206_);
  nor (_19649_, _19648_, _19586_);
  or (_19651_, _19649_, _19647_);
  and (_19652_, _19651_, _03065_);
  or (_19653_, _19578_, _04257_);
  and (_19654_, _19590_, _02342_);
  and (_19655_, _19654_, _19653_);
  or (_19656_, _19655_, _02202_);
  or (_19657_, _19656_, _19652_);
  nor (_19658_, _10913_, _08149_);
  or (_19659_, _19578_, _04953_);
  or (_19660_, _19659_, _19658_);
  and (_19662_, _19660_, _04958_);
  and (_19663_, _19662_, _19657_);
  nor (_19664_, _10789_, _08149_);
  or (_19665_, _19664_, _19578_);
  and (_19666_, _19665_, _02334_);
  or (_19667_, _19666_, _02366_);
  or (_19668_, _19667_, _19663_);
  or (_19669_, _19587_, _02778_);
  and (_19670_, _19669_, _01698_);
  and (_19671_, _19670_, _19668_);
  and (_19673_, _19578_, _01697_);
  or (_19674_, _19673_, _02081_);
  or (_19675_, _19674_, _19671_);
  or (_19676_, _19587_, _02082_);
  and (_19677_, _19676_, _39632_);
  and (_19678_, _19677_, _19675_);
  nor (_19679_, _39632_, _19577_);
  or (_19680_, _19679_, rst);
  or (_41675_, _19680_, _19678_);
  nor (_19681_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_19683_, _19681_, _00001_);
  and (_19684_, _08149_, \oc8051_golden_model_1.P1 [1]);
  nor (_19685_, _08149_, _03161_);
  or (_19686_, _19685_, _19684_);
  or (_19687_, _19686_, _02519_);
  or (_19688_, _03859_, \oc8051_golden_model_1.P1 [1]);
  and (_19689_, _11001_, _03859_);
  not (_19690_, _19689_);
  and (_19691_, _19690_, _19688_);
  or (_19692_, _19691_, _03006_);
  nand (_19694_, _03859_, _01804_);
  and (_19695_, _19694_, _19688_);
  and (_19696_, _19695_, _02062_);
  and (_19697_, _02063_, \oc8051_golden_model_1.P1 [1]);
  or (_19698_, _19697_, _02158_);
  or (_19699_, _19698_, _19696_);
  and (_19700_, _19699_, _02058_);
  and (_19701_, _19700_, _19692_);
  not (_19702_, _04489_);
  and (_19703_, _19702_, \oc8051_golden_model_1.P1 [1]);
  and (_19705_, _11005_, _04489_);
  or (_19706_, _19705_, _19703_);
  and (_19707_, _19706_, _02057_);
  or (_19708_, _19707_, _02155_);
  or (_19709_, _19708_, _19701_);
  and (_19710_, _19709_, _19687_);
  or (_19711_, _19710_, _02153_);
  or (_19712_, _19695_, _02549_);
  and (_19713_, _19712_, _02054_);
  and (_19714_, _19713_, _19711_);
  and (_19716_, _10992_, _04489_);
  or (_19717_, _19716_, _19703_);
  and (_19718_, _19717_, _02053_);
  or (_19719_, _19718_, _19714_);
  or (_19720_, _19719_, _02046_);
  or (_19721_, _19703_, _11020_);
  and (_19722_, _19721_, _19706_);
  or (_19723_, _19722_, _02047_);
  and (_19724_, _19723_, _02043_);
  and (_19725_, _19724_, _19720_);
  and (_19727_, _18858_, _04489_);
  or (_19728_, _19727_, _19703_);
  and (_19729_, _19728_, _02042_);
  or (_19730_, _19729_, _06188_);
  or (_19731_, _19730_, _19725_);
  or (_19732_, _19686_, _05444_);
  and (_19733_, _19732_, _19731_);
  or (_19734_, _19733_, _02031_);
  and (_19735_, _05075_, _03859_);
  or (_19736_, _19684_, _02032_);
  or (_19738_, _19736_, _19735_);
  and (_19739_, _19738_, _02037_);
  and (_19740_, _19739_, _19734_);
  and (_19741_, _18887_, _03859_);
  or (_19742_, _19741_, _19684_);
  and (_19743_, _19742_, _01765_);
  or (_19744_, _19743_, _19740_);
  and (_19745_, _19744_, _02212_);
  or (_19746_, _10989_, _08149_);
  and (_19747_, _19746_, _02210_);
  nand (_19749_, _03859_, _02893_);
  and (_19750_, _19749_, _01994_);
  or (_19751_, _19750_, _19747_);
  and (_19752_, _19751_, _19688_);
  or (_19753_, _19752_, _19745_);
  and (_19754_, _19753_, _03061_);
  or (_19755_, _11113_, _08149_);
  and (_19756_, _19688_, _02331_);
  and (_19757_, _19756_, _19755_);
  or (_19758_, _19757_, _19754_);
  and (_19760_, _19758_, _02208_);
  or (_19761_, _10988_, _08149_);
  and (_19762_, _19688_, _02206_);
  and (_19763_, _19762_, _19761_);
  or (_19764_, _19763_, _19760_);
  and (_19765_, _19764_, _03065_);
  or (_19766_, _19684_, _04209_);
  and (_19767_, _19695_, _02342_);
  and (_19768_, _19767_, _19766_);
  or (_19769_, _19768_, _19765_);
  and (_19771_, _19769_, _02335_);
  or (_19772_, _19694_, _04209_);
  and (_19773_, _19688_, _02334_);
  and (_19774_, _19773_, _19772_);
  or (_19775_, _19774_, _02366_);
  or (_19776_, _19749_, _04209_);
  and (_19777_, _19688_, _02202_);
  and (_19778_, _19777_, _19776_);
  or (_19779_, _19778_, _19775_);
  or (_19780_, _19779_, _19771_);
  or (_19782_, _19691_, _02778_);
  and (_19783_, _19782_, _01698_);
  and (_19784_, _19783_, _19780_);
  and (_19785_, _19717_, _01697_);
  or (_19786_, _19785_, _02081_);
  or (_19787_, _19786_, _19784_);
  or (_19788_, _19684_, _02082_);
  or (_19789_, _19788_, _19689_);
  and (_19790_, _19789_, _39632_);
  and (_19791_, _19790_, _19787_);
  or (_41676_, _19791_, _19683_);
  not (_19793_, \oc8051_golden_model_1.P1 [2]);
  nor (_19794_, _03859_, _19793_);
  nor (_19795_, _08149_, _03624_);
  or (_19796_, _19795_, _19794_);
  or (_19797_, _19796_, _05444_);
  nor (_19798_, _11199_, _08149_);
  or (_19799_, _19798_, _19794_);
  and (_19800_, _19799_, _02158_);
  nor (_19801_, _02062_, _19793_);
  and (_19803_, _03859_, \oc8051_golden_model_1.ACC [2]);
  or (_19804_, _19803_, _19794_);
  and (_19805_, _19804_, _02062_);
  or (_19806_, _19805_, _19801_);
  and (_19807_, _19806_, _03006_);
  or (_19808_, _19807_, _02057_);
  or (_19809_, _19808_, _19800_);
  nor (_19810_, _04489_, _19793_);
  and (_19811_, _11194_, _04489_);
  or (_19812_, _19811_, _19810_);
  or (_19814_, _19812_, _02058_);
  and (_19815_, _19814_, _19809_);
  or (_19816_, _19815_, _02155_);
  or (_19817_, _19796_, _02519_);
  and (_19818_, _19817_, _19816_);
  or (_19819_, _19818_, _02153_);
  or (_19820_, _19804_, _02549_);
  and (_19821_, _19820_, _02054_);
  and (_19822_, _19821_, _19819_);
  and (_19823_, _11192_, _04489_);
  or (_19825_, _19823_, _19810_);
  and (_19826_, _19825_, _02053_);
  or (_19827_, _19826_, _02046_);
  or (_19828_, _19827_, _19822_);
  or (_19829_, _19810_, _11223_);
  and (_19830_, _19829_, _19812_);
  or (_19831_, _19830_, _02047_);
  and (_19832_, _19831_, _02043_);
  and (_19833_, _19832_, _19828_);
  and (_19834_, _18983_, _04489_);
  or (_19836_, _19834_, _19810_);
  and (_19837_, _19836_, _02042_);
  or (_19838_, _19837_, _06188_);
  or (_19839_, _19838_, _19833_);
  and (_19840_, _19839_, _19797_);
  or (_19841_, _19840_, _02031_);
  and (_19842_, _05211_, _03859_);
  or (_19843_, _19794_, _02032_);
  or (_19844_, _19843_, _19842_);
  and (_19845_, _19844_, _02037_);
  and (_19847_, _19845_, _19841_);
  and (_19848_, _19008_, _03859_);
  or (_19849_, _19794_, _19848_);
  and (_19850_, _19849_, _01765_);
  or (_19851_, _19850_, _19847_);
  or (_19852_, _19851_, _07629_);
  and (_19853_, _11189_, _03859_);
  or (_19854_, _19794_, _03059_);
  or (_19855_, _19854_, _19853_);
  and (_19856_, _03859_, _04866_);
  or (_19858_, _19856_, _19794_);
  or (_19859_, _19858_, _01995_);
  and (_19860_, _19859_, _03061_);
  and (_19861_, _19860_, _19855_);
  and (_19862_, _19861_, _19852_);
  and (_19863_, _11315_, _03859_);
  or (_19864_, _19863_, _19794_);
  and (_19865_, _19864_, _02331_);
  or (_19866_, _19865_, _19862_);
  and (_19867_, _19866_, _02208_);
  or (_19869_, _19794_, _04309_);
  and (_19870_, _19858_, _02206_);
  and (_19871_, _19870_, _19869_);
  or (_19872_, _19871_, _19867_);
  and (_19873_, _19872_, _03065_);
  and (_19874_, _19804_, _02342_);
  and (_19875_, _19874_, _19869_);
  or (_19876_, _19875_, _02202_);
  or (_19877_, _19876_, _19873_);
  nor (_19878_, _11187_, _08149_);
  or (_19880_, _19794_, _04953_);
  or (_19881_, _19880_, _19878_);
  and (_19882_, _19881_, _04958_);
  and (_19883_, _19882_, _19877_);
  nor (_19884_, _11314_, _08149_);
  or (_19885_, _19884_, _19794_);
  and (_19886_, _19885_, _02334_);
  or (_19887_, _19886_, _02366_);
  or (_19888_, _19887_, _19883_);
  or (_19889_, _19799_, _02778_);
  and (_19891_, _19889_, _01698_);
  and (_19892_, _19891_, _19888_);
  and (_19893_, _19825_, _01697_);
  or (_19894_, _19893_, _02081_);
  or (_19895_, _19894_, _19892_);
  and (_19896_, _11367_, _03859_);
  or (_19897_, _19794_, _02082_);
  or (_19898_, _19897_, _19896_);
  and (_19899_, _19898_, _39632_);
  and (_19900_, _19899_, _19895_);
  nor (_19902_, _39632_, _19793_);
  or (_19903_, _19902_, rst);
  or (_41678_, _19903_, _19900_);
  and (_19904_, _08149_, \oc8051_golden_model_1.P1 [3]);
  nor (_19905_, _08149_, _03434_);
  or (_19906_, _19905_, _19904_);
  or (_19907_, _19906_, _05444_);
  or (_19908_, _19906_, _02519_);
  nor (_19909_, _11394_, _08149_);
  or (_19910_, _19909_, _19904_);
  or (_19912_, _19910_, _03006_);
  and (_19913_, _03859_, \oc8051_golden_model_1.ACC [3]);
  or (_19914_, _19913_, _19904_);
  and (_19915_, _19914_, _02062_);
  and (_19916_, _02063_, \oc8051_golden_model_1.P1 [3]);
  or (_19917_, _19916_, _02158_);
  or (_19918_, _19917_, _19915_);
  and (_19919_, _19918_, _02058_);
  and (_19920_, _19919_, _19912_);
  and (_19921_, _19702_, \oc8051_golden_model_1.P1 [3]);
  and (_19923_, _11398_, _04489_);
  or (_19924_, _19923_, _19921_);
  and (_19925_, _19924_, _02057_);
  or (_19926_, _19925_, _02155_);
  or (_19927_, _19926_, _19920_);
  and (_19928_, _19927_, _19908_);
  or (_19929_, _19928_, _02153_);
  or (_19930_, _19914_, _02549_);
  and (_19931_, _19930_, _02054_);
  and (_19932_, _19931_, _19929_);
  and (_19934_, _11408_, _04489_);
  or (_19935_, _19934_, _19921_);
  and (_19936_, _19935_, _02053_);
  or (_19937_, _19936_, _02046_);
  or (_19938_, _19937_, _19932_);
  or (_19939_, _19921_, _11415_);
  and (_19940_, _19939_, _19924_);
  or (_19941_, _19940_, _02047_);
  and (_19942_, _19941_, _02043_);
  and (_19943_, _19942_, _19938_);
  and (_19945_, _19106_, _04489_);
  or (_19946_, _19945_, _19921_);
  and (_19947_, _19946_, _02042_);
  or (_19948_, _19947_, _06188_);
  or (_19949_, _19948_, _19943_);
  and (_19950_, _19949_, _19907_);
  or (_19951_, _19950_, _02031_);
  and (_19952_, _05166_, _03859_);
  or (_19953_, _19904_, _02032_);
  or (_19954_, _19953_, _19952_);
  and (_19956_, _19954_, _02037_);
  and (_19957_, _19956_, _19951_);
  and (_19958_, _19131_, _03859_);
  or (_19959_, _19904_, _19958_);
  and (_19960_, _19959_, _01765_);
  or (_19961_, _19960_, _19957_);
  or (_19962_, _19961_, _07629_);
  and (_19963_, _11505_, _03859_);
  or (_19964_, _19904_, _03059_);
  or (_19965_, _19964_, _19963_);
  and (_19967_, _03859_, _04719_);
  or (_19968_, _19967_, _19904_);
  or (_19969_, _19968_, _01995_);
  and (_19970_, _19969_, _03061_);
  and (_19971_, _19970_, _19965_);
  and (_19972_, _19971_, _19962_);
  and (_19973_, _11511_, _03859_);
  or (_19974_, _19973_, _19904_);
  and (_19975_, _19974_, _02331_);
  or (_19976_, _19975_, _19972_);
  and (_19978_, _19976_, _02208_);
  or (_19979_, _19904_, _04153_);
  and (_19980_, _19968_, _02206_);
  and (_19981_, _19980_, _19979_);
  or (_19982_, _19981_, _19978_);
  and (_19983_, _19982_, _03065_);
  and (_19984_, _19914_, _02342_);
  and (_19985_, _19984_, _19979_);
  or (_19986_, _19985_, _02202_);
  or (_19987_, _19986_, _19983_);
  nor (_19989_, _11503_, _08149_);
  or (_19990_, _19904_, _04953_);
  or (_19991_, _19990_, _19989_);
  and (_19992_, _19991_, _04958_);
  and (_19993_, _19992_, _19987_);
  nor (_19994_, _11510_, _08149_);
  or (_19995_, _19994_, _19904_);
  and (_19996_, _19995_, _02334_);
  or (_19997_, _19996_, _02366_);
  or (_19998_, _19997_, _19993_);
  or (_20000_, _19910_, _02778_);
  and (_20001_, _20000_, _01698_);
  and (_20002_, _20001_, _19998_);
  and (_20003_, _19935_, _01697_);
  or (_20004_, _20003_, _02081_);
  or (_20005_, _20004_, _20002_);
  and (_20006_, _11567_, _03859_);
  or (_20007_, _19904_, _02082_);
  or (_20008_, _20007_, _20006_);
  and (_20009_, _20008_, _39632_);
  and (_20011_, _20009_, _20005_);
  nor (_20012_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_20013_, _20012_, _00001_);
  or (_41679_, _20013_, _20011_);
  not (_20014_, \oc8051_golden_model_1.P1 [4]);
  nor (_20015_, _39632_, _20014_);
  or (_20016_, _20015_, rst);
  nor (_20017_, _03859_, _20014_);
  nor (_20018_, _04372_, _08149_);
  or (_20019_, _20018_, _20017_);
  or (_20021_, _20019_, _05444_);
  or (_20022_, _20019_, _02519_);
  nor (_20023_, _11611_, _08149_);
  or (_20024_, _20023_, _20017_);
  or (_20025_, _20024_, _03006_);
  and (_20026_, _03859_, \oc8051_golden_model_1.ACC [4]);
  or (_20027_, _20026_, _20017_);
  and (_20028_, _20027_, _02062_);
  nor (_20029_, _02062_, _20014_);
  or (_20030_, _20029_, _02158_);
  or (_20032_, _20030_, _20028_);
  and (_20033_, _20032_, _02058_);
  and (_20034_, _20033_, _20025_);
  nor (_20035_, _04489_, _20014_);
  and (_20036_, _11597_, _04489_);
  or (_20037_, _20036_, _20035_);
  and (_20038_, _20037_, _02057_);
  or (_20039_, _20038_, _02155_);
  or (_20040_, _20039_, _20034_);
  and (_20041_, _20040_, _20022_);
  or (_20043_, _20041_, _02153_);
  or (_20044_, _20027_, _02549_);
  and (_20045_, _20044_, _02054_);
  and (_20046_, _20045_, _20043_);
  and (_20047_, _11595_, _04489_);
  or (_20048_, _20047_, _20035_);
  and (_20049_, _20048_, _02053_);
  or (_20050_, _20049_, _02046_);
  or (_20051_, _20050_, _20046_);
  or (_20052_, _20035_, _11628_);
  and (_20054_, _20052_, _20037_);
  or (_20055_, _20054_, _02047_);
  and (_20056_, _20055_, _02043_);
  and (_20057_, _20056_, _20051_);
  and (_20058_, _19230_, _04489_);
  or (_20059_, _20058_, _20035_);
  and (_20060_, _20059_, _02042_);
  or (_20061_, _20060_, _06188_);
  or (_20062_, _20061_, _20057_);
  and (_20063_, _20062_, _20021_);
  or (_20065_, _20063_, _02031_);
  and (_20066_, _05303_, _03859_);
  or (_20067_, _20017_, _02032_);
  or (_20068_, _20067_, _20066_);
  and (_20069_, _20068_, _02037_);
  and (_20070_, _20069_, _20065_);
  and (_20071_, _19257_, _03859_);
  or (_20072_, _20017_, _20071_);
  and (_20073_, _20072_, _01765_);
  or (_20074_, _20073_, _20070_);
  or (_20076_, _20074_, _07629_);
  and (_20077_, _11592_, _03859_);
  or (_20078_, _20017_, _03059_);
  or (_20079_, _20078_, _20077_);
  and (_20080_, _04831_, _03859_);
  or (_20081_, _20080_, _20017_);
  or (_20082_, _20081_, _01995_);
  and (_20083_, _20082_, _03061_);
  and (_20084_, _20083_, _20079_);
  and (_20085_, _20084_, _20076_);
  and (_20087_, _11588_, _03859_);
  or (_20088_, _20087_, _20017_);
  and (_20089_, _20088_, _02331_);
  or (_20090_, _20089_, _20085_);
  and (_20091_, _20090_, _02208_);
  or (_20092_, _20017_, _04420_);
  and (_20093_, _20081_, _02206_);
  and (_20094_, _20093_, _20092_);
  or (_20095_, _20094_, _20091_);
  and (_20096_, _20095_, _03065_);
  and (_20098_, _20027_, _02342_);
  and (_20099_, _20098_, _20092_);
  or (_20100_, _20099_, _02202_);
  or (_20101_, _20100_, _20096_);
  nor (_20102_, _11590_, _08149_);
  or (_20103_, _20017_, _04953_);
  or (_20104_, _20103_, _20102_);
  and (_20105_, _20104_, _04958_);
  and (_20106_, _20105_, _20101_);
  nor (_20107_, _11587_, _08149_);
  or (_20109_, _20107_, _20017_);
  and (_20110_, _20109_, _02334_);
  or (_20111_, _20110_, _02366_);
  or (_20112_, _20111_, _20106_);
  or (_20113_, _20024_, _02778_);
  and (_20114_, _20113_, _01698_);
  and (_20115_, _20114_, _20112_);
  and (_20116_, _20048_, _01697_);
  or (_20117_, _20116_, _02081_);
  or (_20118_, _20117_, _20115_);
  and (_20120_, _11771_, _03859_);
  or (_20121_, _20017_, _02082_);
  or (_20122_, _20121_, _20120_);
  and (_20123_, _20122_, _39632_);
  and (_20124_, _20123_, _20118_);
  or (_41680_, _20124_, _20016_);
  not (_20125_, \oc8051_golden_model_1.P1 [5]);
  nor (_20126_, _03859_, _20125_);
  nor (_20127_, _04057_, _08149_);
  or (_20128_, _20127_, _20126_);
  or (_20130_, _20128_, _05444_);
  or (_20131_, _20128_, _02519_);
  nor (_20132_, _11804_, _08149_);
  or (_20133_, _20132_, _20126_);
  or (_20134_, _20133_, _03006_);
  and (_20135_, _03859_, \oc8051_golden_model_1.ACC [5]);
  or (_20136_, _20135_, _20126_);
  and (_20137_, _20136_, _02062_);
  nor (_20138_, _02062_, _20125_);
  or (_20139_, _20138_, _02158_);
  or (_20141_, _20139_, _20137_);
  and (_20142_, _20141_, _02058_);
  and (_20143_, _20142_, _20134_);
  nor (_20144_, _04489_, _20125_);
  and (_20145_, _11789_, _04489_);
  or (_20146_, _20145_, _20144_);
  and (_20147_, _20146_, _02057_);
  or (_20148_, _20147_, _02155_);
  or (_20149_, _20148_, _20143_);
  and (_20150_, _20149_, _20131_);
  or (_20152_, _20150_, _02153_);
  or (_20153_, _20136_, _02549_);
  and (_20154_, _20153_, _02054_);
  and (_20155_, _20154_, _20152_);
  and (_20156_, _11816_, _04489_);
  or (_20157_, _20156_, _20144_);
  and (_20158_, _20157_, _02053_);
  or (_20159_, _20158_, _02046_);
  or (_20160_, _20159_, _20155_);
  or (_20161_, _20144_, _11823_);
  and (_20163_, _20161_, _20146_);
  or (_20164_, _20163_, _02047_);
  and (_20165_, _20164_, _02043_);
  and (_20166_, _20165_, _20160_);
  and (_20167_, _19358_, _04489_);
  or (_20168_, _20167_, _20144_);
  and (_20169_, _20168_, _02042_);
  or (_20170_, _20169_, _06188_);
  or (_20171_, _20170_, _20166_);
  and (_20172_, _20171_, _20130_);
  or (_20174_, _20172_, _02031_);
  and (_20175_, _05258_, _03859_);
  or (_20176_, _20126_, _02032_);
  or (_20177_, _20176_, _20175_);
  and (_20178_, _20177_, _02037_);
  and (_20179_, _20178_, _20174_);
  and (_20180_, _19394_, _03859_);
  or (_20181_, _20180_, _20126_);
  and (_20182_, _20181_, _01765_);
  or (_20183_, _20182_, _20179_);
  or (_20185_, _20183_, _07629_);
  and (_20186_, _11915_, _03859_);
  or (_20187_, _20126_, _03059_);
  or (_20188_, _20187_, _20186_);
  and (_20189_, _04827_, _03859_);
  or (_20190_, _20189_, _20126_);
  or (_20191_, _20190_, _01995_);
  and (_20192_, _20191_, _03061_);
  and (_20193_, _20192_, _20188_);
  and (_20194_, _20193_, _20185_);
  and (_20196_, _11786_, _03859_);
  or (_20197_, _20196_, _20126_);
  and (_20198_, _20197_, _02331_);
  or (_20199_, _20198_, _20194_);
  and (_20200_, _20199_, _02208_);
  or (_20201_, _20126_, _04104_);
  and (_20202_, _20190_, _02206_);
  and (_20203_, _20202_, _20201_);
  or (_20204_, _20203_, _20200_);
  and (_20205_, _20204_, _03065_);
  and (_20207_, _20136_, _02342_);
  and (_20208_, _20207_, _20201_);
  or (_20209_, _20208_, _02202_);
  or (_20210_, _20209_, _20205_);
  nor (_20211_, _11913_, _08149_);
  or (_20212_, _20126_, _04953_);
  or (_20213_, _20212_, _20211_);
  and (_20214_, _20213_, _04958_);
  and (_20215_, _20214_, _20210_);
  nor (_20216_, _11785_, _08149_);
  or (_20218_, _20216_, _20126_);
  and (_20219_, _20218_, _02334_);
  or (_20220_, _20219_, _02366_);
  or (_20221_, _20220_, _20215_);
  or (_20222_, _20133_, _02778_);
  and (_20223_, _20222_, _01698_);
  and (_20224_, _20223_, _20221_);
  and (_20225_, _20157_, _01697_);
  or (_20226_, _20225_, _02081_);
  or (_20227_, _20226_, _20224_);
  and (_20229_, _11974_, _03859_);
  or (_20230_, _20126_, _02082_);
  or (_20231_, _20230_, _20229_);
  and (_20232_, _20231_, _39632_);
  and (_20233_, _20232_, _20227_);
  nor (_20234_, _39632_, _20125_);
  or (_20235_, _20234_, rst);
  or (_41681_, _20235_, _20233_);
  not (_20236_, \oc8051_golden_model_1.P1 [6]);
  nor (_20237_, _39632_, _20236_);
  or (_20239_, _20237_, rst);
  nor (_20240_, _03859_, _20236_);
  nor (_20241_, _03964_, _08149_);
  or (_20242_, _20241_, _20240_);
  or (_20243_, _20242_, _05444_);
  or (_20244_, _20242_, _02519_);
  nor (_20245_, _11993_, _08149_);
  or (_20246_, _20245_, _20240_);
  or (_20247_, _20246_, _03006_);
  and (_20248_, _03859_, \oc8051_golden_model_1.ACC [6]);
  or (_20250_, _20248_, _20240_);
  and (_20251_, _20250_, _02062_);
  nor (_20252_, _02062_, _20236_);
  or (_20253_, _20252_, _02158_);
  or (_20254_, _20253_, _20251_);
  and (_20255_, _20254_, _02058_);
  and (_20256_, _20255_, _20247_);
  nor (_20257_, _04489_, _20236_);
  and (_20258_, _11990_, _04489_);
  or (_20259_, _20258_, _20257_);
  and (_20261_, _20259_, _02057_);
  or (_20262_, _20261_, _02155_);
  or (_20263_, _20262_, _20256_);
  and (_20264_, _20263_, _20244_);
  or (_20265_, _20264_, _02153_);
  or (_20266_, _20250_, _02549_);
  and (_20267_, _20266_, _02054_);
  and (_20268_, _20267_, _20265_);
  and (_20269_, _12017_, _04489_);
  or (_20270_, _20269_, _20257_);
  and (_20272_, _20270_, _02053_);
  or (_20273_, _20272_, _02046_);
  or (_20274_, _20273_, _20268_);
  or (_20275_, _20257_, _12024_);
  and (_20276_, _20275_, _20259_);
  or (_20277_, _20276_, _02047_);
  and (_20278_, _20277_, _02043_);
  and (_20279_, _20278_, _20274_);
  and (_20280_, _19493_, _04489_);
  or (_20281_, _20280_, _20257_);
  and (_20283_, _20281_, _02042_);
  or (_20284_, _20283_, _06188_);
  or (_20285_, _20284_, _20279_);
  and (_20286_, _20285_, _20243_);
  or (_20287_, _20286_, _02031_);
  and (_20288_, _05029_, _03859_);
  or (_20289_, _20240_, _02032_);
  or (_20290_, _20289_, _20288_);
  and (_20291_, _20290_, _02037_);
  and (_20292_, _20291_, _20287_);
  and (_20294_, _19520_, _03859_);
  or (_20295_, _20294_, _20240_);
  and (_20296_, _20295_, _01765_);
  or (_20297_, _20296_, _20292_);
  or (_20298_, _20297_, _07629_);
  and (_20299_, _12112_, _03859_);
  or (_20300_, _20240_, _03059_);
  or (_20301_, _20300_, _20299_);
  and (_20302_, _12103_, _03859_);
  or (_20303_, _20302_, _20240_);
  or (_20305_, _20303_, _01995_);
  and (_20306_, _20305_, _03061_);
  and (_20307_, _20306_, _20301_);
  and (_20308_, _20307_, _20298_);
  and (_20309_, _12118_, _03859_);
  or (_20310_, _20309_, _20240_);
  and (_20311_, _20310_, _02331_);
  or (_20312_, _20311_, _20308_);
  and (_20313_, _20312_, _02208_);
  or (_20314_, _20240_, _04011_);
  and (_20316_, _20303_, _02206_);
  and (_20317_, _20316_, _20314_);
  or (_20318_, _20317_, _20313_);
  and (_20319_, _20318_, _03065_);
  and (_20320_, _20250_, _02342_);
  and (_20321_, _20320_, _20314_);
  or (_20322_, _20321_, _02202_);
  or (_20323_, _20322_, _20319_);
  nor (_20324_, _12110_, _08149_);
  or (_20325_, _20240_, _04953_);
  or (_20327_, _20325_, _20324_);
  and (_20328_, _20327_, _04958_);
  and (_20329_, _20328_, _20323_);
  nor (_20330_, _12117_, _08149_);
  or (_20331_, _20330_, _20240_);
  and (_20332_, _20331_, _02334_);
  or (_20333_, _20332_, _02366_);
  or (_20334_, _20333_, _20329_);
  or (_20335_, _20246_, _02778_);
  and (_20336_, _20335_, _01698_);
  and (_20338_, _20336_, _20334_);
  and (_20339_, _20270_, _01697_);
  or (_20340_, _20339_, _02081_);
  or (_20341_, _20340_, _20338_);
  and (_20342_, _12178_, _03859_);
  or (_20343_, _20240_, _02082_);
  or (_20344_, _20343_, _20342_);
  and (_20345_, _20344_, _39632_);
  and (_20346_, _20345_, _20341_);
  or (_41682_, _20346_, _20239_);
  not (_20348_, \oc8051_golden_model_1.P2 [0]);
  nor (_20349_, _03830_, _20348_);
  and (_20350_, _10792_, _03830_);
  or (_20351_, _20350_, _20349_);
  and (_20352_, _20351_, _02331_);
  and (_20353_, _03830_, _03002_);
  or (_20354_, _20353_, _20349_);
  or (_20355_, _20354_, _05444_);
  nor (_20356_, _04257_, _08250_);
  or (_20357_, _20356_, _20349_);
  and (_20359_, _20357_, _02158_);
  nor (_20360_, _02062_, _20348_);
  and (_20361_, _03830_, \oc8051_golden_model_1.ACC [0]);
  or (_20362_, _20361_, _20349_);
  and (_20363_, _20362_, _02062_);
  or (_20364_, _20363_, _20360_);
  and (_20365_, _20364_, _03006_);
  or (_20366_, _20365_, _02057_);
  or (_20367_, _20366_, _20359_);
  and (_20368_, _10814_, _04492_);
  nor (_20370_, _04492_, _20348_);
  or (_20371_, _20370_, _02058_);
  or (_20372_, _20371_, _20368_);
  and (_20373_, _20372_, _02519_);
  and (_20374_, _20373_, _20367_);
  and (_20375_, _20354_, _02155_);
  or (_20376_, _20375_, _02153_);
  or (_20377_, _20376_, _20374_);
  or (_20378_, _20362_, _02549_);
  and (_20379_, _20378_, _02054_);
  and (_20381_, _20379_, _20377_);
  and (_20382_, _20349_, _02053_);
  or (_20383_, _20382_, _02046_);
  or (_20384_, _20383_, _20381_);
  or (_20385_, _20357_, _02047_);
  and (_20386_, _20385_, _02043_);
  and (_20387_, _20386_, _20384_);
  and (_20388_, _18739_, _04492_);
  or (_20389_, _20388_, _20370_);
  and (_20390_, _20389_, _02042_);
  or (_20392_, _20390_, _06188_);
  or (_20393_, _20392_, _20387_);
  and (_20394_, _20393_, _20355_);
  or (_20395_, _20394_, _02031_);
  and (_20396_, _05120_, _03830_);
  or (_20397_, _20349_, _02032_);
  or (_20398_, _20397_, _20396_);
  and (_20399_, _20398_, _02037_);
  and (_20400_, _20399_, _20395_);
  and (_20401_, _18766_, _03830_);
  or (_20403_, _20401_, _20349_);
  and (_20404_, _20403_, _01765_);
  or (_20405_, _20404_, _20400_);
  or (_20406_, _20405_, _07629_);
  and (_20407_, _10914_, _03830_);
  or (_20408_, _20349_, _03059_);
  or (_20409_, _20408_, _20407_);
  and (_20410_, _03830_, _04837_);
  or (_20411_, _20410_, _20349_);
  or (_20412_, _20411_, _01995_);
  and (_20414_, _20412_, _03061_);
  and (_20415_, _20414_, _20409_);
  and (_20416_, _20415_, _20406_);
  or (_20417_, _20416_, _20352_);
  and (_20418_, _20417_, _02208_);
  nand (_20419_, _20411_, _02206_);
  nor (_20420_, _20419_, _20356_);
  or (_20421_, _20420_, _20418_);
  and (_20422_, _20421_, _03065_);
  or (_20423_, _20349_, _04257_);
  and (_20425_, _20362_, _02342_);
  and (_20426_, _20425_, _20423_);
  or (_20427_, _20426_, _02202_);
  or (_20428_, _20427_, _20422_);
  nor (_20429_, _10913_, _08250_);
  or (_20430_, _20349_, _04953_);
  or (_20431_, _20430_, _20429_);
  and (_20432_, _20431_, _04958_);
  and (_20433_, _20432_, _20428_);
  nor (_20434_, _10789_, _08250_);
  or (_20436_, _20434_, _20349_);
  and (_20437_, _20436_, _02334_);
  or (_20438_, _20437_, _02366_);
  or (_20439_, _20438_, _20433_);
  or (_20440_, _20357_, _02778_);
  and (_20441_, _20440_, _01698_);
  and (_20442_, _20441_, _20439_);
  and (_20443_, _20349_, _01697_);
  or (_20444_, _20443_, _02081_);
  or (_20445_, _20444_, _20442_);
  or (_20447_, _20357_, _02082_);
  and (_20448_, _20447_, _39632_);
  and (_20449_, _20448_, _20445_);
  nor (_20450_, _39632_, _20348_);
  or (_20451_, _20450_, rst);
  or (_41684_, _20451_, _20449_);
  not (_20452_, \oc8051_golden_model_1.P2 [1]);
  nor (_20453_, _03830_, _20452_);
  nor (_20454_, _08250_, _03161_);
  or (_20455_, _20454_, _20453_);
  or (_20457_, _20455_, _02519_);
  or (_20458_, _03830_, \oc8051_golden_model_1.P2 [1]);
  and (_20459_, _11001_, _03830_);
  not (_20460_, _20459_);
  and (_20461_, _20460_, _20458_);
  or (_20462_, _20461_, _03006_);
  nand (_20463_, _03830_, _01804_);
  and (_20464_, _20463_, _20458_);
  and (_20465_, _20464_, _02062_);
  nor (_20466_, _02062_, _20452_);
  or (_20468_, _20466_, _02158_);
  or (_20469_, _20468_, _20465_);
  and (_20470_, _20469_, _02058_);
  and (_20471_, _20470_, _20462_);
  nor (_20472_, _04492_, _20452_);
  and (_20473_, _11005_, _04492_);
  or (_20474_, _20473_, _20472_);
  and (_20475_, _20474_, _02057_);
  or (_20476_, _20475_, _02155_);
  or (_20477_, _20476_, _20471_);
  and (_20479_, _20477_, _20457_);
  or (_20480_, _20479_, _02153_);
  or (_20481_, _20464_, _02549_);
  and (_20482_, _20481_, _02054_);
  and (_20483_, _20482_, _20480_);
  and (_20484_, _10992_, _04492_);
  or (_20485_, _20484_, _20472_);
  and (_20486_, _20485_, _02053_);
  or (_20487_, _20486_, _20483_);
  or (_20488_, _20487_, _02046_);
  or (_20490_, _20472_, _11020_);
  and (_20491_, _20490_, _20474_);
  or (_20492_, _20491_, _02047_);
  and (_20493_, _20492_, _02043_);
  and (_20494_, _20493_, _20488_);
  and (_20495_, _18858_, _04492_);
  or (_20496_, _20495_, _20472_);
  and (_20497_, _20496_, _02042_);
  or (_20498_, _20497_, _06188_);
  or (_20499_, _20498_, _20494_);
  or (_20501_, _20455_, _05444_);
  and (_20502_, _20501_, _20499_);
  or (_20503_, _20502_, _02031_);
  and (_20504_, _05075_, _03830_);
  or (_20505_, _20453_, _02032_);
  or (_20506_, _20505_, _20504_);
  and (_20507_, _20506_, _02037_);
  and (_20508_, _20507_, _20503_);
  and (_20509_, _18887_, _03830_);
  or (_20510_, _20509_, _20453_);
  and (_20512_, _20510_, _01765_);
  or (_20513_, _20512_, _20508_);
  and (_20514_, _20513_, _02212_);
  or (_20515_, _10989_, _08250_);
  and (_20516_, _20515_, _02210_);
  nand (_20517_, _03830_, _02893_);
  and (_20518_, _20517_, _01994_);
  or (_20519_, _20518_, _20516_);
  and (_20520_, _20519_, _20458_);
  or (_20521_, _20520_, _20514_);
  and (_20523_, _20521_, _03061_);
  or (_20524_, _11113_, _08250_);
  and (_20525_, _20458_, _02331_);
  and (_20526_, _20525_, _20524_);
  or (_20527_, _20526_, _20523_);
  and (_20528_, _20527_, _02208_);
  or (_20529_, _10988_, _08250_);
  and (_20530_, _20458_, _02206_);
  and (_20531_, _20530_, _20529_);
  or (_20532_, _20531_, _20528_);
  and (_20534_, _20532_, _03065_);
  or (_20535_, _20453_, _04209_);
  and (_20536_, _20464_, _02342_);
  and (_20537_, _20536_, _20535_);
  or (_20538_, _20537_, _20534_);
  and (_20539_, _20538_, _02335_);
  or (_20540_, _20463_, _04209_);
  and (_20541_, _20458_, _02334_);
  and (_20542_, _20541_, _20540_);
  or (_20543_, _20542_, _02366_);
  or (_20545_, _20517_, _04209_);
  and (_20546_, _20458_, _02202_);
  and (_20547_, _20546_, _20545_);
  or (_20548_, _20547_, _20543_);
  or (_20549_, _20548_, _20539_);
  or (_20550_, _20461_, _02778_);
  and (_20551_, _20550_, _01698_);
  and (_20552_, _20551_, _20549_);
  and (_20553_, _20485_, _01697_);
  or (_20554_, _20553_, _02081_);
  or (_20556_, _20554_, _20552_);
  or (_20557_, _20453_, _02082_);
  or (_20558_, _20557_, _20459_);
  and (_20559_, _20558_, _39632_);
  and (_20560_, _20559_, _20556_);
  nor (_20561_, _39632_, _20452_);
  or (_20562_, _20561_, rst);
  or (_41685_, _20562_, _20560_);
  not (_20563_, \oc8051_golden_model_1.P2 [2]);
  nor (_20564_, _03830_, _20563_);
  nor (_20566_, _08250_, _03624_);
  or (_20567_, _20566_, _20564_);
  or (_20568_, _20567_, _05444_);
  nor (_20569_, _11199_, _08250_);
  or (_20570_, _20569_, _20564_);
  and (_20571_, _20570_, _02158_);
  nor (_20572_, _02062_, _20563_);
  and (_20573_, _03830_, \oc8051_golden_model_1.ACC [2]);
  or (_20574_, _20573_, _20564_);
  and (_20575_, _20574_, _02062_);
  or (_20577_, _20575_, _20572_);
  and (_20578_, _20577_, _03006_);
  or (_20579_, _20578_, _02057_);
  or (_20580_, _20579_, _20571_);
  nor (_20581_, _04492_, _20563_);
  and (_20582_, _11194_, _04492_);
  or (_20583_, _20582_, _20581_);
  or (_20584_, _20583_, _02058_);
  and (_20585_, _20584_, _20580_);
  or (_20586_, _20585_, _02155_);
  or (_20588_, _20567_, _02519_);
  and (_20589_, _20588_, _20586_);
  or (_20590_, _20589_, _02153_);
  or (_20591_, _20574_, _02549_);
  and (_20592_, _20591_, _02054_);
  and (_20593_, _20592_, _20590_);
  and (_20594_, _11192_, _04492_);
  or (_20595_, _20594_, _20581_);
  and (_20596_, _20595_, _02053_);
  or (_20597_, _20596_, _02046_);
  or (_20599_, _20597_, _20593_);
  or (_20600_, _20581_, _11223_);
  and (_20601_, _20600_, _20583_);
  or (_20602_, _20601_, _02047_);
  and (_20603_, _20602_, _02043_);
  and (_20604_, _20603_, _20599_);
  and (_20605_, _18983_, _04492_);
  or (_20606_, _20605_, _20581_);
  and (_20607_, _20606_, _02042_);
  or (_20608_, _20607_, _06188_);
  or (_20610_, _20608_, _20604_);
  and (_20611_, _20610_, _20568_);
  or (_20612_, _20611_, _02031_);
  and (_20613_, _05211_, _03830_);
  or (_20614_, _20564_, _02032_);
  or (_20615_, _20614_, _20613_);
  and (_20616_, _20615_, _02037_);
  and (_20617_, _20616_, _20612_);
  and (_20618_, _19008_, _03830_);
  or (_20619_, _20564_, _20618_);
  and (_20621_, _20619_, _01765_);
  or (_20622_, _20621_, _20617_);
  or (_20623_, _20622_, _07629_);
  and (_20624_, _11189_, _03830_);
  or (_20625_, _20564_, _03059_);
  or (_20626_, _20625_, _20624_);
  and (_20627_, _03830_, _04866_);
  or (_20628_, _20627_, _20564_);
  or (_20629_, _20628_, _01995_);
  and (_20630_, _20629_, _03061_);
  and (_20632_, _20630_, _20626_);
  and (_20633_, _20632_, _20623_);
  and (_20634_, _11315_, _03830_);
  or (_20635_, _20634_, _20564_);
  and (_20636_, _20635_, _02331_);
  or (_20637_, _20636_, _20633_);
  and (_20638_, _20637_, _02208_);
  or (_20639_, _20564_, _04309_);
  and (_20640_, _20628_, _02206_);
  and (_20641_, _20640_, _20639_);
  or (_20643_, _20641_, _20638_);
  and (_20644_, _20643_, _03065_);
  and (_20645_, _20574_, _02342_);
  and (_20646_, _20645_, _20639_);
  or (_20647_, _20646_, _02202_);
  or (_20648_, _20647_, _20644_);
  nor (_20649_, _11187_, _08250_);
  or (_20650_, _20564_, _04953_);
  or (_20651_, _20650_, _20649_);
  and (_20652_, _20651_, _04958_);
  and (_20654_, _20652_, _20648_);
  nor (_20655_, _11314_, _08250_);
  or (_20656_, _20655_, _20564_);
  and (_20657_, _20656_, _02334_);
  or (_20658_, _20657_, _02366_);
  or (_20659_, _20658_, _20654_);
  or (_20660_, _20570_, _02778_);
  and (_20661_, _20660_, _01698_);
  and (_20662_, _20661_, _20659_);
  and (_20663_, _20595_, _01697_);
  or (_20665_, _20663_, _02081_);
  or (_20666_, _20665_, _20662_);
  and (_20667_, _11367_, _03830_);
  or (_20668_, _20564_, _02082_);
  or (_20669_, _20668_, _20667_);
  and (_20670_, _20669_, _39632_);
  and (_20671_, _20670_, _20666_);
  nor (_20672_, _39632_, _20563_);
  or (_20673_, _20672_, rst);
  or (_41686_, _20673_, _20671_);
  not (_20675_, \oc8051_golden_model_1.P2 [3]);
  nor (_20676_, _39632_, _20675_);
  or (_20677_, _20676_, rst);
  nor (_20678_, _03830_, _20675_);
  nor (_20679_, _08250_, _03434_);
  or (_20680_, _20679_, _20678_);
  or (_20681_, _20680_, _05444_);
  or (_20682_, _20680_, _02519_);
  nor (_20683_, _11394_, _08250_);
  or (_20684_, _20683_, _20678_);
  or (_20686_, _20684_, _03006_);
  and (_20687_, _03830_, \oc8051_golden_model_1.ACC [3]);
  or (_20688_, _20687_, _20678_);
  and (_20689_, _20688_, _02062_);
  nor (_20690_, _02062_, _20675_);
  or (_20691_, _20690_, _02158_);
  or (_20692_, _20691_, _20689_);
  and (_20693_, _20692_, _02058_);
  and (_20694_, _20693_, _20686_);
  nor (_20695_, _04492_, _20675_);
  and (_20697_, _11398_, _04492_);
  or (_20698_, _20697_, _20695_);
  and (_20699_, _20698_, _02057_);
  or (_20700_, _20699_, _02155_);
  or (_20701_, _20700_, _20694_);
  and (_20702_, _20701_, _20682_);
  or (_20703_, _20702_, _02153_);
  or (_20704_, _20688_, _02549_);
  and (_20705_, _20704_, _02054_);
  and (_20706_, _20705_, _20703_);
  and (_20708_, _11408_, _04492_);
  or (_20709_, _20708_, _20695_);
  and (_20710_, _20709_, _02053_);
  or (_20711_, _20710_, _02046_);
  or (_20712_, _20711_, _20706_);
  or (_20713_, _20695_, _11415_);
  and (_20714_, _20713_, _20698_);
  or (_20715_, _20714_, _02047_);
  and (_20716_, _20715_, _02043_);
  and (_20717_, _20716_, _20712_);
  and (_20719_, _19106_, _04492_);
  or (_20720_, _20719_, _20695_);
  and (_20721_, _20720_, _02042_);
  or (_20722_, _20721_, _06188_);
  or (_20723_, _20722_, _20717_);
  and (_20724_, _20723_, _20681_);
  or (_20725_, _20724_, _02031_);
  and (_20726_, _05166_, _03830_);
  or (_20727_, _20678_, _02032_);
  or (_20728_, _20727_, _20726_);
  and (_20730_, _20728_, _02037_);
  and (_20731_, _20730_, _20725_);
  and (_20732_, _19131_, _03830_);
  or (_20733_, _20678_, _20732_);
  and (_20734_, _20733_, _01765_);
  or (_20735_, _20734_, _20731_);
  or (_20736_, _20735_, _07629_);
  and (_20737_, _11505_, _03830_);
  or (_20738_, _20678_, _03059_);
  or (_20739_, _20738_, _20737_);
  and (_20741_, _03830_, _04719_);
  or (_20742_, _20741_, _20678_);
  or (_20743_, _20742_, _01995_);
  and (_20744_, _20743_, _03061_);
  and (_20745_, _20744_, _20739_);
  and (_20746_, _20745_, _20736_);
  and (_20747_, _11511_, _03830_);
  or (_20748_, _20747_, _20678_);
  and (_20749_, _20748_, _02331_);
  or (_20750_, _20749_, _20746_);
  and (_20752_, _20750_, _02208_);
  or (_20753_, _20678_, _04153_);
  and (_20754_, _20742_, _02206_);
  and (_20755_, _20754_, _20753_);
  or (_20756_, _20755_, _20752_);
  and (_20757_, _20756_, _03065_);
  and (_20758_, _20688_, _02342_);
  and (_20759_, _20758_, _20753_);
  or (_20760_, _20759_, _02202_);
  or (_20761_, _20760_, _20757_);
  nor (_20763_, _11503_, _08250_);
  or (_20764_, _20678_, _04953_);
  or (_20765_, _20764_, _20763_);
  and (_20766_, _20765_, _04958_);
  and (_20767_, _20766_, _20761_);
  nor (_20768_, _11510_, _08250_);
  or (_20769_, _20768_, _20678_);
  and (_20770_, _20769_, _02334_);
  or (_20771_, _20770_, _02366_);
  or (_20772_, _20771_, _20767_);
  or (_20774_, _20684_, _02778_);
  and (_20775_, _20774_, _01698_);
  and (_20776_, _20775_, _20772_);
  and (_20777_, _20709_, _01697_);
  or (_20778_, _20777_, _02081_);
  or (_20779_, _20778_, _20776_);
  and (_20780_, _11567_, _03830_);
  or (_20781_, _20678_, _02082_);
  or (_20782_, _20781_, _20780_);
  and (_20783_, _20782_, _39632_);
  and (_20785_, _20783_, _20779_);
  or (_41687_, _20785_, _20677_);
  not (_20786_, \oc8051_golden_model_1.P2 [4]);
  nor (_20787_, _03830_, _20786_);
  nor (_20788_, _04372_, _08250_);
  or (_20789_, _20788_, _20787_);
  or (_20790_, _20789_, _05444_);
  or (_20791_, _20789_, _02519_);
  nor (_20792_, _11611_, _08250_);
  or (_20793_, _20792_, _20787_);
  or (_20795_, _20793_, _03006_);
  and (_20796_, _03830_, \oc8051_golden_model_1.ACC [4]);
  or (_20797_, _20796_, _20787_);
  and (_20798_, _20797_, _02062_);
  nor (_20799_, _02062_, _20786_);
  or (_20800_, _20799_, _02158_);
  or (_20801_, _20800_, _20798_);
  and (_20802_, _20801_, _02058_);
  and (_20803_, _20802_, _20795_);
  nor (_20804_, _04492_, _20786_);
  and (_20806_, _11597_, _04492_);
  or (_20807_, _20806_, _20804_);
  and (_20808_, _20807_, _02057_);
  or (_20809_, _20808_, _02155_);
  or (_20810_, _20809_, _20803_);
  and (_20811_, _20810_, _20791_);
  or (_20812_, _20811_, _02153_);
  or (_20813_, _20797_, _02549_);
  and (_20814_, _20813_, _02054_);
  and (_20815_, _20814_, _20812_);
  and (_20817_, _11595_, _04492_);
  or (_20818_, _20817_, _20804_);
  and (_20819_, _20818_, _02053_);
  or (_20820_, _20819_, _02046_);
  or (_20821_, _20820_, _20815_);
  or (_20822_, _20804_, _11628_);
  and (_20823_, _20822_, _20807_);
  or (_20824_, _20823_, _02047_);
  and (_20825_, _20824_, _02043_);
  and (_20826_, _20825_, _20821_);
  and (_20828_, _19230_, _04492_);
  or (_20829_, _20828_, _20804_);
  and (_20830_, _20829_, _02042_);
  or (_20831_, _20830_, _06188_);
  or (_20832_, _20831_, _20826_);
  and (_20833_, _20832_, _20790_);
  or (_20834_, _20833_, _02031_);
  and (_20835_, _05303_, _03830_);
  or (_20836_, _20787_, _02032_);
  or (_20837_, _20836_, _20835_);
  and (_20839_, _20837_, _02037_);
  and (_20840_, _20839_, _20834_);
  and (_20841_, _19257_, _03830_);
  or (_20842_, _20787_, _20841_);
  and (_20843_, _20842_, _01765_);
  or (_20844_, _20843_, _20840_);
  or (_20845_, _20844_, _07629_);
  and (_20846_, _11592_, _03830_);
  or (_20847_, _20787_, _03059_);
  or (_20848_, _20847_, _20846_);
  and (_20850_, _04831_, _03830_);
  or (_20851_, _20850_, _20787_);
  or (_20852_, _20851_, _01995_);
  and (_20853_, _20852_, _03061_);
  and (_20854_, _20853_, _20848_);
  and (_20855_, _20854_, _20845_);
  and (_20856_, _11588_, _03830_);
  or (_20857_, _20856_, _20787_);
  and (_20858_, _20857_, _02331_);
  or (_20859_, _20858_, _20855_);
  and (_20861_, _20859_, _02208_);
  or (_20862_, _20787_, _04420_);
  and (_20863_, _20851_, _02206_);
  and (_20864_, _20863_, _20862_);
  or (_20865_, _20864_, _20861_);
  and (_20866_, _20865_, _03065_);
  and (_20867_, _20797_, _02342_);
  and (_20868_, _20867_, _20862_);
  or (_20869_, _20868_, _02202_);
  or (_20870_, _20869_, _20866_);
  nor (_20872_, _11590_, _08250_);
  or (_20873_, _20787_, _04953_);
  or (_20874_, _20873_, _20872_);
  and (_20875_, _20874_, _04958_);
  and (_20876_, _20875_, _20870_);
  nor (_20877_, _11587_, _08250_);
  or (_20878_, _20877_, _20787_);
  and (_20879_, _20878_, _02334_);
  or (_20880_, _20879_, _02366_);
  or (_20881_, _20880_, _20876_);
  or (_20883_, _20793_, _02778_);
  and (_20884_, _20883_, _01698_);
  and (_20885_, _20884_, _20881_);
  and (_20886_, _20818_, _01697_);
  or (_20887_, _20886_, _02081_);
  or (_20888_, _20887_, _20885_);
  and (_20889_, _11771_, _03830_);
  or (_20890_, _20787_, _02082_);
  or (_20891_, _20890_, _20889_);
  and (_20892_, _20891_, _39632_);
  and (_20894_, _20892_, _20888_);
  nor (_20895_, _39632_, _20786_);
  or (_20896_, _20895_, rst);
  or (_41688_, _20896_, _20894_);
  not (_20897_, \oc8051_golden_model_1.P2 [5]);
  nor (_20898_, _03830_, _20897_);
  nor (_20899_, _04057_, _08250_);
  or (_20900_, _20899_, _20898_);
  or (_20901_, _20900_, _05444_);
  or (_20902_, _20900_, _02519_);
  nor (_20904_, _11804_, _08250_);
  or (_20905_, _20904_, _20898_);
  or (_20906_, _20905_, _03006_);
  and (_20907_, _03830_, \oc8051_golden_model_1.ACC [5]);
  or (_20908_, _20907_, _20898_);
  and (_20909_, _20908_, _02062_);
  nor (_20910_, _02062_, _20897_);
  or (_20911_, _20910_, _02158_);
  or (_20912_, _20911_, _20909_);
  and (_20913_, _20912_, _02058_);
  and (_20915_, _20913_, _20906_);
  nor (_20916_, _04492_, _20897_);
  and (_20917_, _11789_, _04492_);
  or (_20918_, _20917_, _20916_);
  and (_20919_, _20918_, _02057_);
  or (_20920_, _20919_, _02155_);
  or (_20921_, _20920_, _20915_);
  and (_20922_, _20921_, _20902_);
  or (_20923_, _20922_, _02153_);
  or (_20924_, _20908_, _02549_);
  and (_20926_, _20924_, _02054_);
  and (_20927_, _20926_, _20923_);
  and (_20928_, _11816_, _04492_);
  or (_20929_, _20928_, _20916_);
  and (_20930_, _20929_, _02053_);
  or (_20931_, _20930_, _02046_);
  or (_20932_, _20931_, _20927_);
  or (_20933_, _20916_, _11823_);
  and (_20934_, _20933_, _20918_);
  or (_20935_, _20934_, _02047_);
  and (_20937_, _20935_, _02043_);
  and (_20938_, _20937_, _20932_);
  and (_20939_, _19358_, _04492_);
  or (_20940_, _20939_, _20916_);
  and (_20941_, _20940_, _02042_);
  or (_20942_, _20941_, _06188_);
  or (_20943_, _20942_, _20938_);
  and (_20944_, _20943_, _20901_);
  or (_20945_, _20944_, _02031_);
  and (_20946_, _05258_, _03830_);
  or (_20948_, _20898_, _02032_);
  or (_20949_, _20948_, _20946_);
  and (_20950_, _20949_, _02037_);
  and (_20951_, _20950_, _20945_);
  and (_20952_, _19394_, _03830_);
  or (_20953_, _20952_, _20898_);
  and (_20954_, _20953_, _01765_);
  or (_20955_, _20954_, _20951_);
  or (_20956_, _20955_, _07629_);
  and (_20957_, _11915_, _03830_);
  or (_20959_, _20898_, _03059_);
  or (_20960_, _20959_, _20957_);
  and (_20961_, _04827_, _03830_);
  or (_20962_, _20961_, _20898_);
  or (_20963_, _20962_, _01995_);
  and (_20964_, _20963_, _03061_);
  and (_20965_, _20964_, _20960_);
  and (_20966_, _20965_, _20956_);
  and (_20967_, _11786_, _03830_);
  or (_20968_, _20967_, _20898_);
  and (_20970_, _20968_, _02331_);
  or (_20971_, _20970_, _20966_);
  and (_20972_, _20971_, _02208_);
  or (_20973_, _20898_, _04104_);
  and (_20974_, _20962_, _02206_);
  and (_20975_, _20974_, _20973_);
  or (_20976_, _20975_, _20972_);
  and (_20977_, _20976_, _03065_);
  and (_20978_, _20908_, _02342_);
  and (_20979_, _20978_, _20973_);
  or (_20981_, _20979_, _02202_);
  or (_20982_, _20981_, _20977_);
  nor (_20983_, _11913_, _08250_);
  or (_20984_, _20898_, _04953_);
  or (_20985_, _20984_, _20983_);
  and (_20986_, _20985_, _04958_);
  and (_20987_, _20986_, _20982_);
  nor (_20988_, _11785_, _08250_);
  or (_20989_, _20988_, _20898_);
  and (_20990_, _20989_, _02334_);
  or (_20992_, _20990_, _02366_);
  or (_20993_, _20992_, _20987_);
  or (_20994_, _20905_, _02778_);
  and (_20995_, _20994_, _01698_);
  and (_20996_, _20995_, _20993_);
  and (_20997_, _20929_, _01697_);
  or (_20998_, _20997_, _02081_);
  or (_20999_, _20998_, _20996_);
  and (_21000_, _11974_, _03830_);
  or (_21001_, _20898_, _02082_);
  or (_21003_, _21001_, _21000_);
  and (_21004_, _21003_, _39632_);
  and (_21005_, _21004_, _20999_);
  nor (_21006_, _39632_, _20897_);
  or (_21007_, _21006_, rst);
  or (_41689_, _21007_, _21005_);
  not (_21008_, \oc8051_golden_model_1.P2 [6]);
  nor (_21009_, _03830_, _21008_);
  nor (_21010_, _03964_, _08250_);
  or (_21011_, _21010_, _21009_);
  or (_21013_, _21011_, _05444_);
  or (_21014_, _21011_, _02519_);
  nor (_21015_, _11993_, _08250_);
  or (_21016_, _21015_, _21009_);
  or (_21017_, _21016_, _03006_);
  and (_21018_, _03830_, \oc8051_golden_model_1.ACC [6]);
  or (_21019_, _21018_, _21009_);
  and (_21020_, _21019_, _02062_);
  nor (_21021_, _02062_, _21008_);
  or (_21022_, _21021_, _02158_);
  or (_21024_, _21022_, _21020_);
  and (_21025_, _21024_, _02058_);
  and (_21026_, _21025_, _21017_);
  nor (_21027_, _04492_, _21008_);
  and (_21028_, _11990_, _04492_);
  or (_21029_, _21028_, _21027_);
  and (_21030_, _21029_, _02057_);
  or (_21031_, _21030_, _02155_);
  or (_21032_, _21031_, _21026_);
  and (_21033_, _21032_, _21014_);
  or (_21035_, _21033_, _02153_);
  or (_21036_, _21019_, _02549_);
  and (_21037_, _21036_, _02054_);
  and (_21038_, _21037_, _21035_);
  and (_21039_, _12017_, _04492_);
  or (_21040_, _21039_, _21027_);
  and (_21041_, _21040_, _02053_);
  or (_21042_, _21041_, _02046_);
  or (_21043_, _21042_, _21038_);
  or (_21044_, _21027_, _12024_);
  and (_21046_, _21044_, _21029_);
  or (_21047_, _21046_, _02047_);
  and (_21048_, _21047_, _02043_);
  and (_21049_, _21048_, _21043_);
  and (_21050_, _19493_, _04492_);
  or (_21051_, _21050_, _21027_);
  and (_21052_, _21051_, _02042_);
  or (_21053_, _21052_, _06188_);
  or (_21054_, _21053_, _21049_);
  and (_21055_, _21054_, _21013_);
  or (_21057_, _21055_, _02031_);
  and (_21058_, _05029_, _03830_);
  or (_21059_, _21009_, _02032_);
  or (_21060_, _21059_, _21058_);
  and (_21061_, _21060_, _02037_);
  and (_21062_, _21061_, _21057_);
  and (_21063_, _19520_, _03830_);
  or (_21064_, _21063_, _21009_);
  and (_21065_, _21064_, _01765_);
  or (_21066_, _21065_, _21062_);
  or (_21068_, _21066_, _07629_);
  and (_21069_, _12112_, _03830_);
  or (_21070_, _21009_, _03059_);
  or (_21071_, _21070_, _21069_);
  and (_21072_, _12103_, _03830_);
  or (_21073_, _21072_, _21009_);
  or (_21074_, _21073_, _01995_);
  and (_21075_, _21074_, _03061_);
  and (_21076_, _21075_, _21071_);
  and (_21077_, _21076_, _21068_);
  and (_21079_, _12118_, _03830_);
  or (_21080_, _21079_, _21009_);
  and (_21081_, _21080_, _02331_);
  or (_21082_, _21081_, _21077_);
  and (_21083_, _21082_, _02208_);
  or (_21084_, _21009_, _04011_);
  and (_21085_, _21073_, _02206_);
  and (_21086_, _21085_, _21084_);
  or (_21087_, _21086_, _21083_);
  and (_21088_, _21087_, _03065_);
  and (_21090_, _21019_, _02342_);
  and (_21091_, _21090_, _21084_);
  or (_21092_, _21091_, _02202_);
  or (_21093_, _21092_, _21088_);
  nor (_21094_, _12110_, _08250_);
  or (_21095_, _21009_, _04953_);
  or (_21096_, _21095_, _21094_);
  and (_21097_, _21096_, _04958_);
  and (_21098_, _21097_, _21093_);
  nor (_21099_, _12117_, _08250_);
  or (_21101_, _21099_, _21009_);
  and (_21102_, _21101_, _02334_);
  or (_21103_, _21102_, _02366_);
  or (_21104_, _21103_, _21098_);
  or (_21105_, _21016_, _02778_);
  and (_21106_, _21105_, _01698_);
  and (_21107_, _21106_, _21104_);
  and (_21108_, _21040_, _01697_);
  or (_21109_, _21108_, _02081_);
  or (_21110_, _21109_, _21107_);
  and (_21112_, _12178_, _03830_);
  or (_21113_, _21009_, _02082_);
  or (_21114_, _21113_, _21112_);
  and (_21115_, _21114_, _39632_);
  and (_21116_, _21115_, _21110_);
  nor (_21117_, _39632_, _21008_);
  or (_21118_, _21117_, rst);
  or (_41690_, _21118_, _21116_);
  not (_21119_, \oc8051_golden_model_1.P3 [0]);
  nor (_21120_, _39632_, _21119_);
  or (_21122_, _21120_, rst);
  nor (_21123_, _04257_, _08358_);
  nor (_21124_, _03820_, _21119_);
  and (_21125_, _03820_, _04837_);
  or (_21126_, _21125_, _21124_);
  nand (_21127_, _21126_, _02206_);
  nor (_21128_, _21127_, _21123_);
  and (_21129_, _10792_, _03820_);
  or (_21130_, _21129_, _21124_);
  and (_21131_, _21130_, _02331_);
  and (_21133_, _03820_, _03002_);
  or (_21134_, _21133_, _21124_);
  or (_21135_, _21134_, _05444_);
  or (_21136_, _21124_, _21123_);
  or (_21137_, _21136_, _03006_);
  and (_21138_, _03820_, \oc8051_golden_model_1.ACC [0]);
  or (_21139_, _21138_, _21124_);
  and (_21140_, _21139_, _02062_);
  nor (_21141_, _02062_, _21119_);
  or (_21142_, _21141_, _02158_);
  or (_21144_, _21142_, _21140_);
  and (_21145_, _21144_, _02058_);
  and (_21146_, _21145_, _21137_);
  nor (_21147_, _04467_, _21119_);
  and (_21148_, _10814_, _04467_);
  or (_21149_, _21148_, _21147_);
  and (_21150_, _21149_, _02057_);
  or (_21151_, _21150_, _21146_);
  and (_21152_, _21151_, _02519_);
  and (_21153_, _21134_, _02155_);
  or (_21155_, _21153_, _02153_);
  or (_21156_, _21155_, _21152_);
  or (_21157_, _21139_, _02549_);
  and (_21158_, _21157_, _02054_);
  and (_21159_, _21158_, _21156_);
  and (_21160_, _21124_, _02053_);
  or (_21161_, _21160_, _02046_);
  or (_21162_, _21161_, _21159_);
  or (_21163_, _21136_, _02047_);
  and (_21164_, _21163_, _02043_);
  and (_21166_, _21164_, _21162_);
  and (_21167_, _18739_, _04467_);
  or (_21168_, _21167_, _21147_);
  and (_21169_, _21168_, _02042_);
  or (_21170_, _21169_, _06188_);
  or (_21171_, _21170_, _21166_);
  and (_21172_, _21171_, _21135_);
  or (_21173_, _21172_, _02031_);
  and (_21174_, _05120_, _03820_);
  or (_21175_, _21124_, _02032_);
  or (_21177_, _21175_, _21174_);
  and (_21178_, _21177_, _02037_);
  and (_21179_, _21178_, _21173_);
  and (_21180_, _18766_, _03820_);
  or (_21181_, _21180_, _21124_);
  and (_21182_, _21181_, _01765_);
  or (_21183_, _21182_, _21179_);
  or (_21184_, _21183_, _07629_);
  and (_21185_, _10914_, _03820_);
  or (_21186_, _21124_, _03059_);
  or (_21188_, _21186_, _21185_);
  or (_21189_, _21126_, _01995_);
  and (_21190_, _21189_, _03061_);
  and (_21191_, _21190_, _21188_);
  and (_21192_, _21191_, _21184_);
  or (_21193_, _21192_, _21131_);
  and (_21194_, _21193_, _02208_);
  or (_21195_, _21194_, _21128_);
  and (_21196_, _21195_, _03065_);
  or (_21197_, _21124_, _04257_);
  and (_21199_, _21139_, _02342_);
  and (_21200_, _21199_, _21197_);
  or (_21201_, _21200_, _02202_);
  or (_21202_, _21201_, _21196_);
  nor (_21203_, _10913_, _08358_);
  or (_21204_, _21124_, _04953_);
  or (_21205_, _21204_, _21203_);
  and (_21206_, _21205_, _04958_);
  and (_21207_, _21206_, _21202_);
  nor (_21208_, _10789_, _08358_);
  or (_21210_, _21208_, _21124_);
  and (_21211_, _21210_, _02334_);
  or (_21212_, _21211_, _02366_);
  or (_21213_, _21212_, _21207_);
  or (_21214_, _21136_, _02778_);
  and (_21215_, _21214_, _01698_);
  and (_21216_, _21215_, _21213_);
  and (_21217_, _21124_, _01697_);
  or (_21218_, _21217_, _02081_);
  or (_21219_, _21218_, _21216_);
  or (_21221_, _21136_, _02082_);
  and (_21222_, _21221_, _39632_);
  and (_21223_, _21222_, _21219_);
  or (_41692_, _21223_, _21122_);
  or (_21224_, _11113_, _08358_);
  or (_21225_, _03820_, \oc8051_golden_model_1.P3 [1]);
  and (_21226_, _21225_, _02331_);
  and (_21227_, _21226_, _21224_);
  not (_21228_, \oc8051_golden_model_1.P3 [1]);
  nor (_21229_, _03820_, _21228_);
  nor (_21231_, _08358_, _03161_);
  or (_21232_, _21231_, _21229_);
  or (_21233_, _21232_, _02519_);
  and (_21234_, _11001_, _03820_);
  not (_21235_, _21234_);
  and (_21236_, _21235_, _21225_);
  or (_21237_, _21236_, _03006_);
  nand (_21238_, _03820_, _01804_);
  and (_21239_, _21238_, _21225_);
  and (_21240_, _21239_, _02062_);
  nor (_21242_, _02062_, _21228_);
  or (_21243_, _21242_, _02158_);
  or (_21244_, _21243_, _21240_);
  and (_21245_, _21244_, _02058_);
  and (_21246_, _21245_, _21237_);
  nor (_21247_, _04467_, _21228_);
  and (_21248_, _11005_, _04467_);
  or (_21249_, _21248_, _21247_);
  and (_21250_, _21249_, _02057_);
  or (_21251_, _21250_, _02155_);
  or (_21253_, _21251_, _21246_);
  and (_21254_, _21253_, _21233_);
  or (_21255_, _21254_, _02153_);
  or (_21256_, _21239_, _02549_);
  and (_21257_, _21256_, _02054_);
  and (_21258_, _21257_, _21255_);
  and (_21259_, _10992_, _04467_);
  or (_21260_, _21259_, _21247_);
  and (_21261_, _21260_, _02053_);
  or (_21262_, _21261_, _02046_);
  or (_21264_, _21262_, _21258_);
  or (_21265_, _21247_, _11020_);
  and (_21266_, _21265_, _21249_);
  or (_21267_, _21266_, _02047_);
  and (_21268_, _21267_, _02043_);
  and (_21269_, _21268_, _21264_);
  and (_21270_, _18858_, _04467_);
  or (_21271_, _21270_, _21247_);
  and (_21272_, _21271_, _02042_);
  or (_21273_, _21272_, _06188_);
  or (_21275_, _21273_, _21269_);
  or (_21276_, _21232_, _05444_);
  and (_21277_, _21276_, _21275_);
  or (_21278_, _21277_, _02031_);
  and (_21279_, _05075_, _03820_);
  or (_21280_, _21229_, _02032_);
  or (_21281_, _21280_, _21279_);
  and (_21282_, _21281_, _02037_);
  and (_21283_, _21282_, _21278_);
  or (_21284_, _18887_, _08358_);
  and (_21286_, _21225_, _01765_);
  and (_21287_, _21286_, _21284_);
  or (_21288_, _21287_, _21283_);
  and (_21289_, _21288_, _02212_);
  or (_21290_, _10989_, _08358_);
  and (_21291_, _21290_, _02210_);
  nand (_21292_, _03820_, _02893_);
  and (_21293_, _21292_, _01994_);
  or (_21294_, _21293_, _21291_);
  and (_21295_, _21294_, _21225_);
  or (_21297_, _21295_, _21289_);
  and (_21298_, _21297_, _03061_);
  or (_21299_, _21298_, _21227_);
  and (_21300_, _21299_, _02208_);
  or (_21301_, _10988_, _08358_);
  and (_21302_, _21225_, _02206_);
  and (_21303_, _21302_, _21301_);
  or (_21304_, _21303_, _21300_);
  and (_21305_, _21304_, _03065_);
  or (_21306_, _21229_, _04209_);
  and (_21308_, _21239_, _02342_);
  and (_21309_, _21308_, _21306_);
  or (_21310_, _21309_, _21305_);
  and (_21311_, _21310_, _02335_);
  or (_21312_, _21238_, _04209_);
  and (_21313_, _21225_, _02334_);
  and (_21314_, _21313_, _21312_);
  or (_21315_, _21314_, _02366_);
  or (_21316_, _21292_, _04209_);
  and (_21317_, _21225_, _02202_);
  and (_21319_, _21317_, _21316_);
  or (_21320_, _21319_, _21315_);
  or (_21321_, _21320_, _21311_);
  or (_21322_, _21236_, _02778_);
  and (_21323_, _21322_, _01698_);
  and (_21324_, _21323_, _21321_);
  and (_21325_, _21260_, _01697_);
  or (_21326_, _21325_, _02081_);
  or (_21327_, _21326_, _21324_);
  or (_21328_, _21229_, _02082_);
  or (_21330_, _21328_, _21234_);
  and (_21331_, _21330_, _39632_);
  and (_21332_, _21331_, _21327_);
  nor (_21333_, _39632_, _21228_);
  or (_21334_, _21333_, rst);
  or (_41693_, _21334_, _21332_);
  not (_21335_, \oc8051_golden_model_1.P3 [2]);
  nor (_21336_, _03820_, _21335_);
  and (_21337_, _11315_, _03820_);
  or (_21338_, _21337_, _21336_);
  and (_21340_, _21338_, _02331_);
  nor (_21341_, _08358_, _03624_);
  or (_21342_, _21341_, _21336_);
  or (_21343_, _21342_, _05444_);
  nor (_21344_, _11199_, _08358_);
  or (_21345_, _21344_, _21336_);
  or (_21346_, _21345_, _03006_);
  and (_21347_, _03820_, \oc8051_golden_model_1.ACC [2]);
  or (_21348_, _21347_, _21336_);
  and (_21349_, _21348_, _02062_);
  nor (_21351_, _02062_, _21335_);
  or (_21352_, _21351_, _02158_);
  or (_21353_, _21352_, _21349_);
  and (_21354_, _21353_, _02058_);
  and (_21355_, _21354_, _21346_);
  nor (_21356_, _04467_, _21335_);
  and (_21357_, _11194_, _04467_);
  or (_21358_, _21357_, _21356_);
  and (_21359_, _21358_, _02057_);
  or (_21360_, _21359_, _02155_);
  or (_21362_, _21360_, _21355_);
  or (_21363_, _21342_, _02519_);
  and (_21364_, _21363_, _21362_);
  or (_21365_, _21364_, _02153_);
  or (_21366_, _21348_, _02549_);
  and (_21367_, _21366_, _02054_);
  and (_21368_, _21367_, _21365_);
  and (_21369_, _11192_, _04467_);
  or (_21370_, _21369_, _21356_);
  and (_21371_, _21370_, _02053_);
  or (_21373_, _21371_, _02046_);
  or (_21374_, _21373_, _21368_);
  or (_21375_, _21356_, _11223_);
  and (_21376_, _21375_, _21358_);
  or (_21377_, _21376_, _02047_);
  and (_21378_, _21377_, _02043_);
  and (_21379_, _21378_, _21374_);
  and (_21380_, _18983_, _04467_);
  or (_21381_, _21380_, _21356_);
  and (_21382_, _21381_, _02042_);
  or (_21384_, _21382_, _06188_);
  or (_21385_, _21384_, _21379_);
  and (_21386_, _21385_, _21343_);
  or (_21387_, _21386_, _02031_);
  and (_21388_, _05211_, _03820_);
  or (_21389_, _21336_, _02032_);
  or (_21390_, _21389_, _21388_);
  and (_21391_, _21390_, _02037_);
  and (_21392_, _21391_, _21387_);
  and (_21393_, _19008_, _03820_);
  or (_21395_, _21393_, _21336_);
  and (_21396_, _21395_, _01765_);
  or (_21397_, _21396_, _21392_);
  or (_21398_, _21397_, _07629_);
  and (_21399_, _11189_, _03820_);
  or (_21400_, _21336_, _03059_);
  or (_21401_, _21400_, _21399_);
  and (_21402_, _03820_, _04866_);
  or (_21403_, _21402_, _21336_);
  or (_21404_, _21403_, _01995_);
  and (_21406_, _21404_, _03061_);
  and (_21407_, _21406_, _21401_);
  and (_21408_, _21407_, _21398_);
  or (_21409_, _21408_, _21340_);
  and (_21410_, _21409_, _02208_);
  or (_21411_, _21336_, _04309_);
  and (_21412_, _21403_, _02206_);
  and (_21413_, _21412_, _21411_);
  or (_21414_, _21413_, _21410_);
  and (_21415_, _21414_, _03065_);
  and (_21417_, _21348_, _02342_);
  and (_21418_, _21417_, _21411_);
  or (_21419_, _21418_, _02202_);
  or (_21420_, _21419_, _21415_);
  nor (_21421_, _11187_, _08358_);
  or (_21422_, _21336_, _04953_);
  or (_21423_, _21422_, _21421_);
  and (_21424_, _21423_, _04958_);
  and (_21425_, _21424_, _21420_);
  nor (_21426_, _11314_, _08358_);
  or (_21428_, _21426_, _21336_);
  and (_21429_, _21428_, _02334_);
  or (_21430_, _21429_, _02366_);
  or (_21431_, _21430_, _21425_);
  or (_21432_, _21345_, _02778_);
  and (_21433_, _21432_, _01698_);
  and (_21434_, _21433_, _21431_);
  and (_21435_, _21370_, _01697_);
  or (_21436_, _21435_, _02081_);
  or (_21437_, _21436_, _21434_);
  and (_21439_, _11367_, _03820_);
  or (_21440_, _21336_, _02082_);
  or (_21441_, _21440_, _21439_);
  and (_21442_, _21441_, _39632_);
  and (_21443_, _21442_, _21437_);
  nor (_21444_, _39632_, _21335_);
  or (_21445_, _21444_, rst);
  or (_41694_, _21445_, _21443_);
  nor (_21446_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_21447_, _21446_, _00001_);
  and (_21449_, _08358_, \oc8051_golden_model_1.P3 [3]);
  nor (_21450_, _08358_, _03434_);
  or (_21451_, _21450_, _21449_);
  or (_21452_, _21451_, _05444_);
  or (_21453_, _21451_, _02519_);
  nor (_21454_, _11394_, _08358_);
  or (_21455_, _21454_, _21449_);
  or (_21456_, _21455_, _03006_);
  and (_21457_, _03820_, \oc8051_golden_model_1.ACC [3]);
  or (_21458_, _21457_, _21449_);
  and (_21460_, _21458_, _02062_);
  and (_21461_, _02063_, \oc8051_golden_model_1.P3 [3]);
  or (_21462_, _21461_, _02158_);
  or (_21463_, _21462_, _21460_);
  and (_21464_, _21463_, _02058_);
  and (_21465_, _21464_, _21456_);
  not (_21466_, \oc8051_golden_model_1.P3 [3]);
  nor (_21467_, _04467_, _21466_);
  and (_21468_, _11398_, _04467_);
  or (_21469_, _21468_, _21467_);
  and (_21471_, _21469_, _02057_);
  or (_21472_, _21471_, _02155_);
  or (_21473_, _21472_, _21465_);
  and (_21474_, _21473_, _21453_);
  or (_21475_, _21474_, _02153_);
  or (_21476_, _21458_, _02549_);
  and (_21477_, _21476_, _02054_);
  and (_21478_, _21477_, _21475_);
  and (_21479_, _11408_, _04467_);
  or (_21480_, _21479_, _21467_);
  and (_21482_, _21480_, _02053_);
  or (_21483_, _21482_, _02046_);
  or (_21484_, _21483_, _21478_);
  or (_21485_, _21467_, _11415_);
  and (_21486_, _21485_, _21469_);
  or (_21487_, _21486_, _02047_);
  and (_21488_, _21487_, _02043_);
  and (_21489_, _21488_, _21484_);
  and (_21490_, _19106_, _04467_);
  or (_21491_, _21490_, _21467_);
  and (_21493_, _21491_, _02042_);
  or (_21494_, _21493_, _06188_);
  or (_21495_, _21494_, _21489_);
  and (_21496_, _21495_, _21452_);
  or (_21497_, _21496_, _02031_);
  and (_21498_, _05166_, _03820_);
  or (_21499_, _21449_, _02032_);
  or (_21500_, _21499_, _21498_);
  and (_21501_, _21500_, _02037_);
  and (_21502_, _21501_, _21497_);
  and (_21504_, _19131_, _03820_);
  or (_21505_, _21449_, _21504_);
  and (_21506_, _21505_, _01765_);
  or (_21507_, _21506_, _21502_);
  or (_21508_, _21507_, _07629_);
  and (_21509_, _11505_, _03820_);
  or (_21510_, _21449_, _03059_);
  or (_21511_, _21510_, _21509_);
  and (_21512_, _03820_, _04719_);
  or (_21513_, _21512_, _21449_);
  or (_21515_, _21513_, _01995_);
  and (_21516_, _21515_, _03061_);
  and (_21517_, _21516_, _21511_);
  and (_21518_, _21517_, _21508_);
  and (_21519_, _11511_, _03820_);
  or (_21520_, _21519_, _21449_);
  and (_21521_, _21520_, _02331_);
  or (_21522_, _21521_, _21518_);
  and (_21523_, _21522_, _02208_);
  or (_21524_, _21449_, _04153_);
  and (_21526_, _21513_, _02206_);
  and (_21527_, _21526_, _21524_);
  or (_21528_, _21527_, _21523_);
  and (_21529_, _21528_, _03065_);
  and (_21530_, _21458_, _02342_);
  and (_21531_, _21530_, _21524_);
  or (_21532_, _21531_, _02202_);
  or (_21533_, _21532_, _21529_);
  nor (_21534_, _11503_, _08358_);
  or (_21535_, _21449_, _04953_);
  or (_21537_, _21535_, _21534_);
  and (_21538_, _21537_, _04958_);
  and (_21539_, _21538_, _21533_);
  nor (_21540_, _11510_, _08358_);
  or (_21541_, _21540_, _21449_);
  and (_21542_, _21541_, _02334_);
  or (_21543_, _21542_, _02366_);
  or (_21544_, _21543_, _21539_);
  or (_21545_, _21455_, _02778_);
  and (_21546_, _21545_, _01698_);
  and (_21548_, _21546_, _21544_);
  and (_21549_, _21480_, _01697_);
  or (_21550_, _21549_, _02081_);
  or (_21551_, _21550_, _21548_);
  and (_21552_, _11567_, _03820_);
  or (_21553_, _21449_, _02082_);
  or (_21554_, _21553_, _21552_);
  and (_21555_, _21554_, _39632_);
  and (_21556_, _21555_, _21551_);
  or (_41695_, _21556_, _21447_);
  not (_21558_, \oc8051_golden_model_1.P3 [4]);
  nor (_21559_, _03820_, _21558_);
  nor (_21560_, _04372_, _08358_);
  or (_21561_, _21560_, _21559_);
  or (_21562_, _21561_, _05444_);
  or (_21563_, _21561_, _02519_);
  nor (_21564_, _11611_, _08358_);
  or (_21565_, _21564_, _21559_);
  or (_21566_, _21565_, _03006_);
  and (_21567_, _03820_, \oc8051_golden_model_1.ACC [4]);
  or (_21569_, _21567_, _21559_);
  and (_21570_, _21569_, _02062_);
  nor (_21571_, _02062_, _21558_);
  or (_21572_, _21571_, _02158_);
  or (_21573_, _21572_, _21570_);
  and (_21574_, _21573_, _02058_);
  and (_21575_, _21574_, _21566_);
  nor (_21576_, _04467_, _21558_);
  and (_21577_, _11597_, _04467_);
  or (_21578_, _21577_, _21576_);
  and (_21580_, _21578_, _02057_);
  or (_21581_, _21580_, _02155_);
  or (_21582_, _21581_, _21575_);
  and (_21583_, _21582_, _21563_);
  or (_21584_, _21583_, _02153_);
  or (_21585_, _21569_, _02549_);
  and (_21586_, _21585_, _02054_);
  and (_21587_, _21586_, _21584_);
  and (_21588_, _11595_, _04467_);
  or (_21589_, _21588_, _21576_);
  and (_21591_, _21589_, _02053_);
  or (_21592_, _21591_, _02046_);
  or (_21593_, _21592_, _21587_);
  or (_21594_, _21576_, _11628_);
  and (_21595_, _21594_, _21578_);
  or (_21596_, _21595_, _02047_);
  and (_21597_, _21596_, _02043_);
  and (_21598_, _21597_, _21593_);
  and (_21599_, _19230_, _04467_);
  or (_21600_, _21599_, _21576_);
  and (_21602_, _21600_, _02042_);
  or (_21603_, _21602_, _06188_);
  or (_21604_, _21603_, _21598_);
  and (_21605_, _21604_, _21562_);
  or (_21606_, _21605_, _02031_);
  and (_21607_, _05303_, _03820_);
  or (_21608_, _21559_, _02032_);
  or (_21609_, _21608_, _21607_);
  and (_21610_, _21609_, _02037_);
  and (_21611_, _21610_, _21606_);
  and (_21613_, _19257_, _03820_);
  or (_21614_, _21559_, _21613_);
  and (_21615_, _21614_, _01765_);
  or (_21616_, _21615_, _21611_);
  or (_21617_, _21616_, _07629_);
  and (_21618_, _11592_, _03820_);
  or (_21619_, _21559_, _03059_);
  or (_21620_, _21619_, _21618_);
  and (_21621_, _04831_, _03820_);
  or (_21622_, _21621_, _21559_);
  or (_21624_, _21622_, _01995_);
  and (_21625_, _21624_, _03061_);
  and (_21626_, _21625_, _21620_);
  and (_21627_, _21626_, _21617_);
  and (_21628_, _11588_, _03820_);
  or (_21629_, _21628_, _21559_);
  and (_21630_, _21629_, _02331_);
  or (_21631_, _21630_, _21627_);
  and (_21632_, _21631_, _02208_);
  or (_21633_, _21559_, _04420_);
  and (_21635_, _21622_, _02206_);
  and (_21636_, _21635_, _21633_);
  or (_21637_, _21636_, _21632_);
  and (_21638_, _21637_, _03065_);
  and (_21639_, _21569_, _02342_);
  and (_21640_, _21639_, _21633_);
  or (_21641_, _21640_, _02202_);
  or (_21642_, _21641_, _21638_);
  nor (_21643_, _11590_, _08358_);
  or (_21644_, _21559_, _04953_);
  or (_21646_, _21644_, _21643_);
  and (_21647_, _21646_, _04958_);
  and (_21648_, _21647_, _21642_);
  nor (_21649_, _11587_, _08358_);
  or (_21650_, _21649_, _21559_);
  and (_21651_, _21650_, _02334_);
  or (_21652_, _21651_, _02366_);
  or (_21653_, _21652_, _21648_);
  or (_21654_, _21565_, _02778_);
  and (_21655_, _21654_, _01698_);
  and (_21657_, _21655_, _21653_);
  and (_21658_, _21589_, _01697_);
  or (_21659_, _21658_, _02081_);
  or (_21660_, _21659_, _21657_);
  and (_21661_, _11771_, _03820_);
  or (_21662_, _21559_, _02082_);
  or (_21663_, _21662_, _21661_);
  and (_21664_, _21663_, _39632_);
  and (_21665_, _21664_, _21660_);
  nor (_21666_, _39632_, _21558_);
  or (_21668_, _21666_, rst);
  or (_41697_, _21668_, _21665_);
  not (_21669_, \oc8051_golden_model_1.P3 [5]);
  nor (_21670_, _03820_, _21669_);
  nor (_21671_, _04057_, _08358_);
  or (_21672_, _21671_, _21670_);
  or (_21673_, _21672_, _05444_);
  or (_21674_, _21672_, _02519_);
  nor (_21675_, _11804_, _08358_);
  or (_21676_, _21675_, _21670_);
  or (_21678_, _21676_, _03006_);
  and (_21679_, _03820_, \oc8051_golden_model_1.ACC [5]);
  or (_21680_, _21679_, _21670_);
  and (_21681_, _21680_, _02062_);
  nor (_21682_, _02062_, _21669_);
  or (_21683_, _21682_, _02158_);
  or (_21684_, _21683_, _21681_);
  and (_21685_, _21684_, _02058_);
  and (_21686_, _21685_, _21678_);
  nor (_21687_, _04467_, _21669_);
  and (_21689_, _11789_, _04467_);
  or (_21690_, _21689_, _21687_);
  and (_21691_, _21690_, _02057_);
  or (_21692_, _21691_, _02155_);
  or (_21693_, _21692_, _21686_);
  and (_21694_, _21693_, _21674_);
  or (_21695_, _21694_, _02153_);
  or (_21696_, _21680_, _02549_);
  and (_21697_, _21696_, _02054_);
  and (_21698_, _21697_, _21695_);
  and (_21700_, _11816_, _04467_);
  or (_21701_, _21700_, _21687_);
  and (_21702_, _21701_, _02053_);
  or (_21703_, _21702_, _02046_);
  or (_21704_, _21703_, _21698_);
  or (_21705_, _21687_, _11823_);
  and (_21706_, _21705_, _21690_);
  or (_21707_, _21706_, _02047_);
  and (_21708_, _21707_, _02043_);
  and (_21709_, _21708_, _21704_);
  and (_21711_, _19358_, _04467_);
  or (_21712_, _21711_, _21687_);
  and (_21713_, _21712_, _02042_);
  or (_21714_, _21713_, _06188_);
  or (_21715_, _21714_, _21709_);
  and (_21716_, _21715_, _21673_);
  or (_21717_, _21716_, _02031_);
  and (_21718_, _05258_, _03820_);
  or (_21719_, _21670_, _02032_);
  or (_21720_, _21719_, _21718_);
  and (_21722_, _21720_, _02037_);
  and (_21723_, _21722_, _21717_);
  and (_21724_, _19394_, _03820_);
  or (_21725_, _21724_, _21670_);
  and (_21726_, _21725_, _01765_);
  or (_21727_, _21726_, _21723_);
  or (_21728_, _21727_, _07629_);
  and (_21729_, _11915_, _03820_);
  or (_21730_, _21670_, _03059_);
  or (_21731_, _21730_, _21729_);
  and (_21733_, _04827_, _03820_);
  or (_21734_, _21733_, _21670_);
  or (_21735_, _21734_, _01995_);
  and (_21736_, _21735_, _03061_);
  and (_21737_, _21736_, _21731_);
  and (_21738_, _21737_, _21728_);
  and (_21739_, _11786_, _03820_);
  or (_21740_, _21739_, _21670_);
  and (_21741_, _21740_, _02331_);
  or (_21742_, _21741_, _21738_);
  and (_21744_, _21742_, _02208_);
  or (_21745_, _21670_, _04104_);
  and (_21746_, _21734_, _02206_);
  and (_21747_, _21746_, _21745_);
  or (_21748_, _21747_, _21744_);
  and (_21749_, _21748_, _03065_);
  and (_21750_, _21680_, _02342_);
  and (_21751_, _21750_, _21745_);
  or (_21752_, _21751_, _02202_);
  or (_21753_, _21752_, _21749_);
  nor (_21755_, _11913_, _08358_);
  or (_21756_, _21670_, _04953_);
  or (_21757_, _21756_, _21755_);
  and (_21758_, _21757_, _04958_);
  and (_21759_, _21758_, _21753_);
  nor (_21760_, _11785_, _08358_);
  or (_21761_, _21760_, _21670_);
  and (_21762_, _21761_, _02334_);
  or (_21763_, _21762_, _02366_);
  or (_21764_, _21763_, _21759_);
  or (_21766_, _21676_, _02778_);
  and (_21767_, _21766_, _01698_);
  and (_21768_, _21767_, _21764_);
  and (_21769_, _21701_, _01697_);
  or (_21770_, _21769_, _02081_);
  or (_21771_, _21770_, _21768_);
  and (_21772_, _11974_, _03820_);
  or (_21773_, _21670_, _02082_);
  or (_21774_, _21773_, _21772_);
  and (_21775_, _21774_, _39632_);
  and (_21777_, _21775_, _21771_);
  nor (_21778_, _39632_, _21669_);
  or (_21779_, _21778_, rst);
  or (_41698_, _21779_, _21777_);
  not (_21780_, \oc8051_golden_model_1.P3 [6]);
  nor (_21781_, _39632_, _21780_);
  or (_21782_, _21781_, rst);
  nor (_21783_, _03820_, _21780_);
  nor (_21784_, _03964_, _08358_);
  or (_21785_, _21784_, _21783_);
  or (_21787_, _21785_, _05444_);
  or (_21788_, _21785_, _02519_);
  nor (_21789_, _11993_, _08358_);
  or (_21790_, _21789_, _21783_);
  or (_21791_, _21790_, _03006_);
  and (_21792_, _03820_, \oc8051_golden_model_1.ACC [6]);
  or (_21793_, _21792_, _21783_);
  and (_21794_, _21793_, _02062_);
  nor (_21795_, _02062_, _21780_);
  or (_21796_, _21795_, _02158_);
  or (_21798_, _21796_, _21794_);
  and (_21799_, _21798_, _02058_);
  and (_21800_, _21799_, _21791_);
  nor (_21801_, _04467_, _21780_);
  and (_21802_, _11990_, _04467_);
  or (_21803_, _21802_, _21801_);
  and (_21804_, _21803_, _02057_);
  or (_21805_, _21804_, _02155_);
  or (_21806_, _21805_, _21800_);
  and (_21807_, _21806_, _21788_);
  or (_21809_, _21807_, _02153_);
  or (_21810_, _21793_, _02549_);
  and (_21811_, _21810_, _02054_);
  and (_21812_, _21811_, _21809_);
  and (_21813_, _12017_, _04467_);
  or (_21814_, _21813_, _21801_);
  and (_21815_, _21814_, _02053_);
  or (_21816_, _21815_, _02046_);
  or (_21817_, _21816_, _21812_);
  or (_21818_, _21801_, _12024_);
  and (_21820_, _21818_, _21803_);
  or (_21821_, _21820_, _02047_);
  and (_21822_, _21821_, _02043_);
  and (_21823_, _21822_, _21817_);
  and (_21824_, _19493_, _04467_);
  or (_21825_, _21824_, _21801_);
  and (_21826_, _21825_, _02042_);
  or (_21827_, _21826_, _06188_);
  or (_21828_, _21827_, _21823_);
  and (_21829_, _21828_, _21787_);
  or (_21831_, _21829_, _02031_);
  and (_21832_, _05029_, _03820_);
  or (_21833_, _21783_, _02032_);
  or (_21834_, _21833_, _21832_);
  and (_21835_, _21834_, _02037_);
  and (_21836_, _21835_, _21831_);
  and (_21837_, _19520_, _03820_);
  or (_21838_, _21837_, _21783_);
  and (_21839_, _21838_, _01765_);
  or (_21840_, _21839_, _21836_);
  or (_21842_, _21840_, _07629_);
  and (_21843_, _12112_, _03820_);
  or (_21844_, _21783_, _03059_);
  or (_21845_, _21844_, _21843_);
  and (_21846_, _12103_, _03820_);
  or (_21847_, _21846_, _21783_);
  or (_21848_, _21847_, _01995_);
  and (_21849_, _21848_, _03061_);
  and (_21850_, _21849_, _21845_);
  and (_21851_, _21850_, _21842_);
  and (_21853_, _12118_, _03820_);
  or (_21854_, _21853_, _21783_);
  and (_21855_, _21854_, _02331_);
  or (_21856_, _21855_, _21851_);
  and (_21857_, _21856_, _02208_);
  or (_21858_, _21783_, _04011_);
  and (_21859_, _21847_, _02206_);
  and (_21860_, _21859_, _21858_);
  or (_21861_, _21860_, _21857_);
  and (_21862_, _21861_, _03065_);
  and (_21864_, _21793_, _02342_);
  and (_21865_, _21864_, _21858_);
  or (_21866_, _21865_, _02202_);
  or (_21867_, _21866_, _21862_);
  nor (_21868_, _12110_, _08358_);
  or (_21869_, _21783_, _04953_);
  or (_21870_, _21869_, _21868_);
  and (_21871_, _21870_, _04958_);
  and (_21872_, _21871_, _21867_);
  nor (_21873_, _12117_, _08358_);
  or (_21875_, _21873_, _21783_);
  and (_21876_, _21875_, _02334_);
  or (_21877_, _21876_, _02366_);
  or (_21878_, _21877_, _21872_);
  or (_21879_, _21790_, _02778_);
  and (_21880_, _21879_, _01698_);
  and (_21881_, _21880_, _21878_);
  and (_21882_, _21814_, _01697_);
  or (_21883_, _21882_, _02081_);
  or (_21884_, _21883_, _21881_);
  and (_21886_, _12178_, _03820_);
  or (_21887_, _21783_, _02082_);
  or (_21888_, _21887_, _21886_);
  and (_21889_, _21888_, _39632_);
  and (_21890_, _21889_, _21884_);
  or (_41699_, _21890_, _21782_);
  not (_21891_, \oc8051_golden_model_1.PSW [0]);
  nor (_21892_, _39632_, _21891_);
  nor (_21893_, _06324_, _06323_);
  nor (_21894_, _21893_, _06231_);
  and (_21896_, _21893_, _06231_);
  nor (_21897_, _21896_, _21894_);
  nor (_21898_, _06248_, _06247_);
  nor (_21899_, _21898_, _14194_);
  and (_21900_, _21898_, _14194_);
  nor (_21901_, _21900_, _21899_);
  and (_21902_, _21901_, _21897_);
  nor (_21903_, _21901_, _21897_);
  nor (_21904_, _21903_, _21902_);
  nor (_21905_, _21904_, _04939_);
  and (_21907_, _21904_, _04939_);
  nor (_21908_, _21907_, _21905_);
  or (_21909_, _21908_, _05337_);
  not (_21910_, _07582_);
  and (_21911_, _14235_, _21910_);
  and (_21912_, _21911_, \oc8051_golden_model_1.ACC [3]);
  nor (_21913_, _21911_, \oc8051_golden_model_1.ACC [3]);
  nor (_21914_, _21913_, _21912_);
  and (_21915_, _21914_, _15145_);
  nor (_21916_, _21914_, _15145_);
  nor (_21918_, _21916_, _21915_);
  and (_21919_, _15461_, _06231_);
  nor (_21920_, _15461_, _06231_);
  nor (_21921_, _21920_, _21919_);
  nor (_21922_, _21921_, _21918_);
  and (_21923_, _21921_, _21918_);
  or (_21924_, _21923_, _21922_);
  nor (_21925_, _21924_, _07588_);
  and (_21926_, _21924_, _07588_);
  nor (_21927_, _21926_, _21925_);
  and (_21929_, _21927_, _07575_);
  nor (_21930_, _21929_, _07580_);
  nor (_21931_, _10629_, _01722_);
  or (_21932_, _21931_, _21908_);
  not (_21933_, _14627_);
  and (_21934_, _21933_, _14281_);
  nor (_21935_, _21933_, _14281_);
  nor (_21936_, _21935_, _21934_);
  not (_21937_, _21936_);
  not (_21938_, _15255_);
  and (_21940_, _21938_, _14914_);
  nor (_21941_, _21938_, _14914_);
  nor (_21942_, _21941_, _21940_);
  and (_21943_, _21942_, _21937_);
  nor (_21944_, _21942_, _21937_);
  nor (_21945_, _21944_, _21943_);
  and (_21946_, _14010_, _13714_);
  nor (_21947_, _14010_, _13714_);
  or (_21948_, _21947_, _21946_);
  and (_21949_, _21948_, _15568_);
  nor (_21951_, _21948_, _15568_);
  nor (_21952_, _21951_, _21949_);
  and (_21953_, _21952_, _21945_);
  nor (_21954_, _21952_, _21945_);
  nor (_21955_, _21954_, _21953_);
  and (_21956_, _21955_, _06896_);
  nor (_21957_, _21955_, _06896_);
  or (_21958_, _21957_, _21956_);
  and (_21959_, _21958_, _02053_);
  and (_21960_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  nor (_21962_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [0]);
  or (_21963_, _21962_, _21960_);
  and (_21964_, _21963_, _13964_);
  nor (_21965_, _21963_, _13964_);
  nor (_21966_, _21965_, _21964_);
  and (_21967_, _14872_, _14603_);
  and (_21968_, _14871_, _14604_);
  nor (_21969_, _21968_, _21967_);
  nor (_21970_, _21969_, _21966_);
  and (_21971_, _21969_, _21966_);
  nor (_21973_, _21971_, _21970_);
  and (_21974_, _21973_, _15215_);
  nor (_21975_, _21973_, _15215_);
  nor (_21976_, _21975_, _21974_);
  nor (_21977_, _15525_, _06843_);
  and (_21978_, _15525_, _06843_);
  nor (_21979_, _21978_, _21977_);
  nor (_21980_, _21979_, _21976_);
  and (_21981_, _21979_, _21976_);
  nor (_21982_, _21981_, _21980_);
  nand (_21984_, _21982_, _06823_);
  nor (_21985_, _07094_, _07036_);
  and (_21986_, _07094_, _07036_);
  nor (_21987_, _21986_, _21985_);
  nor (_21988_, _07082_, _07068_);
  and (_21989_, _07082_, _07068_);
  nor (_21990_, _21989_, _21988_);
  nor (_21991_, _21990_, _21987_);
  and (_21992_, _21990_, _21987_);
  or (_21993_, _21992_, _21991_);
  and (_21995_, _07126_, _07115_);
  nor (_21996_, _21995_, _07127_);
  nor (_21997_, _21996_, _07057_);
  and (_21998_, _21996_, _07057_);
  nor (_21999_, _21998_, _21997_);
  nor (_22000_, _21999_, _21993_);
  and (_22001_, _21999_, _21993_);
  nor (_22002_, _22001_, _22000_);
  nor (_22003_, _22002_, _09067_);
  and (_22004_, _22002_, _09067_);
  or (_22006_, _22004_, _22003_);
  and (_22007_, _22006_, _02160_);
  nor (_22008_, _05365_, _05212_);
  not (_22009_, _22008_);
  nand (_22010_, _22009_, _10983_);
  or (_22011_, _22009_, _10983_);
  and (_22012_, _22011_, _22010_);
  not (_22013_, _22012_);
  nor (_22014_, _05367_, _05304_);
  nand (_22015_, _22014_, _05029_);
  or (_22017_, _22014_, _05029_);
  and (_22018_, _22017_, _22015_);
  nand (_22019_, _22018_, _22013_);
  or (_22020_, _22018_, _22013_);
  nand (_22021_, _22020_, _22019_);
  nor (_22022_, _22021_, _04637_);
  and (_22023_, _22021_, _04637_);
  or (_22024_, _22023_, _22022_);
  or (_22025_, _22024_, _06849_);
  and (_22026_, _05351_, _04057_);
  nor (_22028_, _05351_, _04057_);
  nor (_22029_, _22028_, _22026_);
  nor (_22030_, _05345_, _04526_);
  not (_22031_, _22030_);
  and (_22032_, _10981_, _05343_);
  nor (_22033_, _10981_, _05343_);
  nor (_22034_, _22033_, _22032_);
  and (_22035_, _22034_, _22031_);
  nor (_22036_, _22034_, _22031_);
  nor (_22037_, _22036_, _22035_);
  nor (_22039_, _22037_, _22029_);
  and (_22040_, _22037_, _22029_);
  or (_22041_, _22040_, _22039_);
  nor (_22042_, _22041_, _06852_);
  and (_22043_, _10312_, _09495_);
  and (_22044_, _22043_, _21891_);
  nor (_22045_, _22043_, _21908_);
  or (_22046_, _22045_, _06853_);
  or (_22047_, _22046_, _22044_);
  nand (_22048_, _22047_, _06849_);
  or (_22050_, _22048_, _22042_);
  and (_22051_, _22050_, _06847_);
  and (_22052_, _22051_, _22025_);
  or (_22053_, _22052_, _22007_);
  and (_22054_, _04534_, _01752_);
  and (_22055_, _22054_, _10299_);
  and (_22056_, _22055_, _22053_);
  not (_22057_, _21908_);
  nor (_22058_, _22054_, _22057_);
  or (_22059_, _22058_, _02079_);
  or (_22061_, _22059_, _22056_);
  nor (_22062_, _21898_, \oc8051_golden_model_1.ACC [6]);
  and (_22063_, _21898_, \oc8051_golden_model_1.ACC [6]);
  nor (_22064_, _22063_, _22062_);
  nor (_22065_, _22064_, \oc8051_golden_model_1.ACC [7]);
  and (_22066_, _22064_, \oc8051_golden_model_1.ACC [7]);
  nor (_22067_, _22066_, _22065_);
  and (_22068_, _22067_, _22012_);
  nor (_22069_, _22067_, _22012_);
  or (_22070_, _22069_, _22068_);
  or (_22072_, _22070_, _04550_);
  and (_22073_, _22072_, _03006_);
  and (_22074_, _22073_, _22061_);
  not (_22075_, _14887_);
  and (_22076_, _22075_, _14596_);
  nor (_22077_, _22075_, _14596_);
  nor (_22078_, _22077_, _22076_);
  and (_22079_, _22078_, _15541_);
  nor (_22080_, _22078_, _15541_);
  nor (_22081_, _22080_, _22079_);
  not (_22083_, _13743_);
  nor (_22084_, _13983_, _22083_);
  and (_22085_, _13983_, _22083_);
  nor (_22086_, _22085_, _22084_);
  and (_22087_, _22086_, _14254_);
  nor (_22088_, _22086_, _14254_);
  nor (_22089_, _22088_, _22087_);
  and (_22090_, _22089_, _15230_);
  nor (_22091_, _22089_, _15230_);
  or (_22092_, _22091_, _22090_);
  and (_22094_, _22092_, _06867_);
  nor (_22095_, _22092_, _06867_);
  or (_22096_, _22095_, _22094_);
  and (_22097_, _22096_, _22081_);
  nor (_22098_, _22096_, _22081_);
  or (_22099_, _22098_, _22097_);
  and (_22100_, _22099_, _02158_);
  or (_22101_, _22100_, _06823_);
  or (_22102_, _22101_, _22074_);
  and (_22103_, _22102_, _21984_);
  or (_22105_, _22103_, _08707_);
  nand (_22106_, _22057_, _08707_);
  and (_22107_, _22106_, _02058_);
  and (_22108_, _22107_, _22105_);
  and (_22109_, _13991_, _13749_);
  nor (_22110_, _13991_, _13749_);
  or (_22111_, _22110_, _22109_);
  nor (_22112_, _14608_, _14262_);
  and (_22113_, _14608_, _14262_);
  nor (_22114_, _22113_, _22112_);
  not (_22116_, _22114_);
  and (_22117_, _22116_, _22111_);
  nor (_22118_, _22116_, _22111_);
  nor (_22119_, _22118_, _22117_);
  not (_22120_, _15549_);
  nor (_22121_, _15236_, _14895_);
  and (_22122_, _15236_, _14895_);
  nor (_22123_, _22122_, _22121_);
  nor (_22124_, _22123_, _22120_);
  and (_22125_, _22123_, _22120_);
  nor (_22127_, _22125_, _22124_);
  nor (_22128_, _22127_, _22119_);
  and (_22129_, _22127_, _22119_);
  nor (_22130_, _22129_, _22128_);
  and (_22131_, _22130_, _06875_);
  nor (_22132_, _22130_, _06875_);
  or (_22133_, _22132_, _22131_);
  and (_22134_, _22133_, _02057_);
  or (_22135_, _22134_, _22108_);
  and (_22136_, _22135_, _01745_);
  nor (_22138_, _22057_, _01745_);
  or (_22139_, _22138_, _22136_);
  or (_22140_, _22139_, _02155_);
  and (_22141_, _13959_, _13723_);
  nor (_22142_, _13959_, _13723_);
  nor (_22143_, _22142_, _22141_);
  and (_22144_, _22143_, _14230_);
  nor (_22145_, _22143_, _14230_);
  or (_22146_, _22145_, _22144_);
  nand (_22147_, _22146_, _14556_);
  or (_22149_, _22146_, _14556_);
  and (_22150_, _22149_, _22147_);
  not (_22151_, _15495_);
  nor (_22152_, _15189_, _14867_);
  and (_22153_, _15189_, _14867_);
  nor (_22154_, _22153_, _22152_);
  nor (_22155_, _22154_, _22151_);
  and (_22156_, _22154_, _22151_);
  nor (_22157_, _22156_, _22155_);
  not (_22158_, _22157_);
  nor (_22160_, _22158_, _22150_);
  and (_22161_, _22158_, _22150_);
  nor (_22162_, _22161_, _22160_);
  and (_22163_, _22162_, _06738_);
  nor (_22164_, _22162_, _06738_);
  or (_22165_, _22164_, _22163_);
  or (_22166_, _22165_, _02519_);
  and (_22167_, _22166_, _06820_);
  and (_22168_, _22167_, _22140_);
  not (_22169_, _10452_);
  nand (_22171_, _22041_, _06884_);
  and (_22172_, _22171_, _22169_);
  or (_22173_, _22172_, _22168_);
  or (_22174_, _22024_, _06884_);
  and (_22175_, _22174_, _02549_);
  and (_22176_, _22175_, _22173_);
  and (_22177_, _22006_, _02153_);
  or (_22178_, _22177_, _10462_);
  or (_22179_, _22178_, _22176_);
  or (_22180_, _21908_, _10460_);
  and (_22182_, _22180_, _02054_);
  and (_22183_, _22182_, _22179_);
  or (_22184_, _22183_, _21959_);
  not (_22185_, _10465_);
  nor (_22186_, _10470_, _22185_);
  and (_22187_, _22186_, _22184_);
  and (_22188_, _08692_, _08836_);
  nor (_22189_, _08881_, _02230_);
  and (_22190_, _22189_, _22188_);
  or (_22191_, _22186_, _22057_);
  nand (_22193_, _22191_, _22190_);
  or (_22194_, _22193_, _22187_);
  or (_22195_, _22190_, _21908_);
  and (_22196_, _22195_, _02047_);
  and (_22197_, _22196_, _22194_);
  not (_22198_, _15210_);
  nor (_22199_, _14286_, _14015_);
  and (_22200_, _14286_, _14015_);
  nor (_22201_, _22200_, _22199_);
  nor (_22202_, _22201_, _22198_);
  and (_22204_, _22201_, _22198_);
  nor (_22205_, _22204_, _22202_);
  nor (_22206_, _14578_, _22083_);
  and (_22207_, _14578_, _22083_);
  nor (_22208_, _22207_, _22206_);
  and (_22209_, _22208_, _14919_);
  nor (_22210_, _22208_, _14919_);
  nor (_22211_, _22210_, _22209_);
  nor (_22212_, _15573_, _06901_);
  and (_22213_, _15573_, _06901_);
  nor (_22215_, _22213_, _22212_);
  not (_22216_, _22215_);
  nor (_22217_, _22216_, _22211_);
  and (_22218_, _22216_, _22211_);
  nor (_22219_, _22218_, _22217_);
  not (_22220_, _22219_);
  nand (_22221_, _22220_, _22205_);
  or (_22222_, _22220_, _22205_);
  and (_22223_, _22222_, _02046_);
  and (_22224_, _22223_, _22221_);
  or (_22226_, _22224_, _22197_);
  not (_22227_, _02139_);
  nor (_22228_, _03316_, _02142_);
  and (_22229_, _22228_, _22227_);
  and (_22230_, _22229_, _10501_);
  and (_22231_, _22230_, _22226_);
  nor (_22232_, _02730_, _01754_);
  or (_22233_, _22232_, _10155_);
  nor (_22234_, _22230_, _22057_);
  or (_22235_, _22234_, _22233_);
  or (_22237_, _22235_, _22231_);
  nand (_22238_, _22233_, _22057_);
  and (_22239_, _22238_, _06181_);
  and (_22240_, _22239_, _22237_);
  nor (_22241_, _14020_, _06127_);
  nor (_22242_, _14021_, _13773_);
  nor (_22243_, _22242_, _22241_);
  nor (_22244_, _22243_, _14291_);
  and (_22245_, _22243_, _14291_);
  nor (_22246_, _22245_, _22244_);
  nor (_22248_, _22246_, _14634_);
  and (_22249_, _22246_, _14634_);
  or (_22250_, _22249_, _22248_);
  not (_22251_, _22250_);
  nor (_22252_, _22251_, _14924_);
  and (_22253_, _22251_, _14924_);
  nor (_22254_, _22253_, _22252_);
  nor (_22255_, _22254_, _15262_);
  and (_22256_, _22254_, _15262_);
  or (_22257_, _22256_, _22255_);
  and (_22259_, _22257_, _15578_);
  nor (_22260_, _22257_, _15578_);
  nor (_22261_, _22260_, _22259_);
  or (_22262_, _22261_, _06906_);
  nand (_22263_, _22261_, _06906_);
  and (_22264_, _22263_, _05474_);
  nand (_22265_, _22264_, _22262_);
  nor (_22266_, _02182_, _10513_);
  and (_22267_, _22266_, _07649_);
  and (_22268_, _22267_, _09032_);
  nand (_22270_, _22268_, _22265_);
  or (_22271_, _22270_, _22240_);
  or (_22272_, _22268_, _21908_);
  and (_22273_, _22272_, _06816_);
  and (_22274_, _22273_, _22271_);
  not (_22275_, _14941_);
  not (_22276_, _06924_);
  and (_22277_, _14030_, _22276_);
  or (_22278_, _22277_, _06925_);
  nor (_22279_, _22278_, _14309_);
  and (_22281_, _22278_, _14309_);
  nor (_22282_, _22281_, _22279_);
  and (_22283_, _22282_, _14648_);
  nor (_22284_, _22282_, _14648_);
  or (_22285_, _22284_, _22283_);
  and (_22286_, _22285_, _22275_);
  nor (_22287_, _22285_, _22275_);
  nor (_22288_, _22287_, _22286_);
  or (_22289_, _22288_, _15278_);
  nand (_22290_, _22288_, _15278_);
  and (_22292_, _22290_, _22289_);
  nor (_22293_, _22292_, _15593_);
  and (_22294_, _22292_, _15593_);
  nor (_22295_, _22294_, _22293_);
  nor (_22296_, _22295_, _06938_);
  and (_22297_, _06937_, _06817_);
  and (_22298_, _22297_, _22295_);
  or (_22299_, _22298_, _06815_);
  or (_22300_, _22299_, _22296_);
  or (_22301_, _22300_, _22274_);
  not (_22303_, _07002_);
  and (_22304_, _14038_, _22303_);
  or (_22305_, _22304_, _07003_);
  nor (_22306_, _22305_, _14326_);
  and (_22307_, _22305_, _14326_);
  nor (_22308_, _22307_, _22306_);
  nor (_22309_, _22308_, _14573_);
  and (_22310_, _22308_, _14573_);
  nor (_22311_, _22310_, _22309_);
  or (_22312_, _22311_, _14961_);
  nand (_22314_, _22311_, _14961_);
  and (_22315_, _22314_, _22312_);
  nor (_22316_, _22315_, _15205_);
  and (_22317_, _22315_, _15205_);
  or (_22318_, _22317_, _22316_);
  nor (_22319_, _22318_, _15519_);
  and (_22320_, _22318_, _15519_);
  nor (_22321_, _22320_, _22319_);
  or (_22322_, _22321_, _07013_);
  and (_22323_, _07012_, _06815_);
  nand (_22325_, _22323_, _22321_);
  and (_22326_, _22325_, _02191_);
  and (_22327_, _22326_, _22322_);
  and (_22328_, _22327_, _22301_);
  not (_22329_, _15294_);
  or (_22330_, _07196_, _07186_);
  and (_22331_, _22330_, _07197_);
  nor (_22332_, _22331_, _14339_);
  and (_22333_, _22331_, _14339_);
  nor (_22334_, _22333_, _22332_);
  nor (_22336_, _22334_, _14664_);
  and (_22337_, _22334_, _14664_);
  or (_22338_, _22337_, _22336_);
  and (_22339_, _22338_, _14973_);
  nor (_22340_, _22338_, _14973_);
  or (_22341_, _22340_, _22339_);
  and (_22342_, _22341_, _22329_);
  nor (_22343_, _22341_, _22329_);
  nor (_22344_, _22343_, _22342_);
  and (_22345_, _22344_, _15505_);
  nor (_22347_, _22344_, _15505_);
  nor (_22348_, _22347_, _22345_);
  and (_22349_, _22348_, _07206_);
  nor (_22350_, _22348_, _07206_);
  or (_22351_, _22350_, _22349_);
  and (_22352_, _22351_, _02186_);
  or (_22353_, _22352_, _22328_);
  and (_22354_, _22353_, _06741_);
  not (_22355_, _06792_);
  and (_22356_, _14049_, _22355_);
  nor (_22358_, _14049_, _22355_);
  nor (_22359_, _22358_, _22356_);
  not (_22360_, _22359_);
  nor (_22361_, _22360_, _14352_);
  and (_22362_, _22360_, _14352_);
  nor (_22363_, _22362_, _22361_);
  and (_22364_, _22363_, _14678_);
  nor (_22365_, _22363_, _14678_);
  or (_22366_, _22365_, _22364_);
  or (_22367_, _22366_, _14988_);
  nand (_22369_, _22366_, _14988_);
  and (_22370_, _22369_, _22367_);
  nor (_22371_, _22370_, _15310_);
  and (_22372_, _22370_, _15310_);
  or (_22373_, _22372_, _22371_);
  nor (_22374_, _22373_, _15609_);
  and (_22375_, _22373_, _15609_);
  nor (_22376_, _22375_, _22374_);
  nand (_22377_, _22376_, _06813_);
  or (_22378_, _22376_, _06813_);
  and (_22380_, _22378_, _22377_);
  and (_22381_, _22380_, _06740_);
  or (_22382_, _22381_, _01876_);
  or (_22383_, _22382_, _22354_);
  nor (_22384_, _03798_, _02119_);
  nor (_22385_, _03811_, _03800_);
  nor (_22386_, _03807_, _03826_);
  nor (_22387_, _03816_, _03852_);
  nor (_22388_, _22387_, _22386_);
  and (_22389_, _22387_, _22386_);
  nor (_22391_, _22389_, _22388_);
  nor (_22392_, _22391_, _22385_);
  and (_22393_, _22391_, _22385_);
  nor (_22394_, _22393_, _22392_);
  not (_22395_, _22394_);
  nor (_22396_, _22395_, _22384_);
  and (_22397_, _22395_, _22384_);
  or (_22398_, _22397_, _22396_);
  or (_22399_, _22398_, _01778_);
  and (_22400_, _22399_, _02043_);
  and (_22402_, _22400_, _22383_);
  not (_22403_, _07217_);
  and (_22404_, _14057_, _13792_);
  nor (_22405_, _14057_, _13792_);
  or (_22406_, _22405_, _22404_);
  nor (_22407_, _14686_, _14360_);
  and (_22408_, _14686_, _14360_);
  nor (_22409_, _22408_, _22407_);
  not (_22410_, _22409_);
  and (_22411_, _22410_, _22406_);
  nor (_22413_, _22410_, _22406_);
  nor (_22414_, _22413_, _22411_);
  not (_22415_, _15617_);
  nor (_22416_, _15318_, _14996_);
  and (_22417_, _15318_, _14996_);
  nor (_22418_, _22417_, _22416_);
  nor (_22419_, _22418_, _22415_);
  and (_22420_, _22418_, _22415_);
  nor (_22421_, _22420_, _22419_);
  nor (_22422_, _22421_, _22414_);
  and (_22424_, _22421_, _22414_);
  nor (_22425_, _22424_, _22422_);
  nand (_22426_, _22425_, _22403_);
  and (_22427_, _22425_, _02042_);
  or (_22428_, _22427_, _07218_);
  and (_22429_, _22428_, _22426_);
  nor (_22430_, _02218_, _01767_);
  not (_22431_, _22430_);
  or (_22432_, _22431_, _22429_);
  or (_22433_, _22432_, _22402_);
  or (_22435_, _22430_, _21908_);
  and (_22436_, _22435_, _05444_);
  and (_22437_, _22436_, _22433_);
  and (_22438_, _22165_, _06188_);
  or (_22439_, _22438_, _02031_);
  or (_22440_, _22439_, _22437_);
  and (_22441_, _14064_, _13799_);
  nor (_22442_, _14064_, _13799_);
  nor (_22443_, _22442_, _22441_);
  and (_22444_, _22443_, _14367_);
  nor (_22446_, _22443_, _14367_);
  or (_22447_, _22446_, _22444_);
  and (_22448_, _22447_, _14693_);
  nor (_22449_, _22447_, _14693_);
  or (_22450_, _22449_, _22448_);
  not (_22451_, _15325_);
  and (_22452_, _22451_, _15003_);
  nor (_22453_, _22451_, _15003_);
  nor (_22454_, _22453_, _22452_);
  nand (_22455_, _22454_, _15624_);
  or (_22457_, _22454_, _15624_);
  and (_22458_, _22457_, _22455_);
  nor (_22459_, _22458_, _22450_);
  and (_22460_, _22458_, _22450_);
  or (_22461_, _22460_, _22459_);
  nor (_22462_, _22461_, _07224_);
  and (_22463_, _22461_, _07224_);
  or (_22464_, _22463_, _02032_);
  or (_22465_, _22464_, _22462_);
  and (_22466_, _22465_, _02037_);
  and (_22468_, _22466_, _22440_);
  not (_22469_, _15008_);
  and (_22470_, _14069_, _13720_);
  nor (_22471_, _14069_, _13720_);
  nor (_22472_, _22471_, _22470_);
  not (_22473_, _22472_);
  not (_22474_, _14698_);
  and (_22475_, _22474_, _14372_);
  nor (_22476_, _22474_, _14372_);
  nor (_22477_, _22476_, _22475_);
  and (_22479_, _22477_, _22473_);
  nor (_22480_, _22477_, _22473_);
  or (_22481_, _22480_, _22479_);
  nor (_22482_, _22481_, _22469_);
  and (_22483_, _22481_, _22469_);
  or (_22484_, _22483_, _22482_);
  and (_22485_, _22484_, _15330_);
  nor (_22486_, _22484_, _15330_);
  or (_22487_, _22486_, _22485_);
  and (_22488_, _22487_, _15629_);
  nor (_22490_, _22487_, _15629_);
  or (_22491_, _22490_, _22488_);
  and (_22492_, _22491_, _07229_);
  nor (_22493_, _22491_, _07229_);
  or (_22494_, _22493_, _22492_);
  and (_22495_, _22494_, _01765_);
  or (_22496_, _22495_, _22468_);
  and (_22497_, _22496_, _06560_);
  and (_22498_, _06262_, _15634_);
  nor (_22499_, _06262_, _15634_);
  nor (_22501_, _22499_, _22498_);
  not (_22502_, _22501_);
  nor (_22503_, _06344_, _06295_);
  and (_22504_, _06344_, _06295_);
  nor (_22505_, _22504_, _22503_);
  not (_22506_, _22505_);
  and (_22507_, _22506_, _06398_);
  nor (_22508_, _22506_, _06398_);
  nor (_22509_, _22508_, _22507_);
  and (_22510_, _22509_, _22502_);
  nor (_22512_, _22509_, _22502_);
  nor (_22513_, _22512_, _22510_);
  nor (_22514_, _06479_, _06220_);
  and (_22515_, _06479_, _06220_);
  nor (_22516_, _22515_, _22514_);
  and (_22517_, _22516_, _22513_);
  nor (_22518_, _22516_, _22513_);
  nor (_22519_, _22518_, _22517_);
  nor (_22520_, _22519_, _13176_);
  and (_22521_, _22519_, _13176_);
  or (_22523_, _22521_, _22520_);
  and (_22524_, _22523_, _06202_);
  or (_22525_, _22524_, _22497_);
  and (_22526_, _22525_, _01776_);
  nand (_22527_, _22398_, _01775_);
  nor (_22528_, _04915_, _02124_);
  not (_22529_, _03344_);
  nor (_22530_, _10550_, _01711_);
  and (_22531_, _22530_, _22529_);
  and (_22532_, _22531_, _22528_);
  nand (_22534_, _22532_, _22527_);
  or (_22535_, _22534_, _22526_);
  or (_22536_, _22532_, _21908_);
  nand (_22537_, _22536_, _22535_);
  nor (_22538_, _02730_, _03333_);
  nor (_22539_, _22538_, _03352_);
  nand (_22540_, _22539_, _22537_);
  or (_22541_, _22539_, _21908_);
  and (_22542_, _22541_, _01995_);
  and (_22543_, _22542_, _22540_);
  nor (_22545_, _14079_, _13810_);
  and (_22546_, _14079_, _13810_);
  or (_22547_, _22546_, _22545_);
  nor (_22548_, _14708_, _14382_);
  and (_22549_, _14708_, _14382_);
  nor (_22550_, _22549_, _22548_);
  nor (_22551_, _22550_, _22547_);
  and (_22552_, _22550_, _22547_);
  or (_22553_, _22552_, _22551_);
  nor (_22554_, _15340_, _15018_);
  and (_22556_, _15340_, _15018_);
  nor (_22557_, _22556_, _22554_);
  and (_22558_, _22557_, _15641_);
  nor (_22559_, _22557_, _15641_);
  nor (_22560_, _22559_, _22558_);
  nor (_22561_, _22560_, _22553_);
  and (_22562_, _22560_, _22553_);
  nor (_22563_, _22562_, _22561_);
  and (_22564_, _22563_, _07242_);
  nor (_22565_, _22563_, _07242_);
  or (_22567_, _22565_, _22564_);
  and (_22568_, _22567_, _01994_);
  or (_22569_, _22568_, _22543_);
  and (_22570_, _22569_, _07240_);
  nand (_22571_, _22398_, _07239_);
  and (_22572_, _10600_, _10150_);
  nand (_22573_, _22572_, _22571_);
  or (_22574_, _22573_, _22570_);
  or (_22575_, _22572_, _21908_);
  and (_22576_, _22575_, _10605_);
  and (_22578_, _22576_, _22574_);
  nand (_22579_, _21908_, _10604_);
  nand (_22580_, _22579_, _10146_);
  or (_22581_, _22580_, _22578_);
  nor (_22582_, _14534_, _06632_);
  and (_22583_, _14534_, _06632_);
  nor (_22584_, _22583_, _22582_);
  and (_22585_, _13818_, _06636_);
  nor (_22586_, _22585_, _14302_);
  nor (_22587_, _22586_, _22584_);
  and (_22589_, _22586_, _22584_);
  nor (_22590_, _22589_, _22587_);
  nor (_22591_, _15170_, _06625_);
  and (_22592_, _15170_, _06625_);
  nor (_22593_, _22592_, _22591_);
  nor (_22594_, _22593_, _22590_);
  and (_22595_, _22593_, _22590_);
  nor (_22596_, _22595_, _22594_);
  nand (_22597_, _06620_, _06617_);
  or (_22598_, _06620_, _06617_);
  and (_22600_, _22598_, _22597_);
  nand (_22601_, _22600_, _22596_);
  or (_22602_, _22600_, _22596_);
  and (_22603_, _22602_, _22601_);
  or (_22604_, _22603_, _10146_);
  and (_22605_, _22604_, _22581_);
  or (_22606_, _22605_, _07263_);
  nor (_22607_, _14563_, _07463_);
  and (_22608_, _14563_, _07463_);
  nor (_22609_, _22608_, _22607_);
  and (_22611_, _13827_, _07467_);
  nor (_22612_, _22611_, _14321_);
  nor (_22613_, _22612_, _22609_);
  and (_22614_, _22612_, _22609_);
  nor (_22615_, _22614_, _22613_);
  nor (_22616_, _15193_, _07456_);
  and (_22617_, _15193_, _07456_);
  nor (_22618_, _22617_, _22616_);
  nor (_22619_, _22618_, _22615_);
  and (_22620_, _22618_, _22615_);
  nor (_22622_, _22620_, _22619_);
  nor (_22623_, _22622_, _07451_);
  and (_22624_, _22622_, _07451_);
  or (_22625_, _22624_, _22623_);
  nor (_22626_, _22625_, _07271_);
  and (_22627_, _22625_, _07271_);
  or (_22628_, _22627_, _22626_);
  or (_22629_, _22628_, _07264_);
  and (_22630_, _22629_, _02330_);
  and (_22631_, _22630_, _22606_);
  nor (_22633_, _11511_, _11315_);
  and (_22634_, _11511_, _11315_);
  nor (_22635_, _22634_, _22633_);
  and (_22636_, _11113_, _10792_);
  nor (_22637_, _11113_, _10792_);
  or (_22638_, _22637_, _22636_);
  and (_22639_, _22638_, _22635_);
  nor (_22640_, _22638_, _22635_);
  nor (_22641_, _22640_, _22639_);
  or (_22642_, _22641_, _11588_);
  nand (_22644_, _22641_, _11588_);
  and (_22645_, _22644_, _22642_);
  nor (_22646_, _22645_, _11786_);
  and (_22647_, _22645_, _11786_);
  or (_22648_, _22647_, _22646_);
  nor (_22649_, _22648_, _12118_);
  and (_22650_, _22648_, _12118_);
  nor (_22651_, _22650_, _22649_);
  not (_22652_, _22651_);
  nor (_22653_, _22652_, _04942_);
  and (_22655_, _22652_, _04942_);
  or (_22656_, _22655_, _22653_);
  and (_22657_, _22656_, _02329_);
  or (_22658_, _22657_, _06734_);
  or (_22659_, _22658_, _22631_);
  nor (_22660_, _08898_, _08883_);
  and (_22661_, _08898_, _08883_);
  nor (_22662_, _22661_, _22660_);
  and (_22663_, _08919_, _07552_);
  nor (_22664_, _22663_, _08920_);
  and (_22666_, _22664_, _07549_);
  nor (_22667_, _22664_, _07549_);
  nor (_22668_, _22667_, _22666_);
  nor (_22669_, _22668_, _22662_);
  and (_22670_, _22668_, _22662_);
  nor (_22671_, _22670_, _22669_);
  nand (_22672_, _22671_, _07540_);
  or (_22673_, _22671_, _07540_);
  and (_22674_, _22673_, _22672_);
  or (_22675_, _22674_, _07537_);
  nand (_22677_, _22674_, _07537_);
  and (_22678_, _22677_, _22675_);
  nor (_22679_, _22678_, _07280_);
  and (_22680_, _22678_, _07280_);
  or (_22681_, _22680_, _07281_);
  or (_22682_, _22681_, _22679_);
  and (_22683_, _22682_, _03059_);
  and (_22684_, _22683_, _22659_);
  not (_22685_, _15679_);
  and (_22686_, _13953_, _13716_);
  nor (_22688_, _13953_, _13716_);
  nor (_22689_, _22688_, _22686_);
  not (_22690_, _14545_);
  and (_22691_, _22690_, _14225_);
  nor (_22692_, _22690_, _14225_);
  nor (_22693_, _22692_, _22691_);
  nor (_22694_, _22693_, _22689_);
  and (_22695_, _22693_, _22689_);
  or (_22696_, _22695_, _22694_);
  not (_22697_, _15184_);
  and (_22699_, _22697_, _15048_);
  nor (_22700_, _22697_, _15048_);
  nor (_22701_, _22700_, _22699_);
  and (_22702_, _22701_, _22696_);
  nor (_22703_, _22701_, _22696_);
  nor (_22704_, _22703_, _22702_);
  nor (_22705_, _22704_, _22685_);
  and (_22706_, _22704_, _22685_);
  or (_22707_, _22706_, _22705_);
  and (_22708_, _22707_, _07286_);
  nor (_22710_, _22707_, _07286_);
  or (_22711_, _22710_, _22708_);
  and (_22712_, _22711_, _02210_);
  or (_22713_, _22712_, _22684_);
  and (_22714_, _22713_, _03061_);
  not (_22715_, _21931_);
  nand (_22716_, _21908_, _02331_);
  nor (_22717_, _22716_, _03841_);
  or (_22718_, _22717_, _22715_);
  or (_22719_, _22718_, _22714_);
  nand (_22721_, _22719_, _21932_);
  nand (_22722_, _22721_, _10138_);
  or (_22723_, _06637_, _06634_);
  nand (_22724_, _06637_, _06634_);
  and (_22725_, _22724_, _22723_);
  and (_22726_, _06628_, _06630_);
  nor (_22727_, _06628_, _06630_);
  nor (_22728_, _22727_, _22726_);
  and (_22729_, _22728_, _22725_);
  nor (_22730_, _22728_, _22725_);
  nor (_22732_, _22730_, _22729_);
  not (_22733_, _06621_);
  nor (_22734_, _06623_, _06618_);
  and (_22735_, _06623_, _06618_);
  nor (_22736_, _22735_, _22734_);
  nor (_22737_, _22736_, _22733_);
  and (_22738_, _22736_, _22733_);
  nor (_22739_, _22738_, _22737_);
  and (_22740_, _22739_, _22732_);
  nor (_22741_, _22739_, _22732_);
  or (_22743_, _22741_, _22740_);
  and (_22744_, _22743_, _06616_);
  nor (_22745_, _22743_, _06616_);
  or (_22746_, _22745_, _22744_);
  or (_22747_, _22746_, _10138_);
  and (_22748_, _22747_, _02703_);
  and (_22749_, _22748_, _22722_);
  and (_22750_, _22746_, _02702_);
  or (_22751_, _22750_, _07304_);
  or (_22752_, _22751_, _22749_);
  or (_22754_, _07468_, _07465_);
  nand (_22755_, _07468_, _07465_);
  and (_22756_, _22755_, _22754_);
  not (_22757_, _22756_);
  and (_22758_, _07460_, _07461_);
  nor (_22759_, _07460_, _07461_);
  nor (_22760_, _22759_, _22758_);
  nor (_22761_, _22760_, _22757_);
  and (_22762_, _22760_, _22757_);
  nor (_22763_, _22762_, _22761_);
  nor (_22765_, _07452_, _07454_);
  and (_22766_, _07452_, _07454_);
  nor (_22767_, _22766_, _22765_);
  nor (_22768_, _22767_, _07449_);
  and (_22769_, _22767_, _07449_);
  nor (_22770_, _22769_, _22768_);
  not (_22771_, _22770_);
  and (_22772_, _22771_, _22763_);
  nor (_22773_, _22771_, _22763_);
  nor (_22774_, _22773_, _22772_);
  nor (_22776_, _22774_, _07270_);
  and (_22777_, _22774_, _07270_);
  or (_22778_, _22777_, _22776_);
  or (_22779_, _22778_, _07305_);
  and (_22780_, _22779_, _02341_);
  and (_22781_, _22780_, _22752_);
  nor (_22782_, _11111_, _10791_);
  and (_22783_, _11111_, _10791_);
  nor (_22784_, _22783_, _22782_);
  not (_22785_, _22784_);
  not (_22787_, _11509_);
  and (_22788_, _22787_, _11313_);
  nor (_22789_, _22787_, _11313_);
  nor (_22790_, _22789_, _22788_);
  nor (_22791_, _22790_, _22785_);
  and (_22792_, _22790_, _22785_);
  nor (_22793_, _22792_, _22791_);
  not (_22794_, _12116_);
  nor (_22795_, _11784_, _11586_);
  and (_22796_, _11784_, _11586_);
  nor (_22798_, _22796_, _22795_);
  nor (_22799_, _22798_, _22794_);
  and (_22800_, _22798_, _22794_);
  nor (_22801_, _22800_, _22799_);
  not (_22802_, _22801_);
  nor (_22803_, _22802_, _22793_);
  and (_22804_, _22802_, _22793_);
  nor (_22805_, _22804_, _22803_);
  not (_22806_, _22805_);
  nor (_22807_, _22806_, _04941_);
  and (_22809_, _22806_, _04941_);
  or (_22810_, _22809_, _22807_);
  and (_22811_, _22810_, _02340_);
  or (_22812_, _22811_, _07312_);
  or (_22813_, _22812_, _22781_);
  not (_22814_, _07541_);
  or (_22815_, _07553_, _07550_);
  nand (_22816_, _07553_, _07550_);
  and (_22817_, _22816_, _22815_);
  not (_22818_, _07544_);
  and (_22820_, _22818_, _07546_);
  nor (_22821_, _22818_, _07546_);
  nor (_22822_, _22821_, _22820_);
  not (_22823_, _22822_);
  and (_22824_, _22823_, _22817_);
  nor (_22825_, _22823_, _22817_);
  nor (_22826_, _22825_, _22824_);
  nand (_22827_, _22826_, _22814_);
  or (_22828_, _22826_, _22814_);
  and (_22829_, _22828_, _22827_);
  or (_22831_, _22829_, _07538_);
  nand (_22832_, _22829_, _07538_);
  and (_22833_, _22832_, _22831_);
  or (_22834_, _22833_, _07535_);
  nand (_22835_, _22833_, _07535_);
  and (_22836_, _22835_, _22834_);
  and (_22837_, _22836_, _07279_);
  nor (_22838_, _22836_, _07279_);
  or (_22839_, _22838_, _22837_);
  or (_22840_, _22839_, _07313_);
  and (_22842_, _22840_, _02208_);
  and (_22843_, _22842_, _22813_);
  and (_22844_, _10650_, _09561_);
  nor (_22845_, _14431_, _13854_);
  and (_22846_, _14431_, _13854_);
  nor (_22847_, _22846_, _22845_);
  nor (_22848_, _15704_, _15069_);
  and (_22849_, _15704_, _15069_);
  nor (_22850_, _22849_, _22848_);
  and (_22851_, _22850_, _22847_);
  nor (_22853_, _22850_, _22847_);
  nor (_22854_, _22853_, _22851_);
  nor (_22855_, _15396_, _14757_);
  and (_22856_, _15396_, _14757_);
  nor (_22857_, _22856_, _22855_);
  nor (_22858_, _14123_, _07320_);
  and (_22859_, _14123_, _07320_);
  nor (_22860_, _22859_, _22858_);
  and (_22861_, _22860_, _22857_);
  nor (_22862_, _22860_, _22857_);
  nor (_22864_, _22862_, _22861_);
  not (_22865_, _22864_);
  nand (_22866_, _22865_, _22854_);
  or (_22867_, _22865_, _22854_);
  and (_22868_, _22867_, _02206_);
  nand (_22869_, _22868_, _22866_);
  nand (_22870_, _22869_, _22844_);
  or (_22871_, _22870_, _22843_);
  or (_22872_, _21908_, _22844_);
  and (_22873_, _22872_, _22871_);
  or (_22874_, _22873_, _10654_);
  nor (_22875_, _13826_, _07466_);
  and (_22876_, _13826_, _07466_);
  nor (_22877_, _22876_, _22875_);
  not (_22878_, _22877_);
  and (_22879_, _07458_, _07462_);
  nor (_22880_, _07458_, _07462_);
  nor (_22881_, _22880_, _22879_);
  nor (_22882_, _22881_, _22878_);
  and (_22883_, _22881_, _22878_);
  nor (_22885_, _22883_, _22882_);
  not (_22886_, _07453_);
  nor (_22887_, _07455_, _07450_);
  and (_22888_, _07455_, _07450_);
  nor (_22889_, _22888_, _22887_);
  nor (_22890_, _22889_, _22886_);
  and (_22891_, _22889_, _22886_);
  nor (_22892_, _22891_, _22890_);
  nor (_22893_, _22892_, _22885_);
  and (_22894_, _22892_, _22885_);
  nor (_22896_, _22894_, _22893_);
  nor (_22897_, _22896_, _07269_);
  and (_22898_, _22896_, _07269_);
  or (_22899_, _22898_, _22897_);
  or (_22900_, _22899_, _10127_);
  nor (_22901_, _13817_, _06635_);
  and (_22902_, _13817_, _06635_);
  nor (_22903_, _22902_, _22901_);
  and (_22904_, _22903_, _06631_);
  nor (_22905_, _22903_, _06631_);
  or (_22907_, _22905_, _22904_);
  and (_22908_, _22907_, _06629_);
  nor (_22909_, _22907_, _06629_);
  or (_22910_, _22909_, _22908_);
  not (_22911_, _06622_);
  nor (_22912_, _06624_, _06619_);
  and (_22913_, _06624_, _06619_);
  nor (_22914_, _22913_, _22912_);
  nor (_22915_, _22914_, _22911_);
  and (_22916_, _22914_, _22911_);
  nor (_22918_, _22916_, _22915_);
  nor (_22919_, _22918_, _22910_);
  and (_22920_, _22918_, _22910_);
  nor (_22921_, _22920_, _22919_);
  nor (_22922_, _22921_, _06615_);
  and (_22923_, _22921_, _06615_);
  or (_22924_, _22923_, _22922_);
  or (_22925_, _22924_, _10132_);
  and (_22926_, _22925_, _02337_);
  and (_22927_, _22926_, _22900_);
  and (_22929_, _22927_, _22874_);
  nor (_22930_, _11112_, _10789_);
  and (_22931_, _11112_, _10789_);
  nor (_22932_, _22931_, _22930_);
  and (_22933_, _22932_, _11314_);
  nor (_22934_, _22932_, _11314_);
  or (_22935_, _22934_, _22933_);
  nand (_22936_, _22935_, _11510_);
  or (_22937_, _22935_, _11510_);
  and (_22938_, _22937_, _22936_);
  nor (_22940_, _11785_, _11587_);
  and (_22941_, _11785_, _11587_);
  nor (_22942_, _22941_, _22940_);
  nor (_22943_, _22942_, _12117_);
  and (_22944_, _22942_, _12117_);
  nor (_22945_, _22944_, _22943_);
  and (_22946_, _22945_, _22938_);
  nor (_22947_, _22945_, _22938_);
  nor (_22948_, _22947_, _22946_);
  and (_22949_, _22948_, _04940_);
  nor (_22951_, _22948_, _04940_);
  or (_22952_, _22951_, _22949_);
  and (_22953_, _22952_, _02336_);
  or (_22954_, _22953_, _07338_);
  or (_22955_, _22954_, _22929_);
  nor (_22956_, _08918_, _07551_);
  and (_22957_, _08918_, _07551_);
  nor (_22958_, _22957_, _22956_);
  not (_22959_, _22958_);
  not (_22960_, _07545_);
  and (_22962_, _22960_, _07547_);
  nor (_22963_, _22960_, _07547_);
  nor (_22964_, _22963_, _22962_);
  nor (_22965_, _22964_, _22959_);
  and (_22966_, _22964_, _22959_);
  nor (_22967_, _22966_, _22965_);
  and (_22968_, _22967_, _07542_);
  nor (_22969_, _22967_, _07542_);
  or (_22970_, _22969_, _22968_);
  and (_22971_, _22970_, _07539_);
  nor (_22973_, _22970_, _07539_);
  or (_22974_, _22973_, _22971_);
  and (_22975_, _22974_, _07536_);
  nor (_22976_, _22974_, _07536_);
  or (_22977_, _22976_, _22975_);
  and (_22978_, _22977_, _07278_);
  nor (_22979_, _22977_, _07278_);
  or (_22980_, _22979_, _22978_);
  or (_22981_, _22980_, _07341_);
  and (_22982_, _22981_, _04953_);
  and (_22984_, _22982_, _22955_);
  and (_22985_, _10124_, _10123_);
  nor (_22986_, _14144_, _13880_);
  and (_22987_, _14144_, _13880_);
  or (_22988_, _22987_, _22986_);
  nor (_22989_, _14541_, _14452_);
  and (_22990_, _14541_, _14452_);
  nor (_22991_, _22990_, _22989_);
  nor (_22992_, _22991_, _22988_);
  and (_22993_, _22991_, _22988_);
  nor (_22995_, _22993_, _22992_);
  not (_22996_, _22995_);
  nor (_22997_, _15727_, _15412_);
  and (_22998_, _15727_, _15412_);
  nor (_22999_, _22998_, _22997_);
  not (_23000_, _15090_);
  and (_23001_, _23000_, _07350_);
  nor (_23002_, _23000_, _07350_);
  nor (_23003_, _23002_, _23001_);
  nor (_23004_, _23003_, _22999_);
  and (_23006_, _23003_, _22999_);
  nor (_23007_, _23006_, _23004_);
  nand (_23008_, _23007_, _22996_);
  or (_23009_, _23007_, _22996_);
  and (_23010_, _23009_, _02202_);
  nand (_23011_, _23010_, _23008_);
  nand (_23012_, _23011_, _22985_);
  or (_23013_, _23012_, _22984_);
  or (_23014_, _21908_, _22985_);
  nand (_23015_, _23014_, _23013_);
  nand (_23017_, _23015_, _06729_);
  not (_23018_, _15177_);
  not (_23019_, _14781_);
  nor (_23020_, _06924_, _06706_);
  nor (_23021_, _14149_, _22276_);
  nor (_23022_, _23021_, _23020_);
  nor (_23023_, _23022_, _14457_);
  and (_23024_, _23022_, _14457_);
  nor (_23025_, _23024_, _23023_);
  and (_23026_, _23025_, _23019_);
  nor (_23028_, _23025_, _23019_);
  nor (_23029_, _23028_, _23026_);
  nor (_23030_, _23029_, _15095_);
  and (_23031_, _23029_, _15095_);
  or (_23032_, _23031_, _23030_);
  nor (_23033_, _23032_, _23018_);
  and (_23034_, _23032_, _23018_);
  nor (_23035_, _23034_, _23033_);
  nor (_23036_, _23035_, _15733_);
  and (_23037_, _23035_, _15733_);
  or (_23039_, _23037_, _23036_);
  nand (_23040_, _23039_, _06726_);
  or (_23041_, _23039_, _06726_);
  and (_23042_, _23041_, _23040_);
  and (_23043_, _23042_, _06728_);
  or (_23044_, _23043_, _06730_);
  and (_23045_, _23044_, _23017_);
  and (_23046_, _23042_, _06727_);
  or (_23047_, _23046_, _06654_);
  or (_23048_, _23047_, _23045_);
  not (_23050_, _07380_);
  nor (_23051_, _07002_, _07000_);
  nor (_23052_, _14154_, _22303_);
  nor (_23053_, _23052_, _23051_);
  nor (_23054_, _23053_, _14462_);
  and (_23055_, _23053_, _14462_);
  nor (_23056_, _23055_, _23054_);
  and (_23057_, _23056_, _14786_);
  nor (_23058_, _23056_, _14786_);
  or (_23059_, _23058_, _23057_);
  nor (_23061_, _23059_, _15100_);
  and (_23062_, _23059_, _15100_);
  or (_23063_, _23062_, _23061_);
  nor (_23064_, _23063_, _15419_);
  and (_23065_, _23063_, _15419_);
  or (_23066_, _23065_, _23064_);
  and (_23067_, _23066_, _15738_);
  nor (_23068_, _23066_, _15738_);
  or (_23069_, _23068_, _23067_);
  nor (_23070_, _23069_, _23050_);
  and (_23072_, _23069_, _23050_);
  or (_23073_, _23072_, _07356_);
  or (_23074_, _23073_, _23070_);
  and (_23075_, _23074_, _02346_);
  and (_23076_, _23075_, _23048_);
  not (_23077_, _07411_);
  and (_23078_, _14159_, _07186_);
  nor (_23079_, _14159_, _07186_);
  nor (_23080_, _23079_, _23078_);
  nor (_23081_, _23080_, _14467_);
  and (_23083_, _23080_, _14467_);
  nor (_23084_, _23083_, _23081_);
  and (_23085_, _23084_, _14791_);
  nor (_23086_, _23084_, _14791_);
  or (_23087_, _23086_, _23085_);
  nor (_23088_, _23087_, _15105_);
  and (_23089_, _23087_, _15105_);
  or (_23090_, _23089_, _23088_);
  nor (_23091_, _23090_, _15424_);
  and (_23092_, _23090_, _15424_);
  or (_23094_, _23092_, _23091_);
  and (_23095_, _23094_, _15744_);
  nor (_23096_, _23094_, _15744_);
  or (_23097_, _23096_, _23095_);
  nand (_23098_, _23097_, _23077_);
  or (_23099_, _23097_, _23077_);
  and (_23100_, _23099_, _02345_);
  and (_23101_, _23100_, _23098_);
  or (_23102_, _23101_, _07384_);
  or (_23103_, _23102_, _23076_);
  not (_23105_, _07439_);
  not (_23106_, _15429_);
  nor (_23107_, _13945_, _22355_);
  nor (_23108_, _06792_, _06786_);
  nor (_23109_, _23108_, _23107_);
  nor (_23110_, _23109_, _14472_);
  and (_23111_, _23109_, _14472_);
  nor (_23112_, _23111_, _23110_);
  nor (_23113_, _23112_, _14796_);
  and (_23114_, _23112_, _14796_);
  or (_23116_, _23114_, _23113_);
  and (_23117_, _23116_, _15110_);
  nor (_23118_, _23116_, _15110_);
  or (_23119_, _23118_, _23117_);
  and (_23120_, _23119_, _23106_);
  nor (_23121_, _23119_, _23106_);
  nor (_23122_, _23121_, _23120_);
  nor (_23123_, _23122_, _15749_);
  and (_23124_, _23122_, _15749_);
  or (_23125_, _23124_, _23123_);
  nor (_23127_, _23125_, _23105_);
  and (_23128_, _23125_, _23105_);
  or (_23129_, _23128_, _07417_);
  or (_23130_, _23129_, _23127_);
  and (_23131_, _23130_, _07416_);
  and (_23132_, _23131_, _23103_);
  nor (_23133_, _07191_, _07190_);
  nor (_23134_, _14235_, \oc8051_golden_model_1.ACC [3]);
  and (_23135_, _14235_, \oc8051_golden_model_1.ACC [3]);
  nor (_23136_, _23135_, _23134_);
  and (_23138_, _23136_, _22064_);
  nor (_23139_, _23136_, _22064_);
  nor (_23140_, _23139_, _23138_);
  not (_23141_, _23140_);
  nand (_23142_, _23141_, _23133_);
  or (_23143_, _23141_, _23133_);
  and (_23144_, _23143_, _23142_);
  nand (_23145_, _23144_, _07415_);
  nor (_23146_, _02350_, _01726_);
  and (_23147_, _23146_, _10689_);
  nand (_23149_, _23147_, _23145_);
  or (_23150_, _23149_, _23132_);
  or (_23151_, _23147_, _21908_);
  and (_23152_, _23151_, _06614_);
  and (_23153_, _23152_, _23150_);
  nor (_23154_, _13817_, _06636_);
  and (_23155_, _13817_, _06636_);
  nor (_23156_, _23155_, _23154_);
  and (_23157_, _23156_, _14217_);
  nor (_23158_, _23156_, _14217_);
  nor (_23160_, _23158_, _23157_);
  and (_23161_, _23160_, _14537_);
  nor (_23162_, _23160_, _14537_);
  nor (_23163_, _23162_, _23161_);
  nor (_23164_, _23163_, _15118_);
  and (_23165_, _23163_, _15118_);
  or (_23166_, _23165_, _23164_);
  nor (_23167_, _23166_, _15174_);
  and (_23168_, _23166_, _15174_);
  nor (_23169_, _23168_, _23167_);
  nor (_23171_, _23169_, _15758_);
  and (_23172_, _23169_, _15758_);
  or (_23173_, _23172_, _23171_);
  or (_23174_, _23173_, _06652_);
  nand (_23175_, _23173_, _06652_);
  and (_23176_, _23175_, _09155_);
  and (_23177_, _23176_, _23174_);
  or (_23178_, _23177_, _06609_);
  or (_23179_, _23178_, _23153_);
  nor (_23180_, _13826_, _07467_);
  and (_23182_, _13826_, _07467_);
  nor (_23183_, _23182_, _23180_);
  and (_23184_, _23183_, _14486_);
  nor (_23185_, _23183_, _14486_);
  nor (_23186_, _23185_, _23184_);
  and (_23187_, _23186_, _14807_);
  nor (_23188_, _23186_, _14807_);
  nor (_23189_, _23188_, _23187_);
  nor (_23190_, _23189_, _15123_);
  and (_23191_, _23189_, _15123_);
  or (_23193_, _23191_, _23190_);
  and (_23194_, _23193_, _15441_);
  nor (_23195_, _23193_, _15441_);
  nor (_23196_, _23195_, _23194_);
  and (_23197_, _23196_, _15764_);
  nor (_23198_, _23196_, _15764_);
  nor (_23199_, _23198_, _23197_);
  and (_23200_, _23199_, _07483_);
  nor (_23201_, _23199_, _07483_);
  or (_23202_, _23201_, _23200_);
  or (_23204_, _23202_, _07448_);
  and (_23205_, _23204_, _07488_);
  and (_23206_, _23205_, _23179_);
  nor (_23207_, _14179_, _08874_);
  and (_23208_, _14179_, _08874_);
  or (_23209_, _23208_, _23207_);
  nor (_23210_, _23209_, _14491_);
  and (_23211_, _23209_, _14491_);
  nor (_23212_, _23211_, _23210_);
  and (_23213_, _23212_, _14813_);
  nor (_23215_, _23212_, _14813_);
  nor (_23216_, _23215_, _23213_);
  and (_23217_, _23216_, _15128_);
  nor (_23218_, _23216_, _15128_);
  nor (_23219_, _23218_, _23217_);
  nor (_23220_, _23219_, _15446_);
  and (_23221_, _23219_, _15446_);
  or (_23222_, _23221_, _23220_);
  nor (_23223_, _23222_, _15769_);
  and (_23224_, _23222_, _15769_);
  or (_23226_, _23224_, _23223_);
  not (_23227_, _23226_);
  nor (_23228_, _23227_, _07529_);
  and (_23229_, _23227_, _07529_);
  or (_23230_, _23229_, _23228_);
  and (_23231_, _23230_, _02085_);
  nor (_23232_, _14184_, _08919_);
  nor (_23233_, _23232_, _22663_);
  nor (_23234_, _23233_, _14496_);
  and (_23235_, _23233_, _14496_);
  or (_23237_, _23235_, _23234_);
  nor (_23238_, _23237_, _14819_);
  and (_23239_, _23237_, _14819_);
  nor (_23240_, _23239_, _23238_);
  nor (_23241_, _23240_, _15133_);
  and (_23242_, _23240_, _15133_);
  or (_23243_, _23242_, _23241_);
  nor (_23244_, _23243_, _15451_);
  and (_23245_, _23243_, _15451_);
  or (_23246_, _23245_, _23244_);
  nor (_23248_, _23246_, _15775_);
  and (_23249_, _23246_, _15775_);
  or (_23250_, _23249_, _23248_);
  or (_23251_, _23250_, _07568_);
  nand (_23252_, _23250_, _07568_);
  and (_23253_, _23252_, _07487_);
  nand (_23254_, _23253_, _23251_);
  nor (_23255_, _13706_, _04969_);
  not (_23256_, _23255_);
  or (_23257_, _03274_, _02765_);
  not (_23259_, _23257_);
  and (_23260_, _02247_, _01566_);
  nor (_23261_, _23260_, _02243_);
  and (_23262_, _23261_, _23259_);
  and (_23263_, _01737_, _01695_);
  and (_23264_, _23263_, _05332_);
  not (_23265_, _23264_);
  nor (_23266_, _03084_, _03350_);
  and (_23267_, _23266_, _23265_);
  and (_23268_, _23267_, _23262_);
  and (_23270_, _23268_, _23256_);
  nand (_23271_, _23270_, _23254_);
  or (_23272_, _23271_, _23231_);
  or (_23273_, _23272_, _23206_);
  or (_23274_, _23270_, _21908_);
  and (_23275_, _23274_, _02778_);
  and (_23276_, _23275_, _23273_);
  and (_23277_, _22099_, _02366_);
  or (_23278_, _23277_, _07575_);
  or (_23279_, _23278_, _23276_);
  and (_23281_, _23279_, _21930_);
  and (_23282_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_23283_, _23282_, _06839_);
  or (_23284_, _23140_, _23283_);
  nand (_23285_, _23140_, _23283_);
  and (_23286_, _23285_, _23284_);
  nand (_23287_, _23286_, _07580_);
  nand (_23288_, _23287_, _01990_);
  or (_23289_, _23288_, _23281_);
  or (_23290_, _21908_, _01990_);
  and (_23292_, _23290_, _01698_);
  and (_23293_, _23292_, _23289_);
  and (_23294_, _21958_, _01697_);
  or (_23295_, _23294_, _05338_);
  or (_23296_, _23295_, _23293_);
  nand (_23297_, _23296_, _21909_);
  and (_23298_, _03292_, _05363_);
  nand (_23299_, _23298_, _23297_);
  or (_23300_, _23298_, _21908_);
  and (_23301_, _23300_, _02082_);
  and (_23303_, _23301_, _23299_);
  nor (_23304_, _14204_, _13743_);
  and (_23305_, _14204_, _13743_);
  nor (_23306_, _23305_, _23304_);
  and (_23307_, _23306_, _14519_);
  nor (_23308_, _23306_, _14519_);
  or (_23309_, _23308_, _23307_);
  and (_23310_, _23309_, _14841_);
  nor (_23311_, _23309_, _14841_);
  or (_23312_, _23311_, _23310_);
  and (_23314_, _23312_, _15156_);
  nor (_23315_, _23312_, _15156_);
  or (_23316_, _23315_, _23314_);
  and (_23317_, _23316_, _15473_);
  nor (_23318_, _23316_, _15473_);
  or (_23319_, _23318_, _23317_);
  and (_23320_, _23319_, _15799_);
  nor (_23321_, _23319_, _15799_);
  or (_23322_, _23321_, _23320_);
  and (_23323_, _23322_, _07602_);
  nor (_23325_, _23322_, _07602_);
  or (_23326_, _23325_, _23323_);
  and (_23327_, _23326_, _02081_);
  or (_23328_, _23327_, _23303_);
  and (_23329_, _23328_, _07600_);
  nor (_23330_, _02198_, _01732_);
  nor (_23331_, _10762_, _07606_);
  and (_23332_, _23331_, _23330_);
  not (_23333_, _07607_);
  and (_23334_, _14235_, _23333_);
  and (_23336_, _23334_, _06377_);
  nor (_23337_, _23334_, _06377_);
  nor (_23338_, _23337_, _23336_);
  nor (_23339_, _23338_, _15161_);
  and (_23340_, _23338_, _15161_);
  or (_23341_, _23340_, _23339_);
  and (_23342_, _23341_, _15804_);
  nor (_23343_, _23341_, _15804_);
  nor (_23344_, _23343_, _23342_);
  nor (_23345_, _15478_, _07614_);
  and (_23347_, _15478_, _07614_);
  nor (_23348_, _23347_, _23345_);
  not (_23349_, _23348_);
  nand (_23350_, _23349_, _23344_);
  or (_23351_, _23349_, _23344_);
  and (_23352_, _23351_, _07599_);
  nand (_23353_, _23352_, _23350_);
  nand (_23354_, _23353_, _23332_);
  or (_23355_, _23354_, _23329_);
  or (_23356_, _23332_, _21908_);
  and (_23358_, _23356_, _39632_);
  and (_23359_, _23358_, _23355_);
  or (_23360_, _23359_, _21892_);
  and (_41701_, _23360_, _39026_);
  not (_23361_, \oc8051_golden_model_1.PSW [1]);
  nor (_23362_, _03838_, _23361_);
  nor (_23363_, _08489_, _03161_);
  or (_23364_, _23363_, _23362_);
  or (_23365_, _23364_, _02519_);
  or (_23366_, _03838_, \oc8051_golden_model_1.PSW [1]);
  and (_23368_, _11001_, _03838_);
  not (_23369_, _23368_);
  and (_23370_, _23369_, _23366_);
  or (_23371_, _23370_, _03006_);
  nand (_23372_, _03838_, _01804_);
  and (_23373_, _23372_, _23366_);
  and (_23374_, _23373_, _02062_);
  nor (_23375_, _02062_, _23361_);
  or (_23376_, _23375_, _02158_);
  or (_23377_, _23376_, _23374_);
  and (_23379_, _23377_, _02058_);
  and (_23380_, _23379_, _23371_);
  nor (_23381_, _04476_, _23361_);
  and (_23382_, _11005_, _04476_);
  or (_23383_, _23382_, _23381_);
  and (_23384_, _23383_, _02057_);
  or (_23385_, _23384_, _02155_);
  or (_23386_, _23385_, _23380_);
  and (_23387_, _23386_, _23365_);
  or (_23388_, _23387_, _02153_);
  or (_23390_, _23373_, _02549_);
  and (_23391_, _23390_, _02054_);
  and (_23392_, _23391_, _23388_);
  and (_23393_, _10992_, _04476_);
  or (_23394_, _23393_, _23381_);
  and (_23395_, _23394_, _02053_);
  or (_23396_, _23395_, _23392_);
  or (_23397_, _23396_, _02046_);
  or (_23398_, _23381_, _11020_);
  and (_23399_, _23398_, _23383_);
  or (_23400_, _23399_, _02047_);
  and (_23401_, _23400_, _02043_);
  and (_23402_, _23401_, _23397_);
  not (_23403_, _04476_);
  nor (_23404_, _11038_, _23403_);
  or (_23405_, _23404_, _23381_);
  and (_23406_, _23405_, _02042_);
  or (_23407_, _23406_, _06188_);
  or (_23408_, _23407_, _23402_);
  or (_23409_, _23364_, _05444_);
  and (_23411_, _23409_, _23408_);
  or (_23412_, _23411_, _02031_);
  and (_23413_, _05075_, _03838_);
  or (_23414_, _23362_, _02032_);
  or (_23415_, _23414_, _23413_);
  and (_23416_, _23415_, _02037_);
  and (_23417_, _23416_, _23412_);
  nor (_23418_, _11096_, _08489_);
  or (_23419_, _23418_, _23362_);
  and (_23420_, _23419_, _01765_);
  or (_23422_, _23420_, _23417_);
  and (_23423_, _23422_, _02212_);
  or (_23424_, _10989_, _08489_);
  and (_23425_, _23424_, _02210_);
  nand (_23426_, _03838_, _02893_);
  and (_23427_, _23426_, _01994_);
  or (_23428_, _23427_, _23425_);
  and (_23429_, _23428_, _23366_);
  or (_23430_, _23429_, _23423_);
  and (_23431_, _23430_, _03061_);
  or (_23433_, _11113_, _08489_);
  and (_23434_, _23366_, _02331_);
  and (_23435_, _23434_, _23433_);
  or (_23436_, _23435_, _23431_);
  and (_23437_, _23436_, _02208_);
  or (_23438_, _10988_, _08489_);
  and (_23439_, _23366_, _02206_);
  and (_23440_, _23439_, _23438_);
  or (_23441_, _23440_, _23437_);
  and (_23442_, _23441_, _03065_);
  or (_23444_, _23362_, _04209_);
  and (_23445_, _23373_, _02342_);
  and (_23446_, _23445_, _23444_);
  or (_23447_, _23446_, _23442_);
  and (_23448_, _23447_, _02335_);
  or (_23449_, _23372_, _04209_);
  and (_23450_, _23366_, _02334_);
  and (_23451_, _23450_, _23449_);
  or (_23452_, _23451_, _02366_);
  or (_23453_, _23426_, _04209_);
  and (_23455_, _23366_, _02202_);
  and (_23456_, _23455_, _23453_);
  or (_23457_, _23456_, _23452_);
  or (_23458_, _23457_, _23448_);
  or (_23459_, _23370_, _02778_);
  and (_23460_, _23459_, _01698_);
  and (_23461_, _23460_, _23458_);
  and (_23462_, _23394_, _01697_);
  or (_23463_, _23462_, _02081_);
  or (_23464_, _23463_, _23461_);
  or (_23466_, _23368_, _23362_);
  or (_23467_, _23466_, _02082_);
  and (_23468_, _23467_, _23464_);
  or (_23469_, _23468_, _39633_);
  or (_23470_, _39632_, \oc8051_golden_model_1.PSW [1]);
  and (_23471_, _23470_, _39026_);
  and (_41702_, _23471_, _23469_);
  nand (_23472_, _06649_, _08459_);
  and (_23473_, _23472_, _08461_);
  nor (_23474_, _08459_, _06657_);
  nor (_23476_, _06658_, \oc8051_golden_model_1.ACC [7]);
  nor (_23477_, _23474_, _23476_);
  and (_23478_, _23477_, _08476_);
  nor (_23479_, _23478_, _23474_);
  and (_23480_, _23479_, _06726_);
  and (_23481_, _23474_, _06723_);
  or (_23482_, _23481_, _06730_);
  or (_23483_, _23482_, _23480_);
  not (_23484_, \oc8051_golden_model_1.PSW [2]);
  nor (_23485_, _03838_, _23484_);
  nor (_23487_, _11298_, _08489_);
  or (_23488_, _23487_, _23485_);
  and (_23489_, _23488_, _01765_);
  nor (_23490_, _08489_, _03624_);
  or (_23491_, _23490_, _23485_);
  or (_23492_, _23491_, _05444_);
  nor (_23493_, _06943_, \oc8051_golden_model_1.ACC [7]);
  nor (_23494_, _06942_, _09162_);
  nor (_23495_, _23494_, _23493_);
  and (_23496_, _23495_, _08502_);
  nor (_23497_, _23495_, _08502_);
  or (_23498_, _23497_, _23496_);
  and (_23499_, _23498_, _07012_);
  nor (_23500_, _23498_, _07012_);
  or (_23501_, _23500_, _06941_);
  or (_23502_, _23501_, _23499_);
  nor (_23503_, _23477_, _06663_);
  nor (_23504_, _09050_, _06659_);
  or (_23505_, _23504_, _23503_);
  or (_23506_, _23505_, _06934_);
  nand (_23508_, _23505_, _06934_);
  and (_23509_, _23508_, _23506_);
  and (_23510_, _23509_, _06817_);
  nor (_23511_, _04476_, _23484_);
  and (_23512_, _11192_, _04476_);
  or (_23513_, _23512_, _23511_);
  and (_23514_, _23513_, _02053_);
  nor (_23515_, _11199_, _08489_);
  or (_23516_, _23515_, _23485_);
  and (_23517_, _23516_, _02158_);
  nor (_23519_, _02062_, _23484_);
  and (_23520_, _03838_, \oc8051_golden_model_1.ACC [2]);
  or (_23521_, _23520_, _23485_);
  and (_23522_, _23521_, _02062_);
  or (_23523_, _23522_, _23519_);
  and (_23524_, _23523_, _03006_);
  or (_23525_, _23524_, _02057_);
  or (_23526_, _23525_, _23517_);
  and (_23527_, _11194_, _04476_);
  or (_23528_, _23527_, _23511_);
  or (_23530_, _23528_, _02058_);
  and (_23531_, _23530_, _02519_);
  and (_23532_, _23531_, _23526_);
  and (_23533_, _23491_, _02155_);
  or (_23534_, _23533_, _02153_);
  or (_23535_, _23534_, _23532_);
  or (_23536_, _23521_, _02549_);
  and (_23537_, _23536_, _02054_);
  and (_23538_, _23537_, _23535_);
  or (_23539_, _23538_, _23514_);
  and (_23541_, _23539_, _02047_);
  or (_23542_, _23511_, _11223_);
  and (_23543_, _23528_, _02046_);
  and (_23544_, _23543_, _23542_);
  or (_23545_, _23544_, _05474_);
  or (_23546_, _23545_, _23541_);
  or (_23547_, _12932_, _06184_);
  or (_23548_, _23547_, _13041_);
  or (_23549_, _23548_, _13155_);
  or (_23550_, _23549_, _13272_);
  or (_23552_, _23550_, _13389_);
  or (_23553_, _23552_, _13507_);
  or (_23554_, _23553_, _13624_);
  and (_23555_, _23554_, _06816_);
  and (_23556_, _23555_, _23546_);
  or (_23557_, _23556_, _06815_);
  or (_23558_, _23557_, _23510_);
  and (_23559_, _23558_, _02191_);
  and (_23560_, _23559_, _23502_);
  and (_23561_, _09066_, _07131_);
  nor (_23563_, _09066_, _07131_);
  or (_23564_, _23563_, _23561_);
  nand (_23565_, _23564_, _07203_);
  or (_23566_, _23564_, _07203_);
  and (_23567_, _23566_, _23565_);
  and (_23568_, _23567_, _02186_);
  or (_23569_, _23568_, _06740_);
  or (_23570_, _23569_, _23560_);
  not (_23571_, _06747_);
  and (_23572_, _06810_, _23571_);
  and (_23573_, _23572_, _09082_);
  nor (_23574_, _23572_, _09082_);
  or (_23575_, _23574_, _23573_);
  or (_23576_, _23575_, _06741_);
  and (_23577_, _23576_, _02043_);
  and (_23578_, _23577_, _23570_);
  nor (_23579_, _11241_, _23403_);
  or (_23580_, _23579_, _23511_);
  and (_23581_, _23580_, _02042_);
  or (_23582_, _23581_, _06188_);
  or (_23584_, _23582_, _23578_);
  and (_23585_, _23584_, _23492_);
  or (_23586_, _23585_, _02031_);
  and (_23587_, _05211_, _03838_);
  or (_23588_, _23485_, _02032_);
  or (_23589_, _23588_, _23587_);
  and (_23590_, _23589_, _02037_);
  and (_23591_, _23590_, _23586_);
  or (_23592_, _23591_, _23489_);
  and (_23593_, _23592_, _06560_);
  nor (_23595_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and (_23596_, _23595_, _06230_);
  nand (_23597_, _23596_, _06202_);
  nand (_23598_, _23597_, _02212_);
  or (_23599_, _23598_, _23593_);
  and (_23600_, _11189_, _03838_);
  or (_23601_, _23485_, _03059_);
  or (_23602_, _23601_, _23600_);
  and (_23603_, _03838_, _04866_);
  or (_23604_, _23603_, _23485_);
  or (_23606_, _23604_, _01995_);
  and (_23607_, _23606_, _03061_);
  and (_23608_, _23607_, _23602_);
  and (_23609_, _23608_, _23599_);
  and (_23610_, _11315_, _03838_);
  or (_23611_, _23610_, _23485_);
  and (_23612_, _23611_, _02331_);
  or (_23613_, _23612_, _23609_);
  and (_23614_, _23613_, _02208_);
  or (_23615_, _23485_, _04309_);
  and (_23617_, _23604_, _02206_);
  and (_23618_, _23617_, _23615_);
  or (_23619_, _23618_, _23614_);
  and (_23620_, _23619_, _03065_);
  and (_23621_, _23521_, _02342_);
  and (_23622_, _23621_, _23615_);
  or (_23623_, _23622_, _02202_);
  or (_23624_, _23623_, _23620_);
  nor (_23625_, _11187_, _08489_);
  or (_23626_, _23485_, _04953_);
  or (_23628_, _23626_, _23625_);
  and (_23629_, _23628_, _04958_);
  and (_23630_, _23629_, _23624_);
  nor (_23631_, _11314_, _08489_);
  or (_23632_, _23631_, _23485_);
  and (_23633_, _23632_, _02334_);
  or (_23634_, _23633_, _07348_);
  or (_23635_, _23634_, _23630_);
  and (_23636_, _23635_, _23483_);
  or (_23637_, _23636_, _06654_);
  and (_23639_, _23494_, _07377_);
  and (_23640_, _23495_, _08464_);
  nor (_23641_, _23640_, _23494_);
  and (_23642_, _23641_, _07380_);
  or (_23643_, _23642_, _23639_);
  or (_23644_, _23643_, _07356_);
  and (_23645_, _23644_, _02346_);
  and (_23646_, _23645_, _23637_);
  nor (_23647_, _07408_, \oc8051_golden_model_1.ACC [7]);
  or (_23648_, _23647_, _07130_);
  and (_23649_, _07408_, \oc8051_golden_model_1.ACC [7]);
  or (_23650_, _23649_, _07132_);
  and (_23651_, _23650_, _23648_);
  or (_23652_, _23561_, _07384_);
  or (_23653_, _23652_, _23651_);
  and (_23654_, _23653_, _07386_);
  or (_23655_, _23654_, _23646_);
  nor (_23656_, _06745_, _09176_);
  nor (_23657_, _06746_, \oc8051_golden_model_1.ACC [7]);
  nor (_23658_, _23657_, _23656_);
  and (_23660_, _23658_, _09149_);
  nor (_23661_, _23660_, _23656_);
  and (_23662_, _23661_, _07439_);
  nor (_23663_, _23661_, _07439_);
  or (_23664_, _23663_, _23662_);
  or (_23665_, _23664_, _07417_);
  and (_23666_, _23665_, _06614_);
  and (_23667_, _23666_, _23655_);
  or (_23668_, _23667_, _23473_);
  and (_23669_, _23668_, _07448_);
  nand (_23671_, _07480_, _09162_);
  and (_23672_, _23671_, _09164_);
  or (_23673_, _23672_, _23669_);
  and (_23674_, _23673_, _07488_);
  nor (_23675_, _09170_, _02087_);
  or (_23676_, _07526_, _07490_);
  and (_23677_, _23676_, _23675_);
  nor (_23678_, _07565_, _07278_);
  nor (_23679_, _23678_, _08458_);
  and (_23680_, _23679_, _09177_);
  or (_23682_, _23680_, _02366_);
  or (_23683_, _23682_, _23677_);
  or (_23684_, _23683_, _23674_);
  or (_23685_, _23516_, _02778_);
  and (_23686_, _23685_, _01698_);
  and (_23687_, _23686_, _23684_);
  and (_23688_, _23513_, _01697_);
  or (_23689_, _23688_, _02081_);
  or (_23690_, _23689_, _23687_);
  and (_23691_, _11367_, _03838_);
  or (_23693_, _23691_, _23485_);
  or (_23694_, _23693_, _02082_);
  and (_23695_, _23694_, _23690_);
  or (_23696_, _23695_, _39633_);
  or (_23697_, _39632_, \oc8051_golden_model_1.PSW [2]);
  and (_23698_, _23697_, _39026_);
  and (_41703_, _23698_, _23696_);
  not (_23699_, \oc8051_golden_model_1.PSW [3]);
  nor (_23700_, _03838_, _23699_);
  and (_23701_, _03838_, _04719_);
  nor (_23703_, _23701_, _23700_);
  and (_23704_, _23703_, _01994_);
  nor (_23705_, _08489_, _03434_);
  nor (_23706_, _23705_, _23700_);
  and (_23707_, _23706_, _06188_);
  and (_23708_, _03838_, \oc8051_golden_model_1.ACC [3]);
  nor (_23709_, _23708_, _23700_);
  nor (_23710_, _23709_, _02063_);
  nor (_23711_, _02062_, _23699_);
  or (_23712_, _23711_, _23710_);
  and (_23714_, _23712_, _03006_);
  nor (_23715_, _11394_, _08489_);
  nor (_23716_, _23715_, _23700_);
  nor (_23717_, _23716_, _03006_);
  or (_23718_, _23717_, _23714_);
  and (_23719_, _23718_, _02058_);
  nor (_23720_, _04476_, _23699_);
  and (_23721_, _11398_, _04476_);
  nor (_23722_, _23721_, _23720_);
  nor (_23723_, _23722_, _02058_);
  or (_23724_, _23723_, _23719_);
  and (_23725_, _23724_, _02519_);
  nor (_23726_, _23706_, _02519_);
  or (_23727_, _23726_, _23725_);
  and (_23728_, _23727_, _02549_);
  nor (_23729_, _23709_, _02549_);
  or (_23730_, _23729_, _23728_);
  and (_23731_, _23730_, _02054_);
  and (_23732_, _11408_, _04476_);
  nor (_23733_, _23732_, _23720_);
  nor (_23735_, _23733_, _02054_);
  or (_23736_, _23735_, _02046_);
  or (_23737_, _23736_, _23731_);
  nor (_23738_, _23720_, _11415_);
  nor (_23739_, _23738_, _23722_);
  or (_23740_, _23739_, _02047_);
  and (_23741_, _23740_, _02043_);
  and (_23742_, _23741_, _23737_);
  nor (_23743_, _11433_, _23403_);
  nor (_23744_, _23743_, _23720_);
  nor (_23746_, _23744_, _02043_);
  nor (_23747_, _23746_, _06188_);
  not (_23748_, _23747_);
  nor (_23749_, _23748_, _23742_);
  nor (_23750_, _23749_, _23707_);
  nor (_23751_, _23750_, _02031_);
  and (_23752_, _05166_, _03838_);
  nor (_23753_, _23700_, _02032_);
  not (_23754_, _23753_);
  nor (_23755_, _23754_, _23752_);
  or (_23757_, _23755_, _01765_);
  nor (_23758_, _23757_, _23751_);
  nor (_23759_, _11490_, _08489_);
  nor (_23760_, _23700_, _23759_);
  nor (_23761_, _23760_, _02037_);
  or (_23762_, _23761_, _01994_);
  nor (_23763_, _23762_, _23758_);
  nor (_23764_, _23763_, _23704_);
  or (_23765_, _23764_, _02210_);
  and (_23766_, _11505_, _03838_);
  or (_23768_, _23766_, _23700_);
  or (_23769_, _23768_, _03059_);
  and (_23770_, _23769_, _03061_);
  and (_23771_, _23770_, _23765_);
  and (_23772_, _11511_, _03838_);
  nor (_23773_, _23772_, _23700_);
  nor (_23774_, _23773_, _03061_);
  nor (_23775_, _23774_, _23771_);
  nor (_23776_, _23775_, _02206_);
  nor (_23777_, _23700_, _04153_);
  not (_23779_, _23777_);
  nor (_23780_, _23703_, _02208_);
  and (_23781_, _23780_, _23779_);
  nor (_23782_, _23781_, _23776_);
  nor (_23783_, _23782_, _02342_);
  or (_23784_, _23777_, _03065_);
  nor (_23785_, _23784_, _23709_);
  or (_23786_, _23785_, _02202_);
  nor (_23787_, _23786_, _23783_);
  nor (_23788_, _11503_, _08489_);
  or (_23790_, _23700_, _04953_);
  nor (_23791_, _23790_, _23788_);
  or (_23792_, _23791_, _02334_);
  nor (_23793_, _23792_, _23787_);
  nor (_23794_, _11510_, _08489_);
  nor (_23795_, _23794_, _23700_);
  nor (_23796_, _23795_, _04958_);
  or (_23797_, _23796_, _23793_);
  and (_23798_, _23797_, _02778_);
  nor (_23799_, _23716_, _02778_);
  or (_23800_, _23799_, _23798_);
  and (_23801_, _23800_, _01698_);
  nor (_23802_, _23733_, _01698_);
  or (_23803_, _23802_, _23801_);
  and (_23804_, _23803_, _02082_);
  and (_23805_, _11567_, _03838_);
  nor (_23806_, _23805_, _23700_);
  nor (_23807_, _23806_, _02082_);
  or (_23808_, _23807_, _23804_);
  or (_23809_, _23808_, _39633_);
  or (_23811_, _39632_, \oc8051_golden_model_1.PSW [3]);
  and (_23812_, _23811_, _39026_);
  and (_41704_, _23812_, _23809_);
  not (_23813_, \oc8051_golden_model_1.PSW [4]);
  nor (_23814_, _03838_, _23813_);
  and (_23815_, _04831_, _03838_);
  nor (_23816_, _23815_, _23814_);
  and (_23817_, _23816_, _01994_);
  nor (_23818_, _04372_, _08489_);
  nor (_23819_, _23818_, _23814_);
  and (_23821_, _23819_, _06188_);
  and (_23822_, _03838_, \oc8051_golden_model_1.ACC [4]);
  nor (_23823_, _23822_, _23814_);
  nor (_23824_, _23823_, _02063_);
  nor (_23825_, _02062_, _23813_);
  or (_23826_, _23825_, _23824_);
  and (_23827_, _23826_, _03006_);
  nor (_23828_, _11611_, _08489_);
  nor (_23829_, _23828_, _23814_);
  nor (_23830_, _23829_, _03006_);
  or (_23832_, _23830_, _23827_);
  and (_23833_, _23832_, _02058_);
  nor (_23834_, _04476_, _23813_);
  and (_23835_, _11597_, _04476_);
  nor (_23836_, _23835_, _23834_);
  nor (_23837_, _23836_, _02058_);
  or (_23838_, _23837_, _23833_);
  and (_23839_, _23838_, _02519_);
  nor (_23840_, _23819_, _02519_);
  or (_23841_, _23840_, _23839_);
  and (_23843_, _23841_, _02549_);
  nor (_23844_, _23823_, _02549_);
  or (_23845_, _23844_, _23843_);
  and (_23846_, _23845_, _02054_);
  and (_23847_, _11595_, _04476_);
  nor (_23848_, _23847_, _23834_);
  nor (_23849_, _23848_, _02054_);
  or (_23850_, _23849_, _23846_);
  and (_23851_, _23850_, _02047_);
  nor (_23852_, _23834_, _11628_);
  nor (_23854_, _23852_, _23836_);
  and (_23855_, _23854_, _02046_);
  or (_23856_, _23855_, _23851_);
  and (_23857_, _23856_, _02043_);
  nor (_23858_, _11646_, _23403_);
  nor (_23859_, _23858_, _23834_);
  nor (_23860_, _23859_, _02043_);
  nor (_23861_, _23860_, _06188_);
  not (_23862_, _23861_);
  nor (_23863_, _23862_, _23857_);
  nor (_23865_, _23863_, _23821_);
  nor (_23866_, _23865_, _02031_);
  and (_23867_, _05303_, _03838_);
  nor (_23868_, _23814_, _02032_);
  not (_23869_, _23868_);
  nor (_23870_, _23869_, _23867_);
  or (_23871_, _23870_, _01765_);
  nor (_23872_, _23871_, _23866_);
  nor (_23873_, _11704_, _08489_);
  nor (_23874_, _23814_, _23873_);
  nor (_23875_, _23874_, _02037_);
  or (_23876_, _23875_, _01994_);
  nor (_23877_, _23876_, _23872_);
  nor (_23878_, _23877_, _23817_);
  or (_23879_, _23878_, _02210_);
  and (_23880_, _11592_, _03838_);
  or (_23881_, _23880_, _23814_);
  or (_23882_, _23881_, _03059_);
  and (_23883_, _23882_, _03061_);
  and (_23884_, _23883_, _23879_);
  and (_23886_, _11588_, _03838_);
  nor (_23887_, _23886_, _23814_);
  nor (_23888_, _23887_, _03061_);
  nor (_23889_, _23888_, _23884_);
  nor (_23890_, _23889_, _02206_);
  nor (_23891_, _23814_, _04420_);
  not (_23892_, _23891_);
  nor (_23893_, _23816_, _02208_);
  and (_23894_, _23893_, _23892_);
  nor (_23895_, _23894_, _23890_);
  nor (_23897_, _23895_, _02342_);
  or (_23898_, _23891_, _03065_);
  nor (_23899_, _23898_, _23823_);
  or (_23900_, _23899_, _02202_);
  nor (_23901_, _23900_, _23897_);
  nor (_23902_, _11590_, _08489_);
  or (_23903_, _23814_, _04953_);
  nor (_23904_, _23903_, _23902_);
  or (_23905_, _23904_, _02334_);
  nor (_23906_, _23905_, _23901_);
  nor (_23908_, _11587_, _08489_);
  nor (_23909_, _23908_, _23814_);
  nor (_23910_, _23909_, _04958_);
  or (_23911_, _23910_, _23906_);
  and (_23912_, _23911_, _02778_);
  nor (_23913_, _23829_, _02778_);
  or (_23914_, _23913_, _23912_);
  and (_23915_, _23914_, _01698_);
  nor (_23916_, _23848_, _01698_);
  or (_23917_, _23916_, _23915_);
  and (_23919_, _23917_, _02082_);
  and (_23920_, _11771_, _03838_);
  nor (_23921_, _23920_, _23814_);
  nor (_23922_, _23921_, _02082_);
  or (_23923_, _23922_, _23919_);
  or (_23924_, _23923_, _39633_);
  or (_23925_, _39632_, \oc8051_golden_model_1.PSW [4]);
  and (_23926_, _23925_, _39026_);
  and (_41705_, _23926_, _23924_);
  not (_23927_, \oc8051_golden_model_1.PSW [5]);
  nor (_23929_, _03838_, _23927_);
  and (_23930_, _04827_, _03838_);
  nor (_23931_, _23930_, _23929_);
  and (_23932_, _23931_, _01994_);
  nor (_23933_, _04057_, _08489_);
  nor (_23934_, _23933_, _23929_);
  and (_23935_, _23934_, _06188_);
  and (_23936_, _03838_, \oc8051_golden_model_1.ACC [5]);
  nor (_23937_, _23936_, _23929_);
  nor (_23938_, _23937_, _02063_);
  nor (_23940_, _02062_, _23927_);
  or (_23941_, _23940_, _23938_);
  and (_23942_, _23941_, _03006_);
  nor (_23943_, _11804_, _08489_);
  nor (_23944_, _23943_, _23929_);
  nor (_23945_, _23944_, _03006_);
  or (_23946_, _23945_, _23942_);
  and (_23947_, _23946_, _02058_);
  nor (_23948_, _04476_, _23927_);
  and (_23949_, _11789_, _04476_);
  nor (_23950_, _23949_, _23948_);
  nor (_23951_, _23950_, _02058_);
  or (_23952_, _23951_, _23947_);
  and (_23953_, _23952_, _02519_);
  nor (_23954_, _23934_, _02519_);
  or (_23955_, _23954_, _23953_);
  and (_23956_, _23955_, _02549_);
  nor (_23957_, _23937_, _02549_);
  or (_23958_, _23957_, _23956_);
  and (_23959_, _23958_, _02054_);
  and (_23961_, _11816_, _04476_);
  nor (_23962_, _23961_, _23948_);
  nor (_23963_, _23962_, _02054_);
  or (_23964_, _23963_, _23959_);
  and (_23965_, _23964_, _02047_);
  nor (_23966_, _23948_, _11823_);
  nor (_23967_, _23966_, _23950_);
  and (_23968_, _23967_, _02046_);
  or (_23969_, _23968_, _23965_);
  and (_23970_, _23969_, _02043_);
  nor (_23972_, _11841_, _23403_);
  nor (_23973_, _23972_, _23948_);
  nor (_23974_, _23973_, _02043_);
  nor (_23975_, _23974_, _06188_);
  not (_23976_, _23975_);
  nor (_23977_, _23976_, _23970_);
  nor (_23978_, _23977_, _23935_);
  nor (_23979_, _23978_, _02031_);
  and (_23980_, _05258_, _03838_);
  nor (_23981_, _23929_, _02032_);
  not (_23983_, _23981_);
  nor (_23984_, _23983_, _23980_);
  or (_23985_, _23984_, _01765_);
  nor (_23986_, _23985_, _23979_);
  nor (_23987_, _11900_, _08489_);
  nor (_23988_, _23987_, _23929_);
  nor (_23989_, _23988_, _02037_);
  or (_23990_, _23989_, _01994_);
  nor (_23991_, _23990_, _23986_);
  nor (_23992_, _23991_, _23932_);
  or (_23994_, _23992_, _02210_);
  and (_23995_, _11915_, _03838_);
  or (_23996_, _23995_, _23929_);
  or (_23997_, _23996_, _03059_);
  and (_23998_, _23997_, _03061_);
  and (_23999_, _23998_, _23994_);
  and (_24000_, _11786_, _03838_);
  nor (_24001_, _24000_, _23929_);
  nor (_24002_, _24001_, _03061_);
  nor (_24003_, _24002_, _23999_);
  nor (_24005_, _24003_, _02206_);
  nor (_24006_, _23929_, _04104_);
  not (_24007_, _24006_);
  nor (_24008_, _23931_, _02208_);
  and (_24009_, _24008_, _24007_);
  nor (_24010_, _24009_, _24005_);
  nor (_24011_, _24010_, _02342_);
  or (_24012_, _24006_, _03065_);
  nor (_24013_, _24012_, _23937_);
  or (_24014_, _24013_, _02202_);
  nor (_24016_, _24014_, _24011_);
  nor (_24017_, _11913_, _08489_);
  or (_24018_, _23929_, _04953_);
  nor (_24019_, _24018_, _24017_);
  or (_24020_, _24019_, _02334_);
  nor (_24021_, _24020_, _24016_);
  nor (_24022_, _11785_, _08489_);
  nor (_24023_, _24022_, _23929_);
  nor (_24024_, _24023_, _04958_);
  or (_24025_, _24024_, _24021_);
  and (_24027_, _24025_, _02778_);
  nor (_24028_, _23944_, _02778_);
  or (_24029_, _24028_, _24027_);
  and (_24030_, _24029_, _01698_);
  nor (_24031_, _23962_, _01698_);
  or (_24032_, _24031_, _24030_);
  and (_24033_, _24032_, _02082_);
  and (_24034_, _11974_, _03838_);
  nor (_24035_, _24034_, _23929_);
  nor (_24036_, _24035_, _02082_);
  or (_24038_, _24036_, _24033_);
  or (_24039_, _24038_, _39633_);
  or (_24040_, _39632_, \oc8051_golden_model_1.PSW [5]);
  and (_24041_, _24040_, _39026_);
  and (_41706_, _24041_, _24039_);
  nor (_24042_, _07474_, _07448_);
  and (_24043_, _06643_, _09155_);
  not (_24044_, _07402_);
  nor (_24045_, _24044_, _07098_);
  nor (_24046_, _24045_, _02346_);
  nor (_24048_, _06730_, _06678_);
  and (_24049_, _24048_, _06717_);
  nor (_24050_, _03838_, _14600_);
  nor (_24051_, _03964_, _08489_);
  nor (_24052_, _24051_, _24050_);
  and (_24053_, _24052_, _06188_);
  or (_24054_, _07005_, _06961_);
  and (_24055_, _24054_, _06815_);
  and (_24056_, _03838_, \oc8051_golden_model_1.ACC [6]);
  nor (_24057_, _24056_, _24050_);
  nor (_24059_, _24057_, _02063_);
  nor (_24060_, _02062_, _14600_);
  or (_24061_, _24060_, _24059_);
  and (_24062_, _24061_, _03006_);
  nor (_24063_, _11993_, _08489_);
  nor (_24064_, _24063_, _24050_);
  nor (_24065_, _24064_, _03006_);
  or (_24066_, _24065_, _24062_);
  and (_24067_, _24066_, _02058_);
  nor (_24068_, _04476_, _14600_);
  and (_24070_, _11990_, _04476_);
  nor (_24071_, _24070_, _24068_);
  nor (_24072_, _24071_, _02058_);
  or (_24073_, _24072_, _24067_);
  and (_24074_, _24073_, _02519_);
  nor (_24075_, _24052_, _02519_);
  or (_24076_, _24075_, _24074_);
  and (_24077_, _24076_, _02549_);
  nor (_24078_, _24057_, _02549_);
  or (_24079_, _24078_, _24077_);
  and (_24081_, _24079_, _02054_);
  and (_24082_, _12017_, _04476_);
  nor (_24083_, _24082_, _24068_);
  nor (_24084_, _24083_, _02054_);
  nor (_24085_, _24084_, _24081_);
  nor (_24086_, _24085_, _02046_);
  nor (_24087_, _24068_, _12024_);
  or (_24088_, _24071_, _02047_);
  nor (_24089_, _24088_, _24087_);
  nor (_24090_, _24089_, _06817_);
  not (_24092_, _24090_);
  nor (_24093_, _24092_, _24086_);
  or (_24094_, _06816_, _06678_);
  nor (_24095_, _24094_, _06927_);
  or (_24096_, _24095_, _06815_);
  nor (_24097_, _24096_, _24093_);
  or (_24098_, _24097_, _24055_);
  and (_24099_, _24098_, _02191_);
  nor (_24100_, _07199_, _07098_);
  nor (_24101_, _24100_, _02191_);
  nor (_24102_, _24101_, _24099_);
  nor (_24103_, _24102_, _06740_);
  nor (_24104_, _06803_, _06743_);
  nor (_24105_, _24104_, _06741_);
  or (_24106_, _24105_, _24103_);
  and (_24107_, _24106_, _02043_);
  nor (_24108_, _12042_, _23403_);
  nor (_24109_, _24108_, _24068_);
  nor (_24110_, _24109_, _02043_);
  nor (_24111_, _24110_, _06188_);
  not (_24113_, _24111_);
  nor (_24114_, _24113_, _24107_);
  nor (_24115_, _24114_, _24053_);
  nor (_24116_, _24115_, _02031_);
  and (_24117_, _05029_, _03838_);
  nor (_24118_, _24050_, _02032_);
  not (_24119_, _24118_);
  nor (_24120_, _24119_, _24117_);
  nor (_24121_, _24120_, _01765_);
  not (_24122_, _24121_);
  nor (_24124_, _24122_, _24116_);
  nor (_24125_, _12096_, _08489_);
  nor (_24126_, _24125_, _24050_);
  nor (_24127_, _24126_, _02037_);
  or (_24128_, _24127_, _07629_);
  or (_24129_, _24128_, _24124_);
  and (_24130_, _12112_, _03838_);
  or (_24131_, _24050_, _03059_);
  or (_24132_, _24131_, _24130_);
  and (_24133_, _12103_, _03838_);
  nor (_24135_, _24133_, _24050_);
  and (_24136_, _24135_, _01994_);
  nor (_24137_, _24136_, _02331_);
  and (_24138_, _24137_, _24132_);
  and (_24139_, _24138_, _24129_);
  and (_24140_, _12118_, _03838_);
  nor (_24141_, _24140_, _24050_);
  nor (_24142_, _24141_, _03061_);
  nor (_24143_, _24142_, _24139_);
  nor (_24144_, _24143_, _02206_);
  nor (_24146_, _24050_, _04011_);
  not (_24147_, _24146_);
  nor (_24148_, _24135_, _02208_);
  and (_24149_, _24148_, _24147_);
  nor (_24150_, _24149_, _24144_);
  nor (_24151_, _24150_, _02342_);
  or (_24152_, _24146_, _03065_);
  nor (_24153_, _24152_, _24057_);
  or (_24154_, _24153_, _02202_);
  nor (_24155_, _24154_, _24151_);
  nor (_24157_, _12110_, _08489_);
  or (_24158_, _24050_, _04953_);
  or (_24159_, _24158_, _24157_);
  and (_24160_, _24159_, _04958_);
  not (_24161_, _24160_);
  nor (_24162_, _24161_, _24155_);
  nor (_24163_, _12117_, _08489_);
  nor (_24164_, _24163_, _24050_);
  nor (_24165_, _24164_, _04958_);
  nor (_24166_, _24165_, _07348_);
  not (_24168_, _24166_);
  nor (_24169_, _24168_, _24162_);
  nor (_24170_, _24169_, _24049_);
  nor (_24171_, _24170_, _06654_);
  nor (_24172_, _06961_, _07356_);
  nand (_24173_, _24172_, _07371_);
  and (_24174_, _24173_, _02346_);
  not (_24175_, _24174_);
  nor (_24176_, _24175_, _24171_);
  nor (_24177_, _24176_, _24046_);
  nor (_24178_, _24177_, _07384_);
  not (_24179_, _06743_);
  and (_24180_, _07430_, _24179_);
  nor (_24181_, _24180_, _07417_);
  nor (_24182_, _24181_, _09155_);
  not (_24183_, _24182_);
  nor (_24184_, _24183_, _24178_);
  nor (_24185_, _24184_, _24043_);
  nor (_24186_, _24185_, _06609_);
  or (_24187_, _24186_, _02085_);
  nor (_24189_, _24187_, _24042_);
  and (_24190_, _07520_, _02085_);
  or (_24191_, _24190_, _07487_);
  nor (_24192_, _24191_, _24189_);
  nor (_24193_, _07559_, _08458_);
  nor (_24194_, _24193_, _24192_);
  and (_24195_, _24194_, _02778_);
  nor (_24196_, _24064_, _02778_);
  or (_24197_, _24196_, _24195_);
  and (_24198_, _24197_, _01698_);
  nor (_24200_, _24083_, _01698_);
  or (_24201_, _24200_, _24198_);
  and (_24202_, _24201_, _02082_);
  and (_24203_, _12178_, _03838_);
  nor (_24204_, _24203_, _24050_);
  nor (_24205_, _24204_, _02082_);
  or (_24206_, _24205_, _24202_);
  or (_24207_, _24206_, _39633_);
  or (_24208_, _39632_, \oc8051_golden_model_1.PSW [6]);
  and (_24209_, _24208_, _39026_);
  and (_41707_, _24209_, _24207_);
  not (_24211_, \oc8051_golden_model_1.PCON [0]);
  nor (_24212_, _03828_, _24211_);
  nor (_24213_, _04257_, _09201_);
  nor (_24214_, _24213_, _24212_);
  and (_24215_, _24214_, _15890_);
  and (_24216_, _03828_, _04837_);
  nor (_24217_, _24216_, _24212_);
  nor (_24218_, _24217_, _02208_);
  not (_24219_, _24218_);
  nor (_24221_, _24219_, _24213_);
  and (_24222_, _03828_, \oc8051_golden_model_1.ACC [0]);
  nor (_24223_, _24222_, _24212_);
  nor (_24224_, _24223_, _02549_);
  nor (_24225_, _24224_, _06188_);
  nor (_24226_, _24214_, _03006_);
  nor (_24227_, _02062_, _24211_);
  nor (_24228_, _24223_, _02063_);
  nor (_24229_, _24228_, _24227_);
  nor (_24230_, _24229_, _02158_);
  or (_24232_, _24230_, _02155_);
  nor (_24233_, _24232_, _24226_);
  or (_24234_, _24233_, _02153_);
  and (_24235_, _24234_, _24225_);
  and (_24236_, _03828_, _03002_);
  and (_24237_, _05444_, _02519_);
  or (_24238_, _24237_, _24212_);
  nor (_24239_, _24238_, _24236_);
  nor (_24240_, _24239_, _24235_);
  nor (_24241_, _24240_, _02031_);
  and (_24243_, _05120_, _03828_);
  nor (_24244_, _24212_, _02032_);
  not (_24245_, _24244_);
  nor (_24246_, _24245_, _24243_);
  nor (_24247_, _24246_, _24241_);
  nor (_24248_, _24247_, _01765_);
  nor (_24249_, _10898_, _09201_);
  or (_24250_, _24212_, _02037_);
  nor (_24251_, _24250_, _24249_);
  or (_24252_, _24251_, _01994_);
  nor (_24254_, _24252_, _24248_);
  nand (_24255_, _24217_, _03059_);
  and (_24256_, _24255_, _07629_);
  nor (_24257_, _24256_, _24254_);
  and (_24258_, _10914_, _03828_);
  nor (_24259_, _24258_, _24212_);
  and (_24260_, _24259_, _02210_);
  nor (_24261_, _24260_, _24257_);
  and (_24262_, _24261_, _03061_);
  and (_24263_, _10792_, _03828_);
  nor (_24265_, _24263_, _24212_);
  nor (_24266_, _24265_, _03061_);
  or (_24267_, _24266_, _24262_);
  and (_24268_, _24267_, _02208_);
  nor (_24269_, _24268_, _24221_);
  nor (_24270_, _24269_, _02342_);
  and (_24271_, _10791_, _03828_);
  or (_24272_, _24271_, _24212_);
  and (_24273_, _24272_, _02342_);
  or (_24274_, _24273_, _24270_);
  and (_24275_, _24274_, _04953_);
  nor (_24276_, _10913_, _09201_);
  nor (_24277_, _24276_, _24212_);
  nor (_24278_, _24277_, _04953_);
  or (_24279_, _24278_, _24275_);
  and (_24280_, _24279_, _04958_);
  nor (_24281_, _10789_, _09201_);
  nor (_24282_, _24281_, _24212_);
  nor (_24283_, _24282_, _04958_);
  nor (_24284_, _24283_, _15890_);
  not (_24286_, _24284_);
  nor (_24287_, _24286_, _24280_);
  nor (_24288_, _24287_, _24215_);
  or (_24289_, _24288_, _39633_);
  or (_24290_, _39632_, \oc8051_golden_model_1.PCON [0]);
  and (_24291_, _24290_, _39026_);
  and (_41709_, _24291_, _24289_);
  nor (_24292_, _03828_, \oc8051_golden_model_1.PCON [1]);
  not (_24293_, _24292_);
  nor (_24294_, _10988_, _09201_);
  nor (_24296_, _24294_, _02208_);
  and (_24297_, _24296_, _24293_);
  nor (_24298_, _11113_, _09201_);
  nor (_24299_, _24298_, _03061_);
  and (_24300_, _24299_, _24293_);
  and (_24301_, _05075_, _03828_);
  not (_24302_, \oc8051_golden_model_1.PCON [1]);
  nor (_24303_, _03828_, _24302_);
  nor (_24304_, _24303_, _02032_);
  not (_24305_, _24304_);
  nor (_24307_, _24305_, _24301_);
  not (_24308_, _24307_);
  and (_24309_, _03828_, _01804_);
  nor (_24310_, _24309_, _24292_);
  and (_24311_, _24310_, _02153_);
  and (_24312_, _24310_, _02062_);
  nor (_24313_, _02062_, _24302_);
  or (_24314_, _24313_, _24312_);
  and (_24315_, _24314_, _03006_);
  and (_24316_, _11001_, _03828_);
  nor (_24318_, _24316_, _24292_);
  and (_24319_, _24318_, _02158_);
  or (_24320_, _24319_, _24315_);
  and (_24321_, _24320_, _02519_);
  nor (_24322_, _09201_, _03161_);
  nor (_24323_, _24322_, _24303_);
  nor (_24324_, _24323_, _02519_);
  nor (_24325_, _24324_, _24321_);
  nor (_24326_, _24325_, _02153_);
  or (_24327_, _24326_, _06188_);
  nor (_24329_, _24327_, _24311_);
  and (_24330_, _24323_, _06188_);
  nor (_24331_, _24330_, _24329_);
  nor (_24332_, _24331_, _02031_);
  nor (_24333_, _24332_, _01765_);
  and (_24334_, _24333_, _24308_);
  and (_24335_, _11096_, _03828_);
  nor (_24336_, _24335_, _02037_);
  and (_24337_, _24336_, _24293_);
  nor (_24338_, _24337_, _24334_);
  nor (_24340_, _24338_, _07629_);
  nor (_24341_, _10989_, _09201_);
  nor (_24342_, _24341_, _03059_);
  and (_24343_, _03828_, _02893_);
  nor (_24344_, _24343_, _01995_);
  nor (_24345_, _24344_, _24342_);
  nor (_24346_, _24345_, _24292_);
  nor (_24347_, _24346_, _24340_);
  nor (_24348_, _24347_, _02331_);
  nor (_24349_, _24348_, _24300_);
  nor (_24351_, _24349_, _02206_);
  nor (_24352_, _24351_, _24297_);
  nor (_24353_, _24352_, _02342_);
  nor (_24354_, _24303_, _04209_);
  nor (_24355_, _24354_, _03065_);
  and (_24356_, _24355_, _24310_);
  nor (_24357_, _24356_, _24353_);
  or (_24358_, _24357_, _17216_);
  and (_24359_, _24309_, _04208_);
  nor (_24360_, _24359_, _04958_);
  and (_24362_, _24360_, _24293_);
  nor (_24363_, _24362_, _02366_);
  and (_24364_, _24343_, _04208_);
  or (_24365_, _24292_, _04953_);
  or (_24366_, _24365_, _24364_);
  and (_24367_, _24366_, _24363_);
  and (_24368_, _24367_, _24358_);
  nor (_24369_, _24318_, _02778_);
  nor (_24370_, _24369_, _24368_);
  nor (_24371_, _24370_, _02081_);
  nor (_24372_, _24316_, _24303_);
  and (_24373_, _24372_, _02081_);
  nor (_24374_, _24373_, _24371_);
  or (_24375_, _24374_, _39633_);
  or (_24376_, _39632_, \oc8051_golden_model_1.PCON [1]);
  and (_24377_, _24376_, _39026_);
  and (_41710_, _24377_, _24375_);
  not (_24378_, \oc8051_golden_model_1.PCON [2]);
  nor (_24379_, _03828_, _24378_);
  nor (_24380_, _11314_, _09201_);
  nor (_24382_, _24380_, _24379_);
  nor (_24383_, _24382_, _04958_);
  and (_24384_, _11315_, _03828_);
  nor (_24385_, _24384_, _24379_);
  nor (_24386_, _24385_, _03061_);
  and (_24387_, _03828_, _04866_);
  nor (_24388_, _24387_, _24379_);
  and (_24389_, _24388_, _01994_);
  and (_24390_, _03828_, \oc8051_golden_model_1.ACC [2]);
  nor (_24391_, _24390_, _24379_);
  nor (_24393_, _24391_, _02549_);
  nor (_24394_, _24391_, _02063_);
  nor (_24395_, _02062_, _24378_);
  or (_24396_, _24395_, _24394_);
  and (_24397_, _24396_, _03006_);
  nor (_24398_, _11199_, _09201_);
  nor (_24399_, _24398_, _24379_);
  nor (_24400_, _24399_, _03006_);
  or (_24401_, _24400_, _24397_);
  and (_24402_, _24401_, _02519_);
  nor (_24404_, _09201_, _03624_);
  nor (_24405_, _24404_, _24379_);
  nor (_24406_, _24405_, _02519_);
  nor (_24407_, _24406_, _24402_);
  nor (_24408_, _24407_, _02153_);
  or (_24409_, _24408_, _06188_);
  nor (_24410_, _24409_, _24393_);
  and (_24411_, _24405_, _06188_);
  nor (_24412_, _24411_, _24410_);
  nor (_24413_, _24412_, _02031_);
  and (_24415_, _05211_, _03828_);
  nor (_24416_, _24379_, _02032_);
  not (_24417_, _24416_);
  nor (_24418_, _24417_, _24415_);
  or (_24419_, _24418_, _01765_);
  nor (_24420_, _24419_, _24413_);
  nor (_24421_, _11298_, _09201_);
  nor (_24422_, _24421_, _24379_);
  nor (_24423_, _24422_, _02037_);
  or (_24424_, _24423_, _01994_);
  nor (_24426_, _24424_, _24420_);
  nor (_24427_, _24426_, _24389_);
  or (_24428_, _24427_, _02210_);
  and (_24429_, _11189_, _03828_);
  or (_24430_, _24429_, _24379_);
  or (_24431_, _24430_, _03059_);
  and (_24432_, _24431_, _03061_);
  and (_24433_, _24432_, _24428_);
  nor (_24434_, _24433_, _24386_);
  nor (_24435_, _24434_, _02206_);
  nor (_24437_, _24379_, _04309_);
  not (_24438_, _24437_);
  nor (_24439_, _24388_, _02208_);
  and (_24440_, _24439_, _24438_);
  nor (_24441_, _24440_, _24435_);
  nor (_24442_, _24441_, _02342_);
  or (_24443_, _24437_, _03065_);
  nor (_24444_, _24443_, _24391_);
  or (_24445_, _24444_, _02202_);
  nor (_24446_, _24445_, _24442_);
  nor (_24448_, _11187_, _09201_);
  or (_24449_, _24379_, _04953_);
  nor (_24450_, _24449_, _24448_);
  or (_24451_, _24450_, _02334_);
  nor (_24452_, _24451_, _24446_);
  nor (_24453_, _24452_, _24383_);
  nor (_24454_, _24453_, _02366_);
  nor (_24455_, _24399_, _02778_);
  or (_24456_, _24455_, _02081_);
  nor (_24457_, _24456_, _24454_);
  and (_24459_, _11367_, _03828_);
  nor (_24460_, _24459_, _24379_);
  and (_24461_, _24460_, _02081_);
  nor (_24462_, _24461_, _24457_);
  or (_24463_, _24462_, _39633_);
  or (_24464_, _39632_, \oc8051_golden_model_1.PCON [2]);
  and (_24465_, _24464_, _39026_);
  and (_41711_, _24465_, _24463_);
  not (_24466_, \oc8051_golden_model_1.PCON [3]);
  nor (_24467_, _03828_, _24466_);
  nor (_24468_, _11510_, _09201_);
  nor (_24469_, _24468_, _24467_);
  nor (_24470_, _24469_, _04958_);
  nor (_24471_, _24467_, _04153_);
  not (_24472_, _24471_);
  and (_24473_, _03828_, _04719_);
  nor (_24474_, _24473_, _24467_);
  nor (_24475_, _24474_, _02208_);
  and (_24476_, _24475_, _24472_);
  and (_24477_, _11511_, _03828_);
  nor (_24479_, _24477_, _24467_);
  nor (_24480_, _24479_, _03061_);
  nor (_24481_, _09201_, _03434_);
  nor (_24482_, _24481_, _24467_);
  and (_24483_, _24482_, _06188_);
  and (_24484_, _03828_, \oc8051_golden_model_1.ACC [3]);
  nor (_24485_, _24484_, _24467_);
  nor (_24486_, _24485_, _02549_);
  nor (_24487_, _24485_, _02063_);
  nor (_24488_, _02062_, _24466_);
  or (_24490_, _24488_, _24487_);
  and (_24491_, _24490_, _03006_);
  nor (_24492_, _11394_, _09201_);
  nor (_24493_, _24492_, _24467_);
  nor (_24494_, _24493_, _03006_);
  or (_24495_, _24494_, _24491_);
  and (_24496_, _24495_, _02519_);
  nor (_24497_, _24482_, _02519_);
  nor (_24498_, _24497_, _24496_);
  nor (_24499_, _24498_, _02153_);
  or (_24501_, _24499_, _06188_);
  nor (_24502_, _24501_, _24486_);
  nor (_24503_, _24502_, _24483_);
  nor (_24504_, _24503_, _02031_);
  and (_24505_, _05166_, _03828_);
  nor (_24506_, _24467_, _02032_);
  not (_24507_, _24506_);
  nor (_24508_, _24507_, _24505_);
  nor (_24509_, _24508_, _01765_);
  not (_24510_, _24509_);
  nor (_24512_, _24510_, _24504_);
  nor (_24513_, _11490_, _09201_);
  nor (_24514_, _24513_, _24467_);
  nor (_24515_, _24514_, _02037_);
  or (_24516_, _24515_, _07629_);
  or (_24517_, _24516_, _24512_);
  and (_24518_, _11505_, _03828_);
  or (_24519_, _24467_, _03059_);
  or (_24520_, _24519_, _24518_);
  and (_24521_, _24474_, _01994_);
  nor (_24523_, _24521_, _02331_);
  and (_24524_, _24523_, _24520_);
  and (_24525_, _24524_, _24517_);
  nor (_24526_, _24525_, _24480_);
  nor (_24527_, _24526_, _02206_);
  nor (_24528_, _24527_, _24476_);
  nor (_24529_, _24528_, _02342_);
  or (_24530_, _24471_, _03065_);
  nor (_24531_, _24530_, _24485_);
  or (_24532_, _24531_, _02202_);
  nor (_24534_, _24532_, _24529_);
  nor (_24535_, _11503_, _09201_);
  or (_24536_, _24467_, _04953_);
  nor (_24537_, _24536_, _24535_);
  or (_24538_, _24537_, _02334_);
  nor (_24539_, _24538_, _24534_);
  nor (_24540_, _24539_, _24470_);
  nor (_24541_, _24540_, _02366_);
  nor (_24542_, _24493_, _02778_);
  or (_24543_, _24542_, _02081_);
  nor (_24545_, _24543_, _24541_);
  and (_24546_, _11567_, _03828_);
  nor (_24547_, _24546_, _24467_);
  and (_24548_, _24547_, _02081_);
  nor (_24549_, _24548_, _24545_);
  or (_24550_, _24549_, _39633_);
  or (_24551_, _39632_, \oc8051_golden_model_1.PCON [3]);
  and (_24552_, _24551_, _39026_);
  and (_41712_, _24552_, _24550_);
  not (_24553_, \oc8051_golden_model_1.PCON [4]);
  nor (_24555_, _03828_, _24553_);
  nor (_24556_, _11587_, _09201_);
  nor (_24557_, _24556_, _24555_);
  nor (_24558_, _24557_, _04958_);
  and (_24559_, _11588_, _03828_);
  nor (_24560_, _24559_, _24555_);
  nor (_24561_, _24560_, _03061_);
  and (_24562_, _05303_, _03828_);
  or (_24563_, _24562_, _24555_);
  and (_24564_, _24563_, _02031_);
  and (_24565_, _03828_, \oc8051_golden_model_1.ACC [4]);
  nor (_24566_, _24565_, _24555_);
  nor (_24567_, _24566_, _02549_);
  nor (_24568_, _24566_, _02063_);
  nor (_24569_, _02062_, _24553_);
  or (_24570_, _24569_, _24568_);
  and (_24571_, _24570_, _03006_);
  nor (_24572_, _11611_, _09201_);
  nor (_24573_, _24572_, _24555_);
  nor (_24574_, _24573_, _03006_);
  or (_24576_, _24574_, _24571_);
  and (_24577_, _24576_, _02519_);
  nor (_24578_, _04372_, _09201_);
  nor (_24579_, _24578_, _24555_);
  nor (_24580_, _24579_, _02519_);
  nor (_24581_, _24580_, _24577_);
  nor (_24582_, _24581_, _02153_);
  or (_24583_, _24582_, _06188_);
  nor (_24584_, _24583_, _24567_);
  and (_24585_, _24579_, _06188_);
  or (_24587_, _24585_, _02031_);
  nor (_24588_, _24587_, _24584_);
  or (_24589_, _24588_, _24564_);
  and (_24590_, _24589_, _02037_);
  nor (_24591_, _11704_, _09201_);
  nor (_24592_, _24591_, _24555_);
  nor (_24593_, _24592_, _02037_);
  or (_24594_, _24593_, _07629_);
  or (_24595_, _24594_, _24590_);
  and (_24596_, _11592_, _03828_);
  or (_24598_, _24555_, _03059_);
  or (_24599_, _24598_, _24596_);
  and (_24600_, _04831_, _03828_);
  nor (_24601_, _24600_, _24555_);
  and (_24602_, _24601_, _01994_);
  nor (_24603_, _24602_, _02331_);
  and (_24604_, _24603_, _24599_);
  and (_24605_, _24604_, _24595_);
  nor (_24606_, _24605_, _24561_);
  nor (_24607_, _24606_, _02206_);
  nor (_24609_, _24555_, _04420_);
  not (_24610_, _24609_);
  nor (_24611_, _24601_, _02208_);
  and (_24612_, _24611_, _24610_);
  nor (_24613_, _24612_, _24607_);
  nor (_24614_, _24613_, _02342_);
  or (_24615_, _24609_, _03065_);
  nor (_24616_, _24615_, _24566_);
  or (_24617_, _24616_, _02202_);
  nor (_24618_, _24617_, _24614_);
  nor (_24620_, _11590_, _09201_);
  or (_24621_, _24555_, _04953_);
  nor (_24622_, _24621_, _24620_);
  or (_24623_, _24622_, _02334_);
  nor (_24624_, _24623_, _24618_);
  nor (_24625_, _24624_, _24558_);
  nor (_24626_, _24625_, _02366_);
  nor (_24627_, _24573_, _02778_);
  or (_24628_, _24627_, _02081_);
  nor (_24629_, _24628_, _24626_);
  and (_24631_, _11771_, _03828_);
  nor (_24632_, _24631_, _24555_);
  and (_24633_, _24632_, _02081_);
  nor (_24634_, _24633_, _24629_);
  or (_24635_, _24634_, _39633_);
  or (_24636_, _39632_, \oc8051_golden_model_1.PCON [4]);
  and (_24637_, _24636_, _39026_);
  and (_41713_, _24637_, _24635_);
  not (_24638_, \oc8051_golden_model_1.PCON [5]);
  nor (_24639_, _03828_, _24638_);
  nor (_24641_, _11785_, _09201_);
  nor (_24642_, _24641_, _24639_);
  nor (_24643_, _24642_, _04958_);
  and (_24644_, _11786_, _03828_);
  nor (_24645_, _24644_, _24639_);
  nor (_24646_, _24645_, _03061_);
  and (_24647_, _04827_, _03828_);
  nor (_24648_, _24647_, _24639_);
  and (_24649_, _24648_, _01994_);
  and (_24650_, _03828_, \oc8051_golden_model_1.ACC [5]);
  nor (_24652_, _24650_, _24639_);
  nor (_24653_, _24652_, _02549_);
  nor (_24654_, _24652_, _02063_);
  nor (_24655_, _02062_, _24638_);
  or (_24656_, _24655_, _24654_);
  and (_24657_, _24656_, _03006_);
  nor (_24658_, _11804_, _09201_);
  nor (_24659_, _24658_, _24639_);
  nor (_24660_, _24659_, _03006_);
  or (_24661_, _24660_, _24657_);
  and (_24662_, _24661_, _02519_);
  nor (_24663_, _04057_, _09201_);
  nor (_24664_, _24663_, _24639_);
  nor (_24665_, _24664_, _02519_);
  nor (_24666_, _24665_, _24662_);
  nor (_24667_, _24666_, _02153_);
  or (_24668_, _24667_, _06188_);
  nor (_24669_, _24668_, _24653_);
  and (_24670_, _24664_, _06188_);
  nor (_24671_, _24670_, _24669_);
  nor (_24673_, _24671_, _02031_);
  and (_24674_, _05258_, _03828_);
  nor (_24675_, _24639_, _02032_);
  not (_24676_, _24675_);
  nor (_24677_, _24676_, _24674_);
  or (_24678_, _24677_, _01765_);
  nor (_24679_, _24678_, _24673_);
  nor (_24680_, _11900_, _09201_);
  nor (_24681_, _24680_, _24639_);
  nor (_24682_, _24681_, _02037_);
  or (_24684_, _24682_, _01994_);
  nor (_24685_, _24684_, _24679_);
  nor (_24686_, _24685_, _24649_);
  or (_24687_, _24686_, _02210_);
  and (_24688_, _11915_, _03828_);
  or (_24689_, _24688_, _24639_);
  or (_24690_, _24689_, _03059_);
  and (_24691_, _24690_, _03061_);
  and (_24692_, _24691_, _24687_);
  nor (_24693_, _24692_, _24646_);
  nor (_24695_, _24693_, _02206_);
  nor (_24696_, _24639_, _04104_);
  not (_24697_, _24696_);
  nor (_24698_, _24648_, _02208_);
  and (_24699_, _24698_, _24697_);
  nor (_24700_, _24699_, _24695_);
  nor (_24701_, _24700_, _02342_);
  or (_24702_, _24696_, _03065_);
  nor (_24703_, _24702_, _24652_);
  or (_24704_, _24703_, _02202_);
  nor (_24706_, _24704_, _24701_);
  nor (_24707_, _11913_, _09201_);
  or (_24708_, _24639_, _04953_);
  nor (_24709_, _24708_, _24707_);
  or (_24710_, _24709_, _02334_);
  nor (_24711_, _24710_, _24706_);
  nor (_24712_, _24711_, _24643_);
  nor (_24713_, _24712_, _02366_);
  nor (_24714_, _24659_, _02778_);
  or (_24715_, _24714_, _02081_);
  nor (_24717_, _24715_, _24713_);
  and (_24718_, _11974_, _03828_);
  nor (_24719_, _24718_, _24639_);
  and (_24720_, _24719_, _02081_);
  nor (_24721_, _24720_, _24717_);
  or (_24722_, _24721_, _39633_);
  or (_24723_, _39632_, \oc8051_golden_model_1.PCON [5]);
  and (_24724_, _24723_, _39026_);
  and (_41714_, _24724_, _24722_);
  not (_24725_, \oc8051_golden_model_1.PCON [6]);
  nor (_24727_, _03828_, _24725_);
  nor (_24728_, _12117_, _09201_);
  nor (_24729_, _24728_, _24727_);
  nor (_24730_, _24729_, _04958_);
  and (_24731_, _12118_, _03828_);
  nor (_24732_, _24731_, _24727_);
  nor (_24733_, _24732_, _03061_);
  and (_24734_, _12103_, _03828_);
  nor (_24735_, _24734_, _24727_);
  and (_24736_, _24735_, _01994_);
  nor (_24738_, _03964_, _09201_);
  nor (_24739_, _24738_, _24727_);
  and (_24740_, _24739_, _06188_);
  and (_24741_, _03828_, \oc8051_golden_model_1.ACC [6]);
  nor (_24742_, _24741_, _24727_);
  nor (_24743_, _24742_, _02549_);
  nor (_24744_, _24742_, _02063_);
  nor (_24745_, _02062_, _24725_);
  or (_24746_, _24745_, _24744_);
  and (_24747_, _24746_, _03006_);
  nor (_24749_, _11993_, _09201_);
  nor (_24750_, _24749_, _24727_);
  nor (_24751_, _24750_, _03006_);
  or (_24752_, _24751_, _24747_);
  and (_24753_, _24752_, _02519_);
  nor (_24754_, _24739_, _02519_);
  nor (_24755_, _24754_, _24753_);
  nor (_24756_, _24755_, _02153_);
  or (_24757_, _24756_, _06188_);
  nor (_24758_, _24757_, _24743_);
  nor (_24759_, _24758_, _24740_);
  nor (_24760_, _24759_, _02031_);
  and (_24761_, _05029_, _03828_);
  nor (_24762_, _24727_, _02032_);
  not (_24763_, _24762_);
  nor (_24764_, _24763_, _24761_);
  or (_24765_, _24764_, _01765_);
  nor (_24766_, _24765_, _24760_);
  nor (_24767_, _12096_, _09201_);
  nor (_24768_, _24767_, _24727_);
  nor (_24770_, _24768_, _02037_);
  or (_24771_, _24770_, _01994_);
  nor (_24772_, _24771_, _24766_);
  nor (_24773_, _24772_, _24736_);
  or (_24774_, _24773_, _02210_);
  and (_24775_, _12112_, _03828_);
  or (_24776_, _24775_, _24727_);
  or (_24777_, _24776_, _03059_);
  and (_24778_, _24777_, _03061_);
  and (_24779_, _24778_, _24774_);
  nor (_24781_, _24779_, _24733_);
  nor (_24782_, _24781_, _02206_);
  nor (_24783_, _24727_, _04011_);
  not (_24784_, _24783_);
  nor (_24785_, _24735_, _02208_);
  and (_24786_, _24785_, _24784_);
  nor (_24787_, _24786_, _24782_);
  nor (_24788_, _24787_, _02342_);
  or (_24789_, _24783_, _03065_);
  nor (_24790_, _24789_, _24742_);
  or (_24792_, _24790_, _02202_);
  nor (_24793_, _24792_, _24788_);
  nor (_24794_, _12110_, _09201_);
  or (_24795_, _24727_, _04953_);
  nor (_24796_, _24795_, _24794_);
  or (_24797_, _24796_, _02334_);
  nor (_24798_, _24797_, _24793_);
  nor (_24799_, _24798_, _24730_);
  nor (_24800_, _24799_, _02366_);
  nor (_24801_, _24750_, _02778_);
  or (_24803_, _24801_, _02081_);
  nor (_24804_, _24803_, _24800_);
  and (_24805_, _12178_, _03828_);
  nor (_24806_, _24805_, _24727_);
  and (_24807_, _24806_, _02081_);
  nor (_24808_, _24807_, _24804_);
  or (_24809_, _24808_, _39633_);
  or (_24810_, _39632_, \oc8051_golden_model_1.PCON [6]);
  and (_24811_, _24810_, _39026_);
  and (_41715_, _24811_, _24809_);
  not (_24813_, \oc8051_golden_model_1.SBUF [0]);
  nor (_24814_, _03805_, _24813_);
  nor (_24815_, _04257_, _09281_);
  nor (_24816_, _24815_, _24814_);
  and (_24817_, _24816_, _15890_);
  and (_24818_, _03805_, \oc8051_golden_model_1.ACC [0]);
  nor (_24819_, _24818_, _24814_);
  nor (_24820_, _24819_, _02549_);
  nor (_24821_, _24819_, _02063_);
  nor (_24822_, _02062_, _24813_);
  or (_24824_, _24822_, _24821_);
  and (_24825_, _24824_, _03006_);
  nor (_24826_, _24816_, _03006_);
  or (_24827_, _24826_, _24825_);
  and (_24828_, _24827_, _02519_);
  and (_24829_, _03805_, _03002_);
  nor (_24830_, _24829_, _24814_);
  nor (_24831_, _24830_, _02519_);
  nor (_24832_, _24831_, _24828_);
  nor (_24833_, _24832_, _02153_);
  or (_24835_, _24833_, _06188_);
  nor (_24836_, _24835_, _24820_);
  and (_24837_, _24830_, _06188_);
  nor (_24838_, _24837_, _24836_);
  nor (_24839_, _24838_, _02031_);
  and (_24840_, _05120_, _03805_);
  nor (_24841_, _24814_, _02032_);
  not (_24842_, _24841_);
  nor (_24843_, _24842_, _24840_);
  nor (_24844_, _24843_, _24839_);
  nor (_24846_, _24844_, _01765_);
  nor (_24847_, _10898_, _09281_);
  or (_24848_, _24814_, _02037_);
  nor (_24849_, _24848_, _24847_);
  or (_24850_, _24849_, _01994_);
  nor (_24851_, _24850_, _24846_);
  and (_24852_, _03805_, _04837_);
  nor (_24853_, _24852_, _24814_);
  nand (_24854_, _24853_, _03059_);
  and (_24855_, _24854_, _07629_);
  nor (_24856_, _24855_, _24851_);
  and (_24857_, _10914_, _03805_);
  nor (_24858_, _24857_, _24814_);
  and (_24859_, _24858_, _02210_);
  nor (_24860_, _24859_, _24856_);
  and (_24861_, _24860_, _03061_);
  and (_24862_, _10792_, _03805_);
  nor (_24863_, _24862_, _24814_);
  nor (_24864_, _24863_, _03061_);
  or (_24865_, _24864_, _24861_);
  and (_24867_, _24865_, _02208_);
  or (_24868_, _24853_, _02208_);
  nor (_24869_, _24868_, _24815_);
  nor (_24870_, _24869_, _24867_);
  nor (_24871_, _24870_, _02342_);
  and (_24872_, _10791_, _03805_);
  or (_24873_, _24872_, _24814_);
  and (_24874_, _24873_, _02342_);
  or (_24875_, _24874_, _24871_);
  and (_24876_, _24875_, _04953_);
  nor (_24878_, _10913_, _09281_);
  nor (_24879_, _24878_, _24814_);
  nor (_24880_, _24879_, _04953_);
  or (_24881_, _24880_, _24876_);
  and (_24882_, _24881_, _04958_);
  nor (_24883_, _10789_, _09281_);
  nor (_24884_, _24883_, _24814_);
  nor (_24885_, _24884_, _04958_);
  nor (_24886_, _24885_, _15890_);
  not (_24887_, _24886_);
  nor (_24889_, _24887_, _24882_);
  nor (_24890_, _24889_, _24817_);
  or (_24891_, _24890_, _39633_);
  or (_24892_, _39632_, \oc8051_golden_model_1.SBUF [0]);
  and (_24893_, _24892_, _39026_);
  and (_41716_, _24893_, _24891_);
  nor (_24894_, _03805_, \oc8051_golden_model_1.SBUF [1]);
  not (_24895_, _24894_);
  nor (_24896_, _10988_, _09281_);
  nor (_24897_, _24896_, _02208_);
  and (_24898_, _24897_, _24895_);
  nor (_24899_, _11113_, _09281_);
  nor (_24900_, _24899_, _03061_);
  and (_24901_, _24900_, _24895_);
  and (_24902_, _05075_, _03805_);
  not (_24903_, \oc8051_golden_model_1.SBUF [1]);
  nor (_24904_, _03805_, _24903_);
  nor (_24905_, _24904_, _02032_);
  not (_24906_, _24905_);
  nor (_24907_, _24906_, _24902_);
  not (_24909_, _24907_);
  nor (_24910_, _09281_, _03161_);
  nor (_24911_, _24910_, _24904_);
  and (_24912_, _24911_, _06188_);
  and (_24913_, _03805_, _01804_);
  nor (_24914_, _24913_, _24894_);
  and (_24915_, _24914_, _02062_);
  nor (_24916_, _02062_, _24903_);
  or (_24917_, _24916_, _24915_);
  and (_24918_, _24917_, _03006_);
  and (_24920_, _11001_, _03805_);
  nor (_24921_, _24920_, _24894_);
  and (_24922_, _24921_, _02158_);
  or (_24923_, _24922_, _24918_);
  and (_24924_, _24923_, _02519_);
  nor (_24925_, _24911_, _02519_);
  nor (_24926_, _24925_, _24924_);
  nor (_24927_, _24926_, _02153_);
  and (_24928_, _24914_, _02153_);
  nor (_24929_, _24928_, _06188_);
  not (_24931_, _24929_);
  nor (_24932_, _24931_, _24927_);
  nor (_24933_, _24932_, _24912_);
  nor (_24934_, _24933_, _02031_);
  nor (_24935_, _24934_, _01765_);
  and (_24936_, _24935_, _24909_);
  and (_24937_, _11096_, _03805_);
  nor (_24938_, _24937_, _02037_);
  and (_24939_, _24938_, _24895_);
  nor (_24940_, _24939_, _24936_);
  nor (_24941_, _24940_, _07629_);
  nor (_24942_, _10989_, _09281_);
  nor (_24943_, _24942_, _03059_);
  and (_24944_, _03805_, _02893_);
  nor (_24945_, _24944_, _01995_);
  or (_24946_, _24945_, _24943_);
  and (_24947_, _24946_, _24895_);
  nor (_24948_, _24947_, _24941_);
  nor (_24949_, _24948_, _02331_);
  nor (_24950_, _24949_, _24901_);
  nor (_24952_, _24950_, _02206_);
  nor (_24953_, _24952_, _24898_);
  nor (_24954_, _24953_, _02342_);
  nor (_24955_, _24904_, _04209_);
  nor (_24956_, _24955_, _03065_);
  and (_24957_, _24956_, _24914_);
  nor (_24958_, _24957_, _24954_);
  or (_24959_, _24958_, _17216_);
  nand (_24960_, _24913_, _04208_);
  nor (_24961_, _24894_, _04958_);
  and (_24963_, _24961_, _24960_);
  nor (_24964_, _24963_, _02366_);
  and (_24965_, _24944_, _04208_);
  or (_24966_, _24894_, _04953_);
  or (_24967_, _24966_, _24965_);
  and (_24968_, _24967_, _24964_);
  and (_24969_, _24968_, _24959_);
  nor (_24970_, _24921_, _02778_);
  nor (_24971_, _24970_, _24969_);
  nor (_24972_, _24971_, _02081_);
  nor (_24974_, _24920_, _24904_);
  and (_24975_, _24974_, _02081_);
  nor (_24976_, _24975_, _24972_);
  or (_24977_, _24976_, _39633_);
  or (_24978_, _39632_, \oc8051_golden_model_1.SBUF [1]);
  and (_24979_, _24978_, _39026_);
  and (_41717_, _24979_, _24977_);
  not (_24980_, \oc8051_golden_model_1.SBUF [2]);
  nor (_24981_, _03805_, _24980_);
  nor (_24982_, _11314_, _09281_);
  nor (_24983_, _24982_, _24981_);
  nor (_24984_, _24983_, _04958_);
  and (_24985_, _11315_, _03805_);
  nor (_24986_, _24985_, _24981_);
  nor (_24987_, _24986_, _03061_);
  and (_24988_, _03805_, _04866_);
  nor (_24989_, _24988_, _24981_);
  and (_24990_, _24989_, _01994_);
  and (_24991_, _03805_, \oc8051_golden_model_1.ACC [2]);
  nor (_24992_, _24991_, _24981_);
  nor (_24994_, _24992_, _02549_);
  nor (_24995_, _24992_, _02063_);
  nor (_24996_, _02062_, _24980_);
  or (_24997_, _24996_, _24995_);
  and (_24998_, _24997_, _03006_);
  nor (_24999_, _11199_, _09281_);
  nor (_25000_, _24999_, _24981_);
  nor (_25001_, _25000_, _03006_);
  or (_25002_, _25001_, _24998_);
  and (_25003_, _25002_, _02519_);
  nor (_25005_, _09281_, _03624_);
  nor (_25006_, _25005_, _24981_);
  nor (_25007_, _25006_, _02519_);
  nor (_25008_, _25007_, _25003_);
  nor (_25009_, _25008_, _02153_);
  or (_25010_, _25009_, _06188_);
  nor (_25011_, _25010_, _24994_);
  and (_25012_, _25006_, _06188_);
  nor (_25013_, _25012_, _25011_);
  nor (_25014_, _25013_, _02031_);
  and (_25016_, _05211_, _03805_);
  nor (_25017_, _24981_, _02032_);
  not (_25018_, _25017_);
  nor (_25019_, _25018_, _25016_);
  or (_25020_, _25019_, _01765_);
  nor (_25021_, _25020_, _25014_);
  nor (_25022_, _11298_, _09281_);
  nor (_25023_, _25022_, _24981_);
  nor (_25024_, _25023_, _02037_);
  or (_25025_, _25024_, _01994_);
  nor (_25026_, _25025_, _25021_);
  nor (_25027_, _25026_, _24990_);
  or (_25028_, _25027_, _02210_);
  and (_25029_, _11189_, _03805_);
  or (_25030_, _25029_, _24981_);
  or (_25031_, _25030_, _03059_);
  and (_25032_, _25031_, _03061_);
  and (_25033_, _25032_, _25028_);
  nor (_25034_, _25033_, _24987_);
  nor (_25035_, _25034_, _02206_);
  nor (_25037_, _24981_, _04309_);
  not (_25038_, _25037_);
  nor (_25039_, _24989_, _02208_);
  and (_25040_, _25039_, _25038_);
  nor (_25041_, _25040_, _25035_);
  nor (_25042_, _25041_, _02342_);
  or (_25043_, _25037_, _03065_);
  nor (_25044_, _25043_, _24992_);
  or (_25045_, _25044_, _02202_);
  nor (_25046_, _25045_, _25042_);
  nor (_25048_, _11187_, _09281_);
  or (_25049_, _24981_, _04953_);
  nor (_25050_, _25049_, _25048_);
  or (_25051_, _25050_, _02334_);
  nor (_25052_, _25051_, _25046_);
  nor (_25053_, _25052_, _24984_);
  nor (_25054_, _25053_, _02366_);
  nor (_25055_, _25000_, _02778_);
  or (_25056_, _25055_, _02081_);
  nor (_25057_, _25056_, _25054_);
  and (_25059_, _11367_, _03805_);
  nor (_25060_, _25059_, _24981_);
  and (_25061_, _25060_, _02081_);
  nor (_25062_, _25061_, _25057_);
  or (_25063_, _25062_, _39633_);
  or (_25064_, _39632_, \oc8051_golden_model_1.SBUF [2]);
  and (_25065_, _25064_, _39026_);
  and (_41719_, _25065_, _25063_);
  not (_25066_, \oc8051_golden_model_1.SBUF [3]);
  nor (_25067_, _03805_, _25066_);
  nor (_25068_, _11510_, _09281_);
  nor (_25069_, _25068_, _25067_);
  nor (_25070_, _25069_, _04958_);
  nor (_25071_, _25067_, _04153_);
  not (_25072_, _25071_);
  and (_25073_, _03805_, _04719_);
  nor (_25074_, _25073_, _25067_);
  nor (_25075_, _25074_, _02208_);
  and (_25076_, _25075_, _25072_);
  and (_25077_, _11511_, _03805_);
  nor (_25079_, _25077_, _25067_);
  nor (_25080_, _25079_, _03061_);
  nor (_25081_, _09281_, _03434_);
  nor (_25082_, _25081_, _25067_);
  and (_25083_, _25082_, _06188_);
  and (_25084_, _03805_, \oc8051_golden_model_1.ACC [3]);
  nor (_25085_, _25084_, _25067_);
  nor (_25086_, _25085_, _02063_);
  nor (_25087_, _02062_, _25066_);
  or (_25088_, _25087_, _25086_);
  and (_25090_, _25088_, _03006_);
  nor (_25091_, _11394_, _09281_);
  nor (_25092_, _25091_, _25067_);
  nor (_25093_, _25092_, _03006_);
  or (_25094_, _25093_, _25090_);
  and (_25095_, _25094_, _02519_);
  nor (_25096_, _25082_, _02519_);
  nor (_25097_, _25096_, _25095_);
  nor (_25098_, _25097_, _02153_);
  nor (_25099_, _25085_, _02549_);
  nor (_25101_, _25099_, _06188_);
  not (_25102_, _25101_);
  nor (_25103_, _25102_, _25098_);
  nor (_25104_, _25103_, _25083_);
  nor (_25105_, _25104_, _02031_);
  and (_25106_, _05166_, _03805_);
  nor (_25107_, _25067_, _02032_);
  not (_25108_, _25107_);
  nor (_25109_, _25108_, _25106_);
  nor (_25110_, _25109_, _01765_);
  not (_25111_, _25110_);
  nor (_25112_, _25111_, _25105_);
  nor (_25113_, _11490_, _09281_);
  nor (_25114_, _25113_, _25067_);
  nor (_25115_, _25114_, _02037_);
  or (_25116_, _25115_, _07629_);
  or (_25117_, _25116_, _25112_);
  and (_25118_, _11505_, _03805_);
  or (_25119_, _25067_, _03059_);
  or (_25120_, _25119_, _25118_);
  and (_25122_, _25074_, _01994_);
  nor (_25123_, _25122_, _02331_);
  and (_25124_, _25123_, _25120_);
  and (_25125_, _25124_, _25117_);
  nor (_25126_, _25125_, _25080_);
  nor (_25127_, _25126_, _02206_);
  nor (_25128_, _25127_, _25076_);
  nor (_25129_, _25128_, _02342_);
  or (_25130_, _25071_, _03065_);
  nor (_25131_, _25130_, _25085_);
  or (_25133_, _25131_, _02202_);
  nor (_25134_, _25133_, _25129_);
  nor (_25135_, _11503_, _09281_);
  or (_25136_, _25067_, _04953_);
  nor (_25137_, _25136_, _25135_);
  or (_25138_, _25137_, _02334_);
  nor (_25139_, _25138_, _25134_);
  nor (_25140_, _25139_, _25070_);
  nor (_25141_, _25140_, _02366_);
  nor (_25142_, _25092_, _02778_);
  or (_25144_, _25142_, _02081_);
  nor (_25145_, _25144_, _25141_);
  and (_25146_, _11567_, _03805_);
  nor (_25147_, _25146_, _25067_);
  and (_25148_, _25147_, _02081_);
  nor (_25149_, _25148_, _25145_);
  or (_25150_, _25149_, _39633_);
  or (_25151_, _39632_, \oc8051_golden_model_1.SBUF [3]);
  and (_25152_, _25151_, _39026_);
  and (_41720_, _25152_, _25150_);
  not (_25153_, \oc8051_golden_model_1.SBUF [4]);
  nor (_25154_, _03805_, _25153_);
  nor (_25155_, _11587_, _09281_);
  nor (_25156_, _25155_, _25154_);
  nor (_25157_, _25156_, _04958_);
  and (_25158_, _11588_, _03805_);
  nor (_25159_, _25158_, _25154_);
  nor (_25160_, _25159_, _03061_);
  and (_25161_, _05303_, _03805_);
  or (_25162_, _25161_, _25154_);
  and (_25164_, _25162_, _02031_);
  and (_25165_, _03805_, \oc8051_golden_model_1.ACC [4]);
  nor (_25166_, _25165_, _25154_);
  nor (_25167_, _25166_, _02549_);
  nor (_25168_, _25166_, _02063_);
  nor (_25169_, _02062_, _25153_);
  or (_25170_, _25169_, _25168_);
  and (_25171_, _25170_, _03006_);
  nor (_25172_, _11611_, _09281_);
  nor (_25173_, _25172_, _25154_);
  nor (_25175_, _25173_, _03006_);
  or (_25176_, _25175_, _25171_);
  and (_25177_, _25176_, _02519_);
  nor (_25178_, _04372_, _09281_);
  nor (_25179_, _25178_, _25154_);
  nor (_25180_, _25179_, _02519_);
  nor (_25181_, _25180_, _25177_);
  nor (_25182_, _25181_, _02153_);
  or (_25183_, _25182_, _06188_);
  nor (_25184_, _25183_, _25167_);
  and (_25186_, _25179_, _06188_);
  or (_25187_, _25186_, _02031_);
  nor (_25188_, _25187_, _25184_);
  or (_25189_, _25188_, _25164_);
  and (_25190_, _25189_, _02037_);
  nor (_25191_, _11704_, _09281_);
  nor (_25192_, _25191_, _25154_);
  nor (_25193_, _25192_, _02037_);
  or (_25194_, _25193_, _07629_);
  or (_25195_, _25194_, _25190_);
  and (_25197_, _11592_, _03805_);
  or (_25198_, _25154_, _03059_);
  or (_25199_, _25198_, _25197_);
  and (_25200_, _04831_, _03805_);
  nor (_25201_, _25200_, _25154_);
  and (_25202_, _25201_, _01994_);
  nor (_25203_, _25202_, _02331_);
  and (_25204_, _25203_, _25199_);
  and (_25205_, _25204_, _25195_);
  nor (_25206_, _25205_, _25160_);
  nor (_25208_, _25206_, _02206_);
  nor (_25209_, _25154_, _04420_);
  not (_25210_, _25209_);
  nor (_25211_, _25201_, _02208_);
  and (_25212_, _25211_, _25210_);
  nor (_25213_, _25212_, _25208_);
  nor (_25214_, _25213_, _02342_);
  or (_25215_, _25209_, _03065_);
  nor (_25216_, _25215_, _25166_);
  or (_25217_, _25216_, _02202_);
  nor (_25219_, _25217_, _25214_);
  nor (_25220_, _11590_, _09281_);
  or (_25221_, _25154_, _04953_);
  nor (_25222_, _25221_, _25220_);
  or (_25223_, _25222_, _02334_);
  nor (_25224_, _25223_, _25219_);
  nor (_25225_, _25224_, _25157_);
  nor (_25226_, _25225_, _02366_);
  nor (_25227_, _25173_, _02778_);
  or (_25228_, _25227_, _02081_);
  nor (_25230_, _25228_, _25226_);
  and (_25231_, _11771_, _03805_);
  nor (_25232_, _25231_, _25154_);
  and (_25233_, _25232_, _02081_);
  nor (_25234_, _25233_, _25230_);
  or (_25235_, _25234_, _39633_);
  or (_25236_, _39632_, \oc8051_golden_model_1.SBUF [4]);
  and (_25237_, _25236_, _39026_);
  and (_41721_, _25237_, _25235_);
  not (_25238_, \oc8051_golden_model_1.SBUF [5]);
  nor (_25240_, _03805_, _25238_);
  nor (_25241_, _11785_, _09281_);
  nor (_25242_, _25241_, _25240_);
  nor (_25243_, _25242_, _04958_);
  and (_25244_, _11786_, _03805_);
  nor (_25245_, _25244_, _25240_);
  nor (_25246_, _25245_, _03061_);
  and (_25247_, _04827_, _03805_);
  nor (_25248_, _25247_, _25240_);
  and (_25249_, _25248_, _01994_);
  and (_25251_, _03805_, \oc8051_golden_model_1.ACC [5]);
  nor (_25252_, _25251_, _25240_);
  nor (_25253_, _25252_, _02549_);
  nor (_25254_, _25252_, _02063_);
  nor (_25255_, _02062_, _25238_);
  or (_25256_, _25255_, _25254_);
  and (_25257_, _25256_, _03006_);
  nor (_25258_, _11804_, _09281_);
  nor (_25259_, _25258_, _25240_);
  nor (_25260_, _25259_, _03006_);
  or (_25262_, _25260_, _25257_);
  and (_25263_, _25262_, _02519_);
  nor (_25264_, _04057_, _09281_);
  nor (_25265_, _25264_, _25240_);
  nor (_25266_, _25265_, _02519_);
  nor (_25267_, _25266_, _25263_);
  nor (_25268_, _25267_, _02153_);
  or (_25269_, _25268_, _06188_);
  nor (_25270_, _25269_, _25253_);
  and (_25271_, _25265_, _06188_);
  nor (_25273_, _25271_, _25270_);
  nor (_25274_, _25273_, _02031_);
  and (_25275_, _05258_, _03805_);
  nor (_25276_, _25240_, _02032_);
  not (_25277_, _25276_);
  nor (_25278_, _25277_, _25275_);
  or (_25279_, _25278_, _01765_);
  nor (_25280_, _25279_, _25274_);
  nor (_25281_, _11900_, _09281_);
  nor (_25282_, _25281_, _25240_);
  nor (_25284_, _25282_, _02037_);
  or (_25285_, _25284_, _01994_);
  nor (_25286_, _25285_, _25280_);
  nor (_25287_, _25286_, _25249_);
  or (_25288_, _25287_, _02210_);
  and (_25289_, _11915_, _03805_);
  or (_25290_, _25289_, _25240_);
  or (_25291_, _25290_, _03059_);
  and (_25292_, _25291_, _03061_);
  and (_25293_, _25292_, _25288_);
  nor (_25295_, _25293_, _25246_);
  nor (_25296_, _25295_, _02206_);
  nor (_25297_, _25240_, _04104_);
  not (_25298_, _25297_);
  nor (_25299_, _25248_, _02208_);
  and (_25300_, _25299_, _25298_);
  nor (_25301_, _25300_, _25296_);
  nor (_25302_, _25301_, _02342_);
  or (_25303_, _25297_, _03065_);
  nor (_25304_, _25303_, _25252_);
  or (_25306_, _25304_, _02202_);
  nor (_25307_, _25306_, _25302_);
  nor (_25308_, _11913_, _09281_);
  or (_25309_, _25240_, _04953_);
  nor (_25310_, _25309_, _25308_);
  or (_25311_, _25310_, _02334_);
  nor (_25312_, _25311_, _25307_);
  nor (_25313_, _25312_, _25243_);
  nor (_25314_, _25313_, _02366_);
  nor (_25315_, _25259_, _02778_);
  or (_25317_, _25315_, _02081_);
  nor (_25318_, _25317_, _25314_);
  and (_25319_, _11974_, _03805_);
  nor (_25320_, _25319_, _25240_);
  and (_25321_, _25320_, _02081_);
  nor (_25322_, _25321_, _25318_);
  or (_25323_, _25322_, _39633_);
  or (_25324_, _39632_, \oc8051_golden_model_1.SBUF [5]);
  and (_25325_, _25324_, _39026_);
  and (_41722_, _25325_, _25323_);
  not (_25327_, \oc8051_golden_model_1.SBUF [6]);
  nor (_25328_, _03805_, _25327_);
  nor (_25329_, _12117_, _09281_);
  nor (_25330_, _25329_, _25328_);
  nor (_25331_, _25330_, _04958_);
  and (_25332_, _12118_, _03805_);
  nor (_25333_, _25332_, _25328_);
  nor (_25334_, _25333_, _03061_);
  and (_25335_, _12103_, _03805_);
  nor (_25336_, _25335_, _25328_);
  and (_25338_, _25336_, _01994_);
  nor (_25339_, _03964_, _09281_);
  nor (_25340_, _25339_, _25328_);
  and (_25341_, _25340_, _06188_);
  and (_25342_, _03805_, \oc8051_golden_model_1.ACC [6]);
  nor (_25343_, _25342_, _25328_);
  nor (_25344_, _25343_, _02549_);
  nor (_25345_, _25343_, _02063_);
  nor (_25346_, _02062_, _25327_);
  or (_25347_, _25346_, _25345_);
  and (_25349_, _25347_, _03006_);
  nor (_25350_, _11993_, _09281_);
  nor (_25351_, _25350_, _25328_);
  nor (_25352_, _25351_, _03006_);
  or (_25353_, _25352_, _25349_);
  and (_25354_, _25353_, _02519_);
  nor (_25355_, _25340_, _02519_);
  nor (_25356_, _25355_, _25354_);
  nor (_25357_, _25356_, _02153_);
  or (_25358_, _25357_, _06188_);
  nor (_25360_, _25358_, _25344_);
  nor (_25361_, _25360_, _25341_);
  nor (_25362_, _25361_, _02031_);
  and (_25363_, _05029_, _03805_);
  nor (_25364_, _25328_, _02032_);
  not (_25365_, _25364_);
  nor (_25366_, _25365_, _25363_);
  or (_25367_, _25366_, _01765_);
  nor (_25368_, _25367_, _25362_);
  nor (_25369_, _12096_, _09281_);
  nor (_25371_, _25369_, _25328_);
  nor (_25372_, _25371_, _02037_);
  or (_25373_, _25372_, _01994_);
  nor (_25374_, _25373_, _25368_);
  nor (_25375_, _25374_, _25338_);
  or (_25376_, _25375_, _02210_);
  and (_25377_, _12112_, _03805_);
  or (_25378_, _25377_, _25328_);
  or (_25379_, _25378_, _03059_);
  and (_25380_, _25379_, _03061_);
  and (_25382_, _25380_, _25376_);
  nor (_25383_, _25382_, _25334_);
  nor (_25384_, _25383_, _02206_);
  nor (_25385_, _25328_, _04011_);
  not (_25386_, _25385_);
  nor (_25387_, _25336_, _02208_);
  and (_25388_, _25387_, _25386_);
  nor (_25389_, _25388_, _25384_);
  nor (_25390_, _25389_, _02342_);
  or (_25391_, _25385_, _03065_);
  nor (_25392_, _25391_, _25343_);
  or (_25393_, _25392_, _02202_);
  nor (_25394_, _25393_, _25390_);
  nor (_25395_, _12110_, _09281_);
  or (_25396_, _25328_, _04953_);
  nor (_25397_, _25396_, _25395_);
  or (_25398_, _25397_, _02334_);
  nor (_25399_, _25398_, _25394_);
  nor (_25400_, _25399_, _25331_);
  nor (_25401_, _25400_, _02366_);
  nor (_25403_, _25351_, _02778_);
  or (_25404_, _25403_, _02081_);
  nor (_25405_, _25404_, _25401_);
  and (_25406_, _12178_, _03805_);
  nor (_25407_, _25406_, _25328_);
  and (_25408_, _25407_, _02081_);
  nor (_25409_, _25408_, _25405_);
  or (_25410_, _25409_, _39633_);
  or (_25411_, _39632_, \oc8051_golden_model_1.SBUF [6]);
  and (_25412_, _25411_, _39026_);
  and (_41723_, _25412_, _25410_);
  not (_25414_, \oc8051_golden_model_1.SCON [0]);
  nor (_25415_, _03868_, _25414_);
  and (_25416_, _10792_, _03868_);
  nor (_25417_, _25416_, _25415_);
  nor (_25418_, _25417_, _03061_);
  and (_25419_, _03868_, _04837_);
  nor (_25420_, _25419_, _25415_);
  and (_25421_, _25420_, _01994_);
  and (_25422_, _03868_, _03002_);
  nor (_25424_, _25422_, _25415_);
  and (_25425_, _25424_, _06188_);
  and (_25426_, _03868_, \oc8051_golden_model_1.ACC [0]);
  nor (_25427_, _25426_, _25415_);
  nor (_25428_, _25427_, _02063_);
  nor (_25429_, _02062_, _25414_);
  or (_25430_, _25429_, _25428_);
  and (_25431_, _25430_, _03006_);
  nor (_25432_, _04257_, _09360_);
  nor (_25433_, _25432_, _25415_);
  nor (_25435_, _25433_, _03006_);
  or (_25436_, _25435_, _25431_);
  and (_25437_, _25436_, _02058_);
  nor (_25438_, _04471_, _25414_);
  and (_25439_, _10814_, _04471_);
  nor (_25440_, _25439_, _25438_);
  nor (_25441_, _25440_, _02058_);
  nor (_25442_, _25441_, _25437_);
  nor (_25443_, _25442_, _02155_);
  nor (_25444_, _25424_, _02519_);
  or (_25446_, _25444_, _25443_);
  and (_25447_, _25446_, _02549_);
  nor (_25448_, _25427_, _02549_);
  or (_25449_, _25448_, _25447_);
  and (_25450_, _25449_, _02054_);
  and (_25451_, _25415_, _02053_);
  or (_25452_, _25451_, _25450_);
  and (_25453_, _25452_, _02047_);
  nor (_25454_, _25433_, _02047_);
  or (_25455_, _25454_, _25453_);
  and (_25457_, _25455_, _02043_);
  nor (_25458_, _10798_, _09397_);
  nor (_25459_, _25458_, _25438_);
  nor (_25460_, _25459_, _02043_);
  or (_25461_, _25460_, _06188_);
  nor (_25462_, _25461_, _25457_);
  nor (_25463_, _25462_, _25425_);
  nor (_25464_, _25463_, _02031_);
  and (_25465_, _05120_, _03868_);
  nor (_25466_, _25415_, _02032_);
  not (_25468_, _25466_);
  nor (_25469_, _25468_, _25465_);
  or (_25470_, _25469_, _01765_);
  nor (_25471_, _25470_, _25464_);
  nor (_25472_, _10898_, _09360_);
  nor (_25473_, _25472_, _25415_);
  nor (_25474_, _25473_, _02037_);
  or (_25475_, _25474_, _01994_);
  nor (_25476_, _25475_, _25471_);
  nor (_25477_, _25476_, _25421_);
  or (_25479_, _25477_, _02210_);
  and (_25480_, _10914_, _03868_);
  or (_25481_, _25480_, _25415_);
  or (_25482_, _25481_, _03059_);
  and (_25483_, _25482_, _03061_);
  and (_25484_, _25483_, _25479_);
  nor (_25485_, _25484_, _25418_);
  nor (_25486_, _25485_, _02206_);
  or (_25487_, _25420_, _02208_);
  nor (_25488_, _25487_, _25432_);
  nor (_25489_, _25488_, _25486_);
  nor (_25490_, _25489_, _02342_);
  nor (_25491_, _25415_, _04257_);
  or (_25492_, _25491_, _03065_);
  nor (_25493_, _25492_, _25427_);
  or (_25494_, _25493_, _02202_);
  nor (_25495_, _25494_, _25490_);
  nor (_25496_, _10913_, _09360_);
  or (_25497_, _25415_, _04953_);
  nor (_25498_, _25497_, _25496_);
  or (_25500_, _25498_, _02334_);
  nor (_25501_, _25500_, _25495_);
  nor (_25502_, _10789_, _09360_);
  nor (_25503_, _25502_, _25415_);
  nor (_25504_, _25503_, _04958_);
  or (_25505_, _25504_, _25501_);
  and (_25506_, _25505_, _02778_);
  nor (_25507_, _25433_, _02778_);
  or (_25508_, _25507_, _25506_);
  and (_25509_, _25508_, _01698_);
  and (_25511_, _25415_, _01697_);
  nor (_25512_, _25511_, _02081_);
  not (_25513_, _25512_);
  nor (_25514_, _25513_, _25509_);
  and (_25515_, _25433_, _02081_);
  or (_25516_, _25515_, _25514_);
  nand (_25517_, _25516_, _39632_);
  or (_25518_, _39632_, \oc8051_golden_model_1.SCON [0]);
  and (_25519_, _25518_, _39026_);
  and (_41725_, _25519_, _25517_);
  not (_25521_, \oc8051_golden_model_1.SCON [1]);
  nor (_25522_, _03868_, _25521_);
  and (_25523_, _05075_, _03868_);
  or (_25524_, _25523_, _25522_);
  and (_25525_, _25524_, _02031_);
  nor (_25526_, _03868_, \oc8051_golden_model_1.SCON [1]);
  and (_25527_, _03868_, _01804_);
  nor (_25528_, _25527_, _25526_);
  and (_25529_, _25528_, _02062_);
  nor (_25530_, _02062_, _25521_);
  or (_25532_, _25530_, _25529_);
  and (_25533_, _25532_, _03006_);
  and (_25534_, _11001_, _03868_);
  nor (_25535_, _25534_, _25526_);
  and (_25536_, _25535_, _02158_);
  or (_25537_, _25536_, _25533_);
  and (_25538_, _25537_, _02058_);
  nor (_25539_, _04471_, _25521_);
  and (_25540_, _11005_, _04471_);
  nor (_25541_, _25540_, _25539_);
  nor (_25543_, _25541_, _02058_);
  or (_25544_, _25543_, _25538_);
  and (_25545_, _25544_, _02519_);
  nor (_25546_, _09360_, _03161_);
  nor (_25547_, _25546_, _25522_);
  nor (_25548_, _25547_, _02519_);
  or (_25549_, _25548_, _25545_);
  nor (_25550_, _25549_, _02153_);
  nor (_25551_, _25528_, _02549_);
  or (_25552_, _25551_, _02053_);
  nor (_25554_, _25552_, _25550_);
  and (_25555_, _10992_, _04471_);
  nor (_25556_, _25555_, _25539_);
  nor (_25557_, _25556_, _02054_);
  or (_25558_, _25557_, _25554_);
  and (_25559_, _25558_, _02047_);
  nor (_25560_, _25539_, _11020_);
  nor (_25561_, _25560_, _25541_);
  and (_25562_, _25561_, _02046_);
  or (_25563_, _25562_, _25559_);
  and (_25565_, _25563_, _02043_);
  nor (_25566_, _11038_, _09397_);
  nor (_25567_, _25566_, _25539_);
  nor (_25568_, _25567_, _02043_);
  nor (_25569_, _25568_, _06188_);
  not (_25570_, _25569_);
  nor (_25571_, _25570_, _25565_);
  and (_25572_, _25547_, _06188_);
  or (_25573_, _25572_, _02031_);
  nor (_25574_, _25573_, _25571_);
  or (_25576_, _25574_, _25525_);
  and (_25577_, _25576_, _02037_);
  nor (_25578_, _11096_, _09360_);
  nor (_25579_, _25578_, _25522_);
  nor (_25580_, _25579_, _02037_);
  nor (_25581_, _25580_, _25577_);
  nor (_25582_, _25581_, _07629_);
  not (_25583_, _25526_);
  nor (_25584_, _10989_, _09360_);
  nor (_25585_, _25584_, _03059_);
  and (_25587_, _03868_, _02893_);
  nor (_25588_, _25587_, _01995_);
  or (_25589_, _25588_, _25585_);
  and (_25590_, _25589_, _25583_);
  nor (_25591_, _25590_, _25582_);
  nor (_25592_, _25591_, _02331_);
  nor (_25593_, _11113_, _09360_);
  nor (_25594_, _25593_, _03061_);
  and (_25595_, _25594_, _25583_);
  nor (_25596_, _25595_, _25592_);
  nor (_25598_, _25596_, _02206_);
  nor (_25599_, _10988_, _09360_);
  nor (_25600_, _25599_, _02208_);
  and (_25601_, _25600_, _25583_);
  nor (_25602_, _25601_, _25598_);
  nor (_25603_, _25602_, _02342_);
  nor (_25604_, _25522_, _04209_);
  nor (_25605_, _25604_, _03065_);
  and (_25606_, _25605_, _25528_);
  nor (_25607_, _25606_, _25603_);
  or (_25609_, _25607_, _17216_);
  nand (_25610_, _25527_, _04208_);
  nor (_25611_, _25526_, _04958_);
  and (_25612_, _25611_, _25610_);
  nor (_25613_, _25612_, _02366_);
  and (_25614_, _25587_, _04208_);
  or (_25615_, _25526_, _04953_);
  or (_25616_, _25615_, _25614_);
  and (_25617_, _25616_, _25613_);
  and (_25618_, _25617_, _25609_);
  nor (_25620_, _25535_, _02778_);
  or (_25621_, _25620_, _01697_);
  nor (_25622_, _25621_, _25618_);
  nor (_25623_, _25556_, _01698_);
  or (_25624_, _25623_, _02081_);
  nor (_25625_, _25624_, _25622_);
  nor (_25626_, _25534_, _25522_);
  and (_25627_, _25626_, _02081_);
  nor (_25628_, _25627_, _25625_);
  or (_25629_, _25628_, _39633_);
  or (_25630_, _39632_, \oc8051_golden_model_1.SCON [1]);
  and (_25631_, _25630_, _39026_);
  and (_41726_, _25631_, _25629_);
  not (_25632_, \oc8051_golden_model_1.SCON [2]);
  nor (_25633_, _03868_, _25632_);
  and (_25634_, _03868_, _04866_);
  nor (_25635_, _25634_, _25633_);
  and (_25636_, _25635_, _01994_);
  nor (_25637_, _09360_, _03624_);
  nor (_25638_, _25637_, _25633_);
  and (_25640_, _25638_, _06188_);
  and (_25641_, _03868_, \oc8051_golden_model_1.ACC [2]);
  nor (_25642_, _25641_, _25633_);
  nor (_25643_, _25642_, _02063_);
  nor (_25644_, _02062_, _25632_);
  or (_25645_, _25644_, _25643_);
  and (_25646_, _25645_, _03006_);
  nor (_25647_, _11199_, _09360_);
  nor (_25648_, _25647_, _25633_);
  nor (_25649_, _25648_, _03006_);
  or (_25651_, _25649_, _25646_);
  and (_25652_, _25651_, _02058_);
  nor (_25653_, _04471_, _25632_);
  and (_25654_, _11194_, _04471_);
  nor (_25655_, _25654_, _25653_);
  nor (_25656_, _25655_, _02058_);
  or (_25657_, _25656_, _02155_);
  or (_25658_, _25657_, _25652_);
  nand (_25659_, _25638_, _02155_);
  and (_25660_, _25659_, _25658_);
  and (_25662_, _25660_, _02549_);
  nor (_25663_, _25642_, _02549_);
  or (_25664_, _25663_, _25662_);
  and (_25665_, _25664_, _02054_);
  and (_25666_, _11192_, _04471_);
  nor (_25667_, _25666_, _25653_);
  nor (_25668_, _25667_, _02054_);
  or (_25669_, _25668_, _25665_);
  and (_25670_, _25669_, _02047_);
  nor (_25671_, _25653_, _11223_);
  nor (_25673_, _25671_, _25655_);
  and (_25674_, _25673_, _02046_);
  or (_25675_, _25674_, _25670_);
  and (_25676_, _25675_, _02043_);
  nor (_25677_, _11241_, _09397_);
  nor (_25678_, _25677_, _25653_);
  nor (_25679_, _25678_, _02043_);
  nor (_25680_, _25679_, _06188_);
  not (_25681_, _25680_);
  nor (_25682_, _25681_, _25676_);
  nor (_25684_, _25682_, _25640_);
  nor (_25685_, _25684_, _02031_);
  and (_25686_, _05211_, _03868_);
  nor (_25687_, _25633_, _02032_);
  not (_25688_, _25687_);
  nor (_25689_, _25688_, _25686_);
  or (_25690_, _25689_, _01765_);
  nor (_25691_, _25690_, _25685_);
  nor (_25692_, _11298_, _09360_);
  nor (_25693_, _25633_, _25692_);
  nor (_25695_, _25693_, _02037_);
  or (_25696_, _25695_, _01994_);
  nor (_25697_, _25696_, _25691_);
  nor (_25698_, _25697_, _25636_);
  or (_25699_, _25698_, _02210_);
  and (_25700_, _11189_, _03868_);
  or (_25701_, _25700_, _25633_);
  or (_25702_, _25701_, _03059_);
  and (_25703_, _25702_, _03061_);
  and (_25704_, _25703_, _25699_);
  and (_25706_, _11315_, _03868_);
  nor (_25707_, _25706_, _25633_);
  nor (_25708_, _25707_, _03061_);
  nor (_25709_, _25708_, _25704_);
  nor (_25710_, _25709_, _02206_);
  nor (_25711_, _25633_, _04309_);
  not (_25712_, _25711_);
  nor (_25713_, _25635_, _02208_);
  and (_25714_, _25713_, _25712_);
  nor (_25715_, _25714_, _25710_);
  nor (_25716_, _25715_, _02342_);
  or (_25717_, _25711_, _03065_);
  nor (_25718_, _25717_, _25642_);
  or (_25719_, _25718_, _02202_);
  nor (_25720_, _25719_, _25716_);
  nor (_25721_, _11187_, _09360_);
  or (_25722_, _25633_, _04953_);
  nor (_25723_, _25722_, _25721_);
  or (_25724_, _25723_, _02334_);
  nor (_25725_, _25724_, _25720_);
  nor (_25727_, _11314_, _09360_);
  nor (_25728_, _25727_, _25633_);
  nor (_25729_, _25728_, _04958_);
  or (_25730_, _25729_, _25725_);
  and (_25731_, _25730_, _02778_);
  nor (_25732_, _25648_, _02778_);
  or (_25733_, _25732_, _25731_);
  and (_25734_, _25733_, _01698_);
  nor (_25735_, _25667_, _01698_);
  or (_25736_, _25735_, _25734_);
  and (_25738_, _25736_, _02082_);
  and (_25739_, _11367_, _03868_);
  nor (_25740_, _25739_, _25633_);
  nor (_25741_, _25740_, _02082_);
  or (_25742_, _25741_, _25738_);
  or (_25743_, _25742_, _39633_);
  or (_25744_, _39632_, \oc8051_golden_model_1.SCON [2]);
  and (_25745_, _25744_, _39026_);
  and (_41727_, _25745_, _25743_);
  not (_25746_, \oc8051_golden_model_1.SCON [3]);
  nor (_25748_, _03868_, _25746_);
  and (_25749_, _03868_, _04719_);
  nor (_25750_, _25749_, _25748_);
  and (_25751_, _25750_, _01994_);
  nor (_25752_, _09360_, _03434_);
  nor (_25753_, _25752_, _25748_);
  and (_25754_, _25753_, _06188_);
  and (_25755_, _03868_, \oc8051_golden_model_1.ACC [3]);
  nor (_25756_, _25755_, _25748_);
  nor (_25757_, _25756_, _02063_);
  nor (_25759_, _02062_, _25746_);
  or (_25760_, _25759_, _25757_);
  and (_25761_, _25760_, _03006_);
  nor (_25762_, _11394_, _09360_);
  nor (_25763_, _25762_, _25748_);
  nor (_25764_, _25763_, _03006_);
  or (_25765_, _25764_, _25761_);
  and (_25766_, _25765_, _02058_);
  nor (_25767_, _04471_, _25746_);
  and (_25768_, _11398_, _04471_);
  nor (_25770_, _25768_, _25767_);
  nor (_25771_, _25770_, _02058_);
  or (_25772_, _25771_, _25766_);
  and (_25773_, _25772_, _02519_);
  nor (_25774_, _25753_, _02519_);
  or (_25775_, _25774_, _25773_);
  and (_25776_, _25775_, _02549_);
  nor (_25777_, _25756_, _02549_);
  or (_25778_, _25777_, _25776_);
  and (_25779_, _25778_, _02054_);
  and (_25781_, _11408_, _04471_);
  nor (_25782_, _25781_, _25767_);
  nor (_25783_, _25782_, _02054_);
  or (_25784_, _25783_, _25779_);
  and (_25785_, _25784_, _02047_);
  nor (_25786_, _25767_, _11415_);
  nor (_25787_, _25786_, _25770_);
  and (_25788_, _25787_, _02046_);
  or (_25789_, _25788_, _25785_);
  and (_25790_, _25789_, _02043_);
  nor (_25792_, _11433_, _09397_);
  nor (_25793_, _25792_, _25767_);
  nor (_25794_, _25793_, _02043_);
  nor (_25795_, _25794_, _06188_);
  not (_25796_, _25795_);
  nor (_25797_, _25796_, _25790_);
  nor (_25798_, _25797_, _25754_);
  nor (_25799_, _25798_, _02031_);
  and (_25800_, _05166_, _03868_);
  nor (_25801_, _25748_, _02032_);
  not (_25802_, _25801_);
  nor (_25803_, _25802_, _25800_);
  or (_25804_, _25803_, _01765_);
  nor (_25805_, _25804_, _25799_);
  nor (_25806_, _11490_, _09360_);
  nor (_25807_, _25748_, _25806_);
  nor (_25808_, _25807_, _02037_);
  or (_25809_, _25808_, _01994_);
  nor (_25810_, _25809_, _25805_);
  nor (_25811_, _25810_, _25751_);
  or (_25813_, _25811_, _02210_);
  and (_25814_, _11505_, _03868_);
  or (_25815_, _25814_, _25748_);
  or (_25816_, _25815_, _03059_);
  and (_25817_, _25816_, _03061_);
  and (_25818_, _25817_, _25813_);
  and (_25819_, _11511_, _03868_);
  nor (_25820_, _25819_, _25748_);
  nor (_25821_, _25820_, _03061_);
  nor (_25822_, _25821_, _25818_);
  nor (_25824_, _25822_, _02206_);
  nor (_25825_, _25748_, _04153_);
  not (_25826_, _25825_);
  nor (_25827_, _25750_, _02208_);
  and (_25828_, _25827_, _25826_);
  nor (_25829_, _25828_, _25824_);
  nor (_25830_, _25829_, _02342_);
  or (_25831_, _25825_, _03065_);
  nor (_25832_, _25831_, _25756_);
  or (_25833_, _25832_, _02202_);
  nor (_25835_, _25833_, _25830_);
  nor (_25836_, _11503_, _09360_);
  or (_25837_, _25748_, _04953_);
  nor (_25838_, _25837_, _25836_);
  or (_25839_, _25838_, _02334_);
  nor (_25840_, _25839_, _25835_);
  nor (_25841_, _11510_, _09360_);
  nor (_25842_, _25841_, _25748_);
  nor (_25843_, _25842_, _04958_);
  or (_25844_, _25843_, _25840_);
  and (_25846_, _25844_, _02778_);
  nor (_25847_, _25763_, _02778_);
  or (_25848_, _25847_, _25846_);
  and (_25849_, _25848_, _01698_);
  nor (_25850_, _25782_, _01698_);
  nor (_25851_, _25850_, _02081_);
  not (_25852_, _25851_);
  nor (_25853_, _25852_, _25849_);
  and (_25854_, _11567_, _03868_);
  nor (_25855_, _25854_, _25748_);
  and (_25857_, _25855_, _02081_);
  nor (_25858_, _25857_, _25853_);
  or (_25859_, _25858_, _39633_);
  or (_25860_, _39632_, \oc8051_golden_model_1.SCON [3]);
  and (_25861_, _25860_, _39026_);
  and (_41728_, _25861_, _25859_);
  not (_25862_, \oc8051_golden_model_1.SCON [4]);
  nor (_25863_, _03868_, _25862_);
  and (_25864_, _04831_, _03868_);
  nor (_25865_, _25864_, _25863_);
  and (_25867_, _25865_, _01994_);
  nor (_25868_, _04372_, _09360_);
  nor (_25869_, _25868_, _25863_);
  and (_25870_, _25869_, _06188_);
  and (_25871_, _03868_, \oc8051_golden_model_1.ACC [4]);
  nor (_25872_, _25871_, _25863_);
  nor (_25873_, _25872_, _02063_);
  nor (_25874_, _02062_, _25862_);
  or (_25875_, _25874_, _25873_);
  and (_25876_, _25875_, _03006_);
  nor (_25878_, _11611_, _09360_);
  nor (_25879_, _25878_, _25863_);
  nor (_25880_, _25879_, _03006_);
  or (_25881_, _25880_, _25876_);
  and (_25882_, _25881_, _02058_);
  nor (_25883_, _04471_, _25862_);
  and (_25884_, _11597_, _04471_);
  nor (_25885_, _25884_, _25883_);
  nor (_25886_, _25885_, _02058_);
  or (_25887_, _25886_, _25882_);
  and (_25889_, _25887_, _02519_);
  nor (_25890_, _25869_, _02519_);
  or (_25891_, _25890_, _25889_);
  and (_25892_, _25891_, _02549_);
  nor (_25893_, _25872_, _02549_);
  or (_25894_, _25893_, _25892_);
  and (_25895_, _25894_, _02054_);
  and (_25896_, _11595_, _04471_);
  nor (_25897_, _25896_, _25883_);
  nor (_25898_, _25897_, _02054_);
  or (_25899_, _25898_, _25895_);
  and (_25900_, _25899_, _02047_);
  nor (_25901_, _25883_, _11628_);
  nor (_25902_, _25901_, _25885_);
  and (_25903_, _25902_, _02046_);
  or (_25904_, _25903_, _25900_);
  and (_25905_, _25904_, _02043_);
  nor (_25906_, _11646_, _09397_);
  nor (_25907_, _25906_, _25883_);
  nor (_25908_, _25907_, _02043_);
  nor (_25910_, _25908_, _06188_);
  not (_25911_, _25910_);
  nor (_25912_, _25911_, _25905_);
  nor (_25913_, _25912_, _25870_);
  nor (_25914_, _25913_, _02031_);
  and (_25915_, _05303_, _03868_);
  nor (_25916_, _25863_, _02032_);
  not (_25917_, _25916_);
  nor (_25918_, _25917_, _25915_);
  or (_25919_, _25918_, _01765_);
  nor (_25921_, _25919_, _25914_);
  nor (_25922_, _11704_, _09360_);
  nor (_25923_, _25863_, _25922_);
  nor (_25924_, _25923_, _02037_);
  or (_25925_, _25924_, _01994_);
  nor (_25926_, _25925_, _25921_);
  nor (_25927_, _25926_, _25867_);
  or (_25928_, _25927_, _02210_);
  and (_25929_, _11592_, _03868_);
  or (_25930_, _25929_, _25863_);
  or (_25932_, _25930_, _03059_);
  and (_25933_, _25932_, _03061_);
  and (_25934_, _25933_, _25928_);
  and (_25935_, _11588_, _03868_);
  nor (_25936_, _25935_, _25863_);
  nor (_25937_, _25936_, _03061_);
  nor (_25938_, _25937_, _25934_);
  nor (_25939_, _25938_, _02206_);
  nor (_25940_, _25863_, _04420_);
  not (_25941_, _25940_);
  nor (_25943_, _25865_, _02208_);
  and (_25944_, _25943_, _25941_);
  nor (_25945_, _25944_, _25939_);
  nor (_25946_, _25945_, _02342_);
  or (_25947_, _25940_, _03065_);
  nor (_25948_, _25947_, _25872_);
  or (_25949_, _25948_, _02202_);
  nor (_25950_, _25949_, _25946_);
  nor (_25951_, _11590_, _09360_);
  or (_25952_, _25863_, _04953_);
  nor (_25954_, _25952_, _25951_);
  or (_25955_, _25954_, _02334_);
  nor (_25956_, _25955_, _25950_);
  nor (_25957_, _11587_, _09360_);
  nor (_25958_, _25957_, _25863_);
  nor (_25959_, _25958_, _04958_);
  or (_25960_, _25959_, _25956_);
  and (_25961_, _25960_, _02778_);
  nor (_25962_, _25879_, _02778_);
  or (_25963_, _25962_, _25961_);
  and (_25965_, _25963_, _01698_);
  nor (_25966_, _25897_, _01698_);
  or (_25967_, _25966_, _25965_);
  and (_25968_, _25967_, _02082_);
  and (_25969_, _11771_, _03868_);
  nor (_25970_, _25969_, _25863_);
  nor (_25971_, _25970_, _02082_);
  or (_25972_, _25971_, _25968_);
  or (_25973_, _25972_, _39633_);
  or (_25974_, _39632_, \oc8051_golden_model_1.SCON [4]);
  and (_25976_, _25974_, _39026_);
  and (_41729_, _25976_, _25973_);
  not (_25977_, \oc8051_golden_model_1.SCON [5]);
  nor (_25978_, _03868_, _25977_);
  and (_25979_, _04827_, _03868_);
  nor (_25980_, _25979_, _25978_);
  and (_25981_, _25980_, _01994_);
  nor (_25982_, _04057_, _09360_);
  nor (_25983_, _25982_, _25978_);
  and (_25984_, _25983_, _06188_);
  and (_25986_, _03868_, \oc8051_golden_model_1.ACC [5]);
  nor (_25987_, _25986_, _25978_);
  nor (_25988_, _25987_, _02063_);
  nor (_25989_, _02062_, _25977_);
  or (_25990_, _25989_, _25988_);
  and (_25991_, _25990_, _03006_);
  nor (_25992_, _11804_, _09360_);
  nor (_25993_, _25992_, _25978_);
  nor (_25994_, _25993_, _03006_);
  or (_25995_, _25994_, _25991_);
  and (_25997_, _25995_, _02058_);
  nor (_25998_, _04471_, _25977_);
  and (_25999_, _11789_, _04471_);
  nor (_26000_, _25999_, _25998_);
  nor (_26001_, _26000_, _02058_);
  or (_26002_, _26001_, _25997_);
  and (_26003_, _26002_, _02519_);
  nor (_26004_, _25983_, _02519_);
  or (_26005_, _26004_, _26003_);
  and (_26006_, _26005_, _02549_);
  nor (_26008_, _25987_, _02549_);
  or (_26009_, _26008_, _26006_);
  and (_26010_, _26009_, _02054_);
  and (_26011_, _11816_, _04471_);
  nor (_26012_, _26011_, _25998_);
  nor (_26013_, _26012_, _02054_);
  or (_26014_, _26013_, _26010_);
  and (_26015_, _26014_, _02047_);
  nor (_26016_, _25998_, _11823_);
  nor (_26017_, _26016_, _26000_);
  and (_26019_, _26017_, _02046_);
  or (_26020_, _26019_, _26015_);
  and (_26021_, _26020_, _02043_);
  nor (_26022_, _11841_, _09397_);
  nor (_26023_, _26022_, _25998_);
  nor (_26024_, _26023_, _02043_);
  nor (_26025_, _26024_, _06188_);
  not (_26026_, _26025_);
  nor (_26027_, _26026_, _26021_);
  nor (_26028_, _26027_, _25984_);
  nor (_26030_, _26028_, _02031_);
  and (_26031_, _05258_, _03868_);
  nor (_26032_, _25978_, _02032_);
  not (_26033_, _26032_);
  nor (_26034_, _26033_, _26031_);
  or (_26035_, _26034_, _01765_);
  nor (_26036_, _26035_, _26030_);
  nor (_26037_, _11900_, _09360_);
  nor (_26038_, _26037_, _25978_);
  nor (_26039_, _26038_, _02037_);
  or (_26041_, _26039_, _01994_);
  nor (_26042_, _26041_, _26036_);
  nor (_26043_, _26042_, _25981_);
  or (_26044_, _26043_, _02210_);
  and (_26045_, _11915_, _03868_);
  or (_26046_, _26045_, _25978_);
  or (_26047_, _26046_, _03059_);
  and (_26048_, _26047_, _03061_);
  and (_26049_, _26048_, _26044_);
  and (_26050_, _11786_, _03868_);
  nor (_26051_, _26050_, _25978_);
  nor (_26052_, _26051_, _03061_);
  nor (_26053_, _26052_, _26049_);
  nor (_26054_, _26053_, _02206_);
  nor (_26055_, _25978_, _04104_);
  not (_26056_, _26055_);
  nor (_26057_, _25980_, _02208_);
  and (_26058_, _26057_, _26056_);
  nor (_26059_, _26058_, _26054_);
  nor (_26060_, _26059_, _02342_);
  or (_26062_, _26055_, _03065_);
  nor (_26063_, _26062_, _25987_);
  or (_26064_, _26063_, _02202_);
  nor (_26065_, _26064_, _26060_);
  nor (_26066_, _11913_, _09360_);
  or (_26067_, _25978_, _04953_);
  nor (_26068_, _26067_, _26066_);
  or (_26069_, _26068_, _02334_);
  nor (_26070_, _26069_, _26065_);
  nor (_26071_, _11785_, _09360_);
  nor (_26073_, _26071_, _25978_);
  nor (_26074_, _26073_, _04958_);
  or (_26075_, _26074_, _26070_);
  and (_26076_, _26075_, _02778_);
  nor (_26077_, _25993_, _02778_);
  or (_26078_, _26077_, _26076_);
  and (_26079_, _26078_, _01698_);
  nor (_26080_, _26012_, _01698_);
  or (_26081_, _26080_, _26079_);
  and (_26082_, _26081_, _02082_);
  and (_26084_, _11974_, _03868_);
  nor (_26085_, _26084_, _25978_);
  nor (_26086_, _26085_, _02082_);
  or (_26087_, _26086_, _26082_);
  or (_26088_, _26087_, _39633_);
  or (_26089_, _39632_, \oc8051_golden_model_1.SCON [5]);
  and (_26090_, _26089_, _39026_);
  and (_41730_, _26090_, _26088_);
  not (_26091_, \oc8051_golden_model_1.SCON [6]);
  nor (_26092_, _03868_, _26091_);
  and (_26094_, _12103_, _03868_);
  nor (_26095_, _26094_, _26092_);
  and (_26096_, _26095_, _01994_);
  nor (_26097_, _03964_, _09360_);
  nor (_26098_, _26097_, _26092_);
  and (_26099_, _26098_, _06188_);
  and (_26100_, _03868_, \oc8051_golden_model_1.ACC [6]);
  nor (_26101_, _26100_, _26092_);
  nor (_26102_, _26101_, _02063_);
  nor (_26103_, _02062_, _26091_);
  or (_26105_, _26103_, _26102_);
  and (_26106_, _26105_, _03006_);
  nor (_26107_, _11993_, _09360_);
  nor (_26108_, _26107_, _26092_);
  nor (_26109_, _26108_, _03006_);
  or (_26110_, _26109_, _26106_);
  and (_26111_, _26110_, _02058_);
  nor (_26112_, _04471_, _26091_);
  and (_26113_, _11990_, _04471_);
  nor (_26114_, _26113_, _26112_);
  nor (_26116_, _26114_, _02058_);
  or (_26117_, _26116_, _26111_);
  and (_26118_, _26117_, _02519_);
  nor (_26119_, _26098_, _02519_);
  or (_26120_, _26119_, _26118_);
  and (_26121_, _26120_, _02549_);
  nor (_26122_, _26101_, _02549_);
  or (_26123_, _26122_, _26121_);
  and (_26124_, _26123_, _02054_);
  and (_26125_, _12017_, _04471_);
  nor (_26127_, _26125_, _26112_);
  nor (_26128_, _26127_, _02054_);
  or (_26129_, _26128_, _26124_);
  and (_26130_, _26129_, _02047_);
  nor (_26131_, _26112_, _12024_);
  nor (_26132_, _26131_, _26114_);
  and (_26133_, _26132_, _02046_);
  or (_26134_, _26133_, _26130_);
  and (_26135_, _26134_, _02043_);
  nor (_26136_, _12042_, _09397_);
  nor (_26138_, _26136_, _26112_);
  nor (_26139_, _26138_, _02043_);
  nor (_26140_, _26139_, _06188_);
  not (_26141_, _26140_);
  nor (_26142_, _26141_, _26135_);
  nor (_26143_, _26142_, _26099_);
  nor (_26144_, _26143_, _02031_);
  and (_26145_, _05029_, _03868_);
  nor (_26146_, _26092_, _02032_);
  not (_26147_, _26146_);
  nor (_26149_, _26147_, _26145_);
  or (_26150_, _26149_, _01765_);
  nor (_26151_, _26150_, _26144_);
  nor (_26152_, _12096_, _09360_);
  nor (_26153_, _26152_, _26092_);
  nor (_26154_, _26153_, _02037_);
  or (_26155_, _26154_, _01994_);
  nor (_26156_, _26155_, _26151_);
  nor (_26157_, _26156_, _26096_);
  or (_26158_, _26157_, _02210_);
  and (_26160_, _12112_, _03868_);
  or (_26161_, _26160_, _26092_);
  or (_26162_, _26161_, _03059_);
  and (_26163_, _26162_, _03061_);
  and (_26164_, _26163_, _26158_);
  and (_26165_, _12118_, _03868_);
  nor (_26166_, _26165_, _26092_);
  nor (_26167_, _26166_, _03061_);
  nor (_26168_, _26167_, _26164_);
  nor (_26169_, _26168_, _02206_);
  nor (_26171_, _26092_, _04011_);
  not (_26172_, _26171_);
  nor (_26173_, _26095_, _02208_);
  and (_26174_, _26173_, _26172_);
  nor (_26175_, _26174_, _26169_);
  nor (_26176_, _26175_, _02342_);
  or (_26177_, _26171_, _03065_);
  nor (_26178_, _26177_, _26101_);
  or (_26179_, _26178_, _02202_);
  nor (_26180_, _26179_, _26176_);
  nor (_26182_, _12110_, _09360_);
  or (_26183_, _26092_, _04953_);
  nor (_26184_, _26183_, _26182_);
  or (_26185_, _26184_, _02334_);
  nor (_26186_, _26185_, _26180_);
  nor (_26187_, _12117_, _09360_);
  nor (_26188_, _26187_, _26092_);
  nor (_26189_, _26188_, _04958_);
  or (_26190_, _26189_, _26186_);
  and (_26191_, _26190_, _02778_);
  nor (_26193_, _26108_, _02778_);
  or (_26194_, _26193_, _26191_);
  and (_26195_, _26194_, _01698_);
  nor (_26196_, _26127_, _01698_);
  or (_26197_, _26196_, _26195_);
  and (_26198_, _26197_, _02082_);
  and (_26199_, _12178_, _03868_);
  nor (_26200_, _26199_, _26092_);
  nor (_26201_, _26200_, _02082_);
  or (_26202_, _26201_, _26198_);
  or (_26204_, _26202_, _39633_);
  or (_26205_, _39632_, \oc8051_golden_model_1.SCON [6]);
  and (_26206_, _26205_, _39026_);
  and (_41731_, _26206_, _26204_);
  nor (_26207_, _04182_, _01986_);
  nor (_26208_, _04257_, _09531_);
  nor (_26209_, _26208_, _26207_);
  and (_26210_, _26209_, _15890_);
  and (_26211_, _03893_, _04837_);
  nor (_26212_, _26211_, _26207_);
  nor (_26214_, _26212_, _02208_);
  not (_26215_, _26214_);
  nor (_26216_, _26215_, _26208_);
  and (_26217_, _03893_, \oc8051_golden_model_1.ACC [0]);
  nor (_26218_, _26217_, _26207_);
  nor (_26219_, _26218_, _02063_);
  nor (_26220_, _02062_, _01986_);
  or (_26221_, _26220_, _26219_);
  and (_26222_, _26221_, _03006_);
  nor (_26223_, _26209_, _03006_);
  or (_26225_, _26223_, _26222_);
  and (_26226_, _26225_, _02519_);
  or (_26227_, _26226_, _02587_);
  and (_26228_, _26227_, _02549_);
  nor (_26229_, _26218_, _02549_);
  or (_26230_, _26229_, _26228_);
  and (_26231_, _26230_, _03114_);
  nor (_26232_, _06188_, _03031_);
  not (_26233_, _26232_);
  nor (_26234_, _26233_, _26231_);
  or (_26236_, _09531_, _03020_);
  nor (_26237_, _26207_, _05444_);
  and (_26238_, _26237_, _26236_);
  nor (_26239_, _26238_, _26234_);
  nor (_26240_, _26239_, _02031_);
  nor (_26241_, _26207_, _02032_);
  nand (_26242_, _05120_, _04182_);
  and (_26243_, _26242_, _26241_);
  nor (_26244_, _26243_, _26240_);
  nor (_26245_, _26244_, _01765_);
  or (_26247_, _10898_, _09531_);
  nor (_26248_, _26207_, _02037_);
  and (_26249_, _26248_, _26247_);
  or (_26250_, _26249_, _01994_);
  nor (_26251_, _26250_, _26245_);
  nand (_26252_, _26212_, _03059_);
  and (_26253_, _26252_, _07629_);
  nor (_26254_, _26253_, _26251_);
  and (_26255_, _10914_, _03893_);
  nor (_26256_, _26255_, _26207_);
  and (_26258_, _26256_, _02210_);
  nor (_26259_, _26258_, _26254_);
  and (_26260_, _26259_, _03061_);
  and (_26261_, _10792_, _03893_);
  nor (_26262_, _26261_, _26207_);
  nor (_26263_, _26262_, _03061_);
  or (_26264_, _26263_, _26260_);
  and (_26265_, _26264_, _02208_);
  nor (_26266_, _26265_, _26216_);
  nor (_26267_, _26266_, _02342_);
  and (_26269_, _10791_, _03893_);
  or (_26270_, _26269_, _26207_);
  and (_26271_, _26270_, _02342_);
  or (_26272_, _26271_, _26267_);
  and (_26273_, _26272_, _04953_);
  nor (_26274_, _10913_, _09478_);
  nor (_26275_, _26274_, _26207_);
  nor (_26276_, _26275_, _04953_);
  or (_26277_, _26276_, _26273_);
  and (_26278_, _26277_, _04958_);
  nor (_26280_, _10789_, _09531_);
  nor (_26281_, _26280_, _26207_);
  nor (_26282_, _26281_, _04958_);
  nor (_26283_, _26282_, _15890_);
  not (_26284_, _26283_);
  nor (_26285_, _26284_, _26278_);
  nor (_26286_, _26285_, _26210_);
  and (_26287_, _26286_, _39632_);
  nor (_26288_, _39632_, _01986_);
  or (_26289_, _26288_, rst);
  or (_41733_, _26289_, _26287_);
  nor (_26291_, _04182_, _03104_);
  and (_26292_, _11001_, _04182_);
  nor (_26293_, _26292_, _26291_);
  nor (_26294_, _26293_, _02082_);
  nor (_26295_, _23146_, _03104_);
  and (_26296_, _11113_, _03893_);
  or (_26297_, _26296_, _26291_);
  and (_26298_, _26297_, _02331_);
  and (_26299_, _01718_, _03104_);
  and (_26301_, _03893_, \oc8051_golden_model_1.ACC [1]);
  or (_26302_, _26301_, _26291_);
  nor (_26303_, _26302_, _02063_);
  nor (_26304_, _09495_, \oc8051_golden_model_1.SP [1]);
  and (_26305_, _01747_, \oc8051_golden_model_1.SP [1]);
  nor (_26306_, _26305_, _26304_);
  nor (_26307_, _26306_, _26303_);
  and (_26308_, _26307_, _03006_);
  nor (_26309_, _04182_, \oc8051_golden_model_1.SP [1]);
  nor (_26310_, _26309_, _26292_);
  and (_26312_, _26310_, _02158_);
  or (_26313_, _26312_, _26308_);
  and (_26314_, _26313_, _01745_);
  nor (_26315_, _01745_, \oc8051_golden_model_1.SP [1]);
  or (_26316_, _26315_, _02155_);
  or (_26317_, _26316_, _26314_);
  nand (_26318_, _03108_, _02155_);
  and (_26319_, _26318_, _26317_);
  and (_26320_, _26319_, _02549_);
  and (_26321_, _26302_, _02153_);
  or (_26323_, _26321_, _26320_);
  and (_26324_, _26323_, _03114_);
  or (_26325_, _26324_, _09488_);
  nor (_26326_, _26325_, _03113_);
  nor (_26327_, _03311_, _03104_);
  or (_26328_, _26327_, _06188_);
  nor (_26329_, _26328_, _26326_);
  nand (_26330_, _04182_, _03161_);
  nor (_26331_, _26309_, _05444_);
  and (_26332_, _26331_, _26330_);
  nor (_26334_, _26332_, _02031_);
  not (_26335_, _26334_);
  nor (_26336_, _26335_, _26329_);
  nor (_26337_, _26291_, _02032_);
  nand (_26338_, _05075_, _04182_);
  and (_26339_, _26338_, _26337_);
  or (_26340_, _26339_, _01765_);
  nor (_26341_, _26340_, _26336_);
  nor (_26342_, _26309_, _02037_);
  nand (_26343_, _11096_, _03893_);
  and (_26345_, _26343_, _26342_);
  nor (_26346_, _26345_, _26341_);
  nor (_26347_, _26346_, _01994_);
  and (_26348_, _03893_, _04846_);
  or (_26349_, _26348_, _26291_);
  and (_26350_, _26349_, _01994_);
  or (_26351_, _26350_, _26347_);
  and (_26352_, _26351_, _03308_);
  or (_26353_, _26352_, _26299_);
  and (_26354_, _26353_, _03059_);
  nor (_26356_, _10989_, _09478_);
  or (_26357_, _26356_, _03059_);
  nor (_26358_, _26357_, _26309_);
  nor (_26359_, _26358_, _26354_);
  nor (_26360_, _26359_, _02331_);
  nor (_26361_, _26360_, _26298_);
  nor (_26362_, _26361_, _02206_);
  nor (_26363_, _10988_, _09478_);
  or (_26364_, _26363_, _02208_);
  nor (_26365_, _26364_, _26309_);
  nor (_26367_, _26365_, _26362_);
  nor (_26368_, _26367_, _09562_);
  and (_26369_, _01728_, _03104_);
  nor (_26370_, _26291_, _04209_);
  nor (_26371_, _26370_, _03065_);
  and (_26372_, _26371_, _26302_);
  or (_26373_, _26372_, _26369_);
  nor (_26374_, _26373_, _26368_);
  or (_26375_, _26374_, _17216_);
  and (_26376_, _11112_, _03893_);
  or (_26377_, _26376_, _04958_);
  nor (_26378_, _26377_, _26309_);
  and (_26379_, _04182_, _02893_);
  and (_26380_, _26379_, _04208_);
  or (_26381_, _26309_, _04953_);
  or (_26382_, _26381_, _26380_);
  nand (_26383_, _26382_, _23146_);
  nor (_26384_, _26383_, _26378_);
  and (_26385_, _26384_, _26375_);
  nor (_26386_, _26385_, _26295_);
  nor (_26388_, _26386_, _02083_);
  nor (_26389_, _02919_, _02366_);
  not (_26390_, _26389_);
  nor (_26391_, _26390_, _26388_);
  and (_26392_, _26310_, _02366_);
  nor (_26393_, _26392_, _03537_);
  not (_26394_, _26393_);
  nor (_26395_, _26394_, _26391_);
  nor (_26396_, _01990_, _03104_);
  nor (_26397_, _26396_, _02081_);
  not (_26399_, _26397_);
  nor (_26400_, _26399_, _26395_);
  nor (_26401_, _26400_, _26294_);
  nor (_26402_, _26401_, _39633_);
  nor (_26403_, _39632_, _03104_);
  or (_26404_, _26403_, rst);
  or (_41734_, _26404_, _26402_);
  and (_26405_, _05388_, _01726_);
  nor (_26406_, _04182_, _02518_);
  and (_26407_, _11315_, _04182_);
  nor (_26409_, _26407_, _26406_);
  nor (_26410_, _26409_, _03061_);
  and (_26411_, _12587_, _01718_);
  or (_26412_, _09531_, _03624_);
  nor (_26413_, _26406_, _05444_);
  and (_26414_, _26413_, _26412_);
  nor (_26415_, _12587_, _01750_);
  nor (_26416_, _11199_, _09531_);
  nor (_26417_, _26416_, _26406_);
  and (_26418_, _26417_, _02158_);
  and (_26420_, _03893_, \oc8051_golden_model_1.ACC [2]);
  nor (_26421_, _26420_, _26406_);
  or (_26422_, _26421_, _02063_);
  nand (_26423_, _09495_, \oc8051_golden_model_1.SP [2]);
  nor (_26424_, _12587_, _01747_);
  nor (_26425_, _26424_, _02158_);
  and (_26426_, _26425_, _26423_);
  and (_26427_, _26426_, _26422_);
  nor (_26428_, _26427_, _03446_);
  not (_26429_, _26428_);
  nor (_26431_, _26429_, _26418_);
  nor (_26432_, _12587_, _01745_);
  or (_26433_, _26432_, _02155_);
  nor (_26434_, _26433_, _26431_);
  and (_26435_, _04567_, _02155_);
  nor (_26436_, _26435_, _26434_);
  and (_26437_, _26436_, _02549_);
  nor (_26438_, _26421_, _02549_);
  or (_26439_, _26438_, _26437_);
  and (_26440_, _26439_, _03114_);
  or (_26442_, _26440_, _03563_);
  and (_26443_, _26442_, _01750_);
  or (_26444_, _26443_, _26415_);
  and (_26445_, _26444_, _04460_);
  and (_26446_, _05388_, _01767_);
  nor (_26447_, _26446_, _06188_);
  not (_26448_, _26447_);
  nor (_26449_, _26448_, _26445_);
  nor (_26450_, _26449_, _26414_);
  nor (_26451_, _26450_, _02031_);
  nor (_26453_, _26406_, _02032_);
  nand (_26454_, _05211_, _04182_);
  and (_26455_, _26454_, _26453_);
  or (_26456_, _26455_, _01765_);
  nor (_26457_, _26456_, _26451_);
  nor (_26458_, _11298_, _09478_);
  nor (_26459_, _26458_, _26406_);
  nor (_26460_, _26459_, _02037_);
  or (_26461_, _26460_, _01994_);
  or (_26462_, _26461_, _26457_);
  and (_26464_, _03893_, _04866_);
  nor (_26465_, _26464_, _26406_);
  nand (_26466_, _26465_, _01994_);
  and (_26467_, _26466_, _26462_);
  nor (_26468_, _26467_, _01718_);
  nor (_26469_, _26468_, _26411_);
  and (_26470_, _26469_, _03059_);
  and (_26471_, _11189_, _03893_);
  nor (_26472_, _26471_, _26406_);
  nor (_26473_, _26472_, _03059_);
  or (_26475_, _26473_, _26470_);
  and (_26476_, _26475_, _03061_);
  nor (_26477_, _26476_, _26410_);
  nor (_26478_, _26477_, _02206_);
  not (_26479_, _26406_);
  and (_26480_, _26479_, _04308_);
  or (_26481_, _26480_, _02208_);
  nor (_26482_, _26481_, _26465_);
  nor (_26483_, _26482_, _26478_);
  nor (_26484_, _26483_, _09562_);
  and (_26486_, _05388_, _01728_);
  nor (_26487_, _26486_, _02202_);
  or (_26488_, _26421_, _03065_);
  or (_26489_, _26488_, _26480_);
  nand (_26490_, _26489_, _26487_);
  nor (_26491_, _26490_, _26484_);
  nor (_26492_, _11187_, _09478_);
  nor (_26493_, _26492_, _26406_);
  and (_26494_, _26493_, _02202_);
  nor (_26495_, _26494_, _26491_);
  and (_26497_, _26495_, _04958_);
  nor (_26498_, _11314_, _09478_);
  nor (_26499_, _26498_, _26406_);
  nor (_26500_, _26499_, _04958_);
  or (_26501_, _26500_, _26497_);
  and (_26502_, _26501_, _09472_);
  and (_26503_, _12587_, _02350_);
  or (_26504_, _26503_, _26502_);
  and (_26505_, _26504_, _04964_);
  or (_26506_, _26505_, _26405_);
  and (_26508_, _26506_, _02084_);
  and (_26509_, _12587_, _02083_);
  or (_26510_, _26509_, _02366_);
  nor (_26511_, _26510_, _26508_);
  and (_26512_, _26417_, _02366_);
  nor (_26513_, _26512_, _03537_);
  not (_26514_, _26513_);
  nor (_26515_, _26514_, _26511_);
  nor (_26516_, _12587_, _01990_);
  nor (_26517_, _26516_, _02081_);
  not (_26519_, _26517_);
  nor (_26520_, _26519_, _26515_);
  and (_26521_, _11367_, _03893_);
  nor (_26522_, _26521_, _26406_);
  and (_26523_, _26522_, _02081_);
  nor (_26524_, _26523_, _26520_);
  and (_26525_, _26524_, _39632_);
  nor (_26526_, _39632_, _02518_);
  or (_26527_, _26526_, rst);
  or (_41735_, _26527_, _26525_);
  nor (_26529_, _05386_, _01990_);
  and (_26530_, _05386_, _01726_);
  nor (_26531_, _04182_, _02362_);
  and (_26532_, _11511_, _04182_);
  nor (_26533_, _26532_, _26531_);
  nor (_26534_, _26533_, _03061_);
  and (_26535_, _12348_, _01718_);
  nor (_26536_, _09478_, _03434_);
  nor (_26537_, _26536_, _26531_);
  nor (_26538_, _26537_, _05444_);
  or (_26540_, _26538_, _02031_);
  nor (_26541_, _11394_, _09531_);
  nor (_26542_, _26541_, _26531_);
  and (_26543_, _26542_, _02158_);
  and (_26544_, _03893_, \oc8051_golden_model_1.ACC [3]);
  nor (_26545_, _26544_, _26531_);
  or (_26546_, _26545_, _02063_);
  nand (_26547_, _09495_, \oc8051_golden_model_1.SP [3]);
  nor (_26548_, _12348_, _01747_);
  nor (_26549_, _26548_, _02158_);
  and (_26550_, _26549_, _26547_);
  and (_26551_, _26550_, _26546_);
  nor (_26552_, _26551_, _03446_);
  not (_26553_, _26552_);
  nor (_26554_, _26553_, _26543_);
  nor (_26555_, _12348_, _01745_);
  or (_26556_, _26555_, _02155_);
  nor (_26557_, _26556_, _26554_);
  and (_26558_, _04557_, _02155_);
  nor (_26559_, _26558_, _26557_);
  and (_26561_, _26559_, _02549_);
  nor (_26562_, _26545_, _02549_);
  or (_26563_, _26562_, _26561_);
  and (_26564_, _26563_, _03114_);
  or (_26565_, _26564_, _09488_);
  nor (_26566_, _26565_, _03485_);
  nor (_26567_, _05386_, _03311_);
  or (_26568_, _26567_, _06188_);
  nor (_26569_, _26568_, _26566_);
  nor (_26570_, _26569_, _26540_);
  nor (_26572_, _26531_, _02032_);
  nand (_26573_, _05166_, _04182_);
  and (_26574_, _26573_, _26572_);
  or (_26575_, _26574_, _01765_);
  nor (_26576_, _26575_, _26570_);
  nor (_26577_, _11490_, _09478_);
  nor (_26578_, _26577_, _26531_);
  nor (_26579_, _26578_, _02037_);
  or (_26580_, _26579_, _01994_);
  or (_26581_, _26580_, _26576_);
  and (_26583_, _03893_, _04719_);
  nor (_26584_, _26583_, _26531_);
  nand (_26585_, _26584_, _01994_);
  and (_26586_, _26585_, _26581_);
  nor (_26587_, _26586_, _01718_);
  nor (_26588_, _26587_, _26535_);
  and (_26589_, _26588_, _03059_);
  and (_26590_, _11505_, _03893_);
  nor (_26591_, _26590_, _26531_);
  nor (_26592_, _26591_, _03059_);
  or (_26594_, _26592_, _26589_);
  and (_26595_, _26594_, _03061_);
  nor (_26596_, _26595_, _26534_);
  nor (_26597_, _26596_, _02206_);
  not (_26598_, _26531_);
  and (_26599_, _26598_, _04152_);
  or (_26600_, _26599_, _02208_);
  nor (_26601_, _26600_, _26584_);
  nor (_26602_, _26601_, _26597_);
  nor (_26603_, _26602_, _09562_);
  and (_26605_, _05386_, _01728_);
  nor (_26606_, _26605_, _02202_);
  or (_26607_, _26545_, _03065_);
  or (_26608_, _26607_, _26599_);
  nand (_26609_, _26608_, _26606_);
  nor (_26610_, _26609_, _26603_);
  nor (_26611_, _11503_, _09478_);
  nor (_26612_, _26611_, _26531_);
  and (_26613_, _26612_, _02202_);
  nor (_26614_, _26613_, _26610_);
  and (_26616_, _26614_, _04958_);
  nor (_26617_, _11510_, _09478_);
  nor (_26618_, _26617_, _26531_);
  nor (_26619_, _26618_, _04958_);
  or (_26620_, _26619_, _26616_);
  and (_26621_, _26620_, _09472_);
  nor (_26622_, _04554_, _02362_);
  nor (_26623_, _26622_, _04555_);
  nor (_26624_, _26623_, _09472_);
  or (_26625_, _26624_, _26621_);
  and (_26627_, _26625_, _04964_);
  or (_26628_, _26627_, _26530_);
  and (_26629_, _26628_, _02084_);
  nor (_26630_, _26623_, _02084_);
  or (_26631_, _26630_, _26629_);
  and (_26632_, _26631_, _02778_);
  nor (_26633_, _26542_, _02778_);
  nor (_26634_, _26633_, _03537_);
  not (_26635_, _26634_);
  nor (_26636_, _26635_, _26632_);
  nor (_26638_, _26636_, _26529_);
  nor (_26639_, _26638_, _02081_);
  and (_26640_, _11567_, _03893_);
  nor (_26641_, _26640_, _26531_);
  and (_26642_, _26641_, _02081_);
  nor (_26643_, _26642_, _26639_);
  or (_26644_, _26643_, _39633_);
  or (_26645_, _39632_, \oc8051_golden_model_1.SP [3]);
  and (_26646_, _26645_, _39026_);
  and (_41736_, _26646_, _26644_);
  nor (_26648_, _03441_, \oc8051_golden_model_1.SP [4]);
  nor (_26649_, _26648_, _09465_);
  nor (_26650_, _26649_, _01990_);
  nor (_26651_, _04182_, _09510_);
  and (_26652_, _11588_, _04182_);
  nor (_26653_, _26652_, _26651_);
  nor (_26654_, _26653_, _03061_);
  nor (_26655_, _04372_, _09478_);
  nor (_26656_, _26655_, _26651_);
  nor (_26657_, _26656_, _05444_);
  or (_26659_, _26657_, _02031_);
  nor (_26660_, _11611_, _09531_);
  nor (_26661_, _26660_, _26651_);
  and (_26662_, _26661_, _02158_);
  and (_26663_, _03893_, \oc8051_golden_model_1.ACC [4]);
  nor (_26664_, _26663_, _26651_);
  or (_26665_, _26664_, _02063_);
  nand (_26666_, _09495_, \oc8051_golden_model_1.SP [4]);
  not (_26667_, _26649_);
  nor (_26668_, _26667_, _01747_);
  nor (_26669_, _26668_, _02158_);
  and (_26670_, _26669_, _26666_);
  and (_26671_, _26670_, _26665_);
  nor (_26672_, _26671_, _03446_);
  not (_26673_, _26672_);
  nor (_26674_, _26673_, _26662_);
  nor (_26675_, _26667_, _01745_);
  or (_26676_, _26675_, _02155_);
  nor (_26677_, _26676_, _26674_);
  and (_26678_, _09511_, _01986_);
  nor (_26680_, _04556_, _09510_);
  nor (_26681_, _26680_, _26678_);
  and (_26682_, _26681_, _02155_);
  nor (_26683_, _26682_, _26677_);
  and (_26684_, _26683_, _02549_);
  nor (_26685_, _26664_, _02549_);
  or (_26686_, _26685_, _26684_);
  and (_26687_, _26686_, _03114_);
  and (_26688_, _03442_, \oc8051_golden_model_1.SP [4]);
  nor (_26689_, _03442_, \oc8051_golden_model_1.SP [4]);
  nor (_26691_, _26689_, _26688_);
  and (_26692_, _26691_, _02052_);
  nor (_26693_, _26692_, _09488_);
  not (_26694_, _26693_);
  nor (_26695_, _26694_, _26687_);
  nor (_26696_, _26649_, _03311_);
  or (_26697_, _26696_, _06188_);
  nor (_26698_, _26697_, _26695_);
  nor (_26699_, _26698_, _26659_);
  nor (_26700_, _26651_, _02032_);
  nand (_26702_, _05303_, _03893_);
  and (_26703_, _26702_, _26700_);
  or (_26704_, _26703_, _01765_);
  nor (_26705_, _26704_, _26699_);
  nor (_26706_, _11704_, _09478_);
  nor (_26707_, _26706_, _26651_);
  nor (_26708_, _26707_, _02037_);
  or (_26709_, _26708_, _01994_);
  or (_26710_, _26709_, _26705_);
  and (_26711_, _04831_, _03893_);
  nor (_26713_, _26711_, _26651_);
  nand (_26714_, _26713_, _01994_);
  and (_26715_, _26714_, _26710_);
  nor (_26716_, _26715_, _01718_);
  and (_26717_, _26667_, _01718_);
  nor (_26718_, _26717_, _26716_);
  and (_26719_, _26718_, _03059_);
  and (_26720_, _11592_, _03893_);
  nor (_26721_, _26720_, _26651_);
  nor (_26722_, _26721_, _03059_);
  or (_26724_, _26722_, _26719_);
  and (_26725_, _26724_, _03061_);
  nor (_26726_, _26725_, _26654_);
  nor (_26727_, _26726_, _02206_);
  nor (_26728_, _26651_, _04420_);
  not (_26729_, _26728_);
  nor (_26730_, _26713_, _02208_);
  and (_26731_, _26730_, _26729_);
  nor (_26732_, _26731_, _26727_);
  nor (_26733_, _26732_, _09562_);
  and (_26735_, _26649_, _01728_);
  or (_26736_, _26728_, _03065_);
  nor (_26737_, _26736_, _26664_);
  or (_26738_, _26737_, _26735_);
  or (_26739_, _26738_, _02202_);
  nor (_26740_, _26739_, _26733_);
  nor (_26741_, _11590_, _09478_);
  nor (_26742_, _26741_, _26651_);
  and (_26743_, _26742_, _02202_);
  nor (_26744_, _26743_, _26740_);
  and (_26746_, _26744_, _04958_);
  nor (_26747_, _11587_, _09478_);
  nor (_26748_, _26747_, _26651_);
  nor (_26749_, _26748_, _04958_);
  or (_26750_, _26749_, _26746_);
  and (_26751_, _26750_, _09472_);
  nor (_26752_, _04555_, _09510_);
  nor (_26753_, _26752_, _09511_);
  nor (_26754_, _26753_, _09472_);
  or (_26755_, _26754_, _01726_);
  nor (_26757_, _26755_, _26751_);
  and (_26758_, _26667_, _01726_);
  nor (_26759_, _26758_, _26757_);
  and (_26760_, _26759_, _02084_);
  nor (_26761_, _26753_, _02084_);
  or (_26762_, _26761_, _26760_);
  and (_26763_, _26762_, _02778_);
  nor (_26764_, _26661_, _02778_);
  nor (_26765_, _26764_, _03537_);
  not (_26766_, _26765_);
  nor (_26768_, _26766_, _26763_);
  nor (_26769_, _26768_, _26650_);
  nor (_26770_, _26769_, _02081_);
  and (_26771_, _11771_, _03893_);
  nor (_26772_, _26771_, _26651_);
  and (_26773_, _26772_, _02081_);
  nor (_26774_, _26773_, _26770_);
  or (_26775_, _26774_, _39633_);
  or (_26776_, _39632_, \oc8051_golden_model_1.SP [4]);
  and (_26777_, _26776_, _39026_);
  and (_41738_, _26777_, _26775_);
  nor (_26779_, _09465_, \oc8051_golden_model_1.SP [5]);
  nor (_26780_, _26779_, _09466_);
  nor (_26781_, _26780_, _01990_);
  nor (_26782_, _04182_, _09509_);
  and (_26783_, _11786_, _04182_);
  nor (_26784_, _26783_, _26782_);
  nor (_26785_, _26784_, _03061_);
  nor (_26786_, _04057_, _09478_);
  nor (_26787_, _26786_, _26782_);
  nor (_26789_, _26787_, _05444_);
  or (_26790_, _26789_, _02031_);
  nor (_26791_, _11804_, _09531_);
  nor (_26792_, _26791_, _26782_);
  and (_26793_, _26792_, _02158_);
  and (_26794_, _03893_, \oc8051_golden_model_1.ACC [5]);
  nor (_26795_, _26794_, _26782_);
  or (_26796_, _26795_, _02063_);
  nand (_26797_, _09495_, \oc8051_golden_model_1.SP [5]);
  not (_26798_, _26780_);
  nor (_26799_, _26798_, _01747_);
  nor (_26800_, _26799_, _02158_);
  and (_26801_, _26800_, _26797_);
  and (_26802_, _26801_, _26796_);
  nor (_26803_, _26802_, _03446_);
  not (_26804_, _26803_);
  nor (_26805_, _26804_, _26793_);
  nor (_26806_, _26798_, _01745_);
  or (_26807_, _26806_, _02155_);
  nor (_26808_, _26807_, _26805_);
  and (_26810_, _09512_, _01986_);
  nor (_26811_, _26678_, _09509_);
  nor (_26812_, _26811_, _26810_);
  and (_26813_, _26812_, _02155_);
  nor (_26814_, _26813_, _26808_);
  and (_26815_, _26814_, _02549_);
  nor (_26816_, _26795_, _02549_);
  or (_26817_, _26816_, _26815_);
  and (_26818_, _26817_, _03114_);
  and (_26819_, _09466_, \oc8051_golden_model_1.SP [0]);
  nor (_26821_, _26688_, \oc8051_golden_model_1.SP [5]);
  nor (_26822_, _26821_, _26819_);
  and (_26823_, _26822_, _02052_);
  nor (_26824_, _26823_, _09488_);
  not (_26825_, _26824_);
  nor (_26826_, _26825_, _26818_);
  nor (_26827_, _26780_, _03311_);
  or (_26828_, _26827_, _06188_);
  nor (_26829_, _26828_, _26826_);
  nor (_26830_, _26829_, _26790_);
  nor (_26832_, _26782_, _02032_);
  nand (_26833_, _05258_, _04182_);
  and (_26834_, _26833_, _26832_);
  or (_26835_, _26834_, _01765_);
  nor (_26836_, _26835_, _26830_);
  nor (_26837_, _11900_, _09478_);
  nor (_26838_, _26837_, _26782_);
  nor (_26839_, _26838_, _02037_);
  or (_26840_, _26839_, _01994_);
  or (_26841_, _26840_, _26836_);
  and (_26843_, _04827_, _03893_);
  nor (_26844_, _26843_, _26782_);
  nand (_26845_, _26844_, _01994_);
  and (_26846_, _26845_, _26841_);
  nor (_26847_, _26846_, _01718_);
  and (_26848_, _26798_, _01718_);
  nor (_26849_, _26848_, _26847_);
  and (_26850_, _26849_, _03059_);
  and (_26851_, _11915_, _03893_);
  nor (_26852_, _26851_, _26782_);
  nor (_26854_, _26852_, _03059_);
  or (_26855_, _26854_, _26850_);
  and (_26856_, _26855_, _03061_);
  nor (_26857_, _26856_, _26785_);
  nor (_26858_, _26857_, _02206_);
  nor (_26859_, _26782_, _04104_);
  not (_26860_, _26859_);
  nor (_26861_, _26844_, _02208_);
  and (_26862_, _26861_, _26860_);
  nor (_26863_, _26862_, _26858_);
  nor (_26865_, _26863_, _09562_);
  and (_26866_, _26780_, _01728_);
  or (_26867_, _26859_, _03065_);
  nor (_26868_, _26867_, _26795_);
  or (_26869_, _26868_, _26866_);
  or (_26870_, _26869_, _02202_);
  nor (_26871_, _26870_, _26865_);
  nor (_26872_, _11913_, _09478_);
  nor (_26873_, _26872_, _26782_);
  and (_26874_, _26873_, _02202_);
  nor (_26876_, _26874_, _26871_);
  and (_26877_, _26876_, _04958_);
  nor (_26878_, _11785_, _09478_);
  nor (_26879_, _26878_, _26782_);
  nor (_26880_, _26879_, _04958_);
  or (_26881_, _26880_, _26877_);
  and (_26882_, _26881_, _09472_);
  nor (_26883_, _09511_, _09509_);
  nor (_26884_, _26883_, _09512_);
  nor (_26885_, _26884_, _09472_);
  or (_26887_, _26885_, _01726_);
  nor (_26888_, _26887_, _26882_);
  and (_26889_, _26798_, _01726_);
  nor (_26890_, _26889_, _26888_);
  and (_26891_, _26890_, _02084_);
  nor (_26892_, _26884_, _02084_);
  or (_26893_, _26892_, _26891_);
  and (_26894_, _26893_, _02778_);
  nor (_26895_, _26792_, _02778_);
  nor (_26896_, _26895_, _03537_);
  not (_26898_, _26896_);
  nor (_26899_, _26898_, _26894_);
  nor (_26900_, _26899_, _26781_);
  nor (_26901_, _26900_, _02081_);
  and (_26902_, _11974_, _03893_);
  nor (_26903_, _26902_, _26782_);
  and (_26904_, _26903_, _02081_);
  nor (_26905_, _26904_, _26901_);
  or (_26906_, _26905_, _39633_);
  or (_26907_, _39632_, \oc8051_golden_model_1.SP [5]);
  and (_26909_, _26907_, _39026_);
  and (_41739_, _26909_, _26906_);
  nor (_26910_, _04182_, _09508_);
  and (_26911_, _12118_, _04182_);
  nor (_26912_, _26911_, _26910_);
  nor (_26913_, _26912_, _03061_);
  or (_26914_, _03964_, _09531_);
  nor (_26915_, _26910_, _05444_);
  and (_26916_, _26915_, _26914_);
  nor (_26917_, _11993_, _09531_);
  nor (_26919_, _26917_, _26910_);
  and (_26920_, _26919_, _02158_);
  and (_26921_, _03893_, \oc8051_golden_model_1.ACC [6]);
  nor (_26922_, _26921_, _26910_);
  or (_26923_, _26922_, _02063_);
  nand (_26924_, _09495_, \oc8051_golden_model_1.SP [6]);
  nor (_26925_, _09466_, \oc8051_golden_model_1.SP [6]);
  nor (_26926_, _26925_, _09467_);
  not (_26927_, _26926_);
  nor (_26928_, _26927_, _01747_);
  nor (_26930_, _26928_, _02158_);
  and (_26931_, _26930_, _26924_);
  and (_26932_, _26931_, _26923_);
  nor (_26933_, _26932_, _03446_);
  not (_26934_, _26933_);
  nor (_26935_, _26934_, _26920_);
  nor (_26936_, _26927_, _01745_);
  or (_26937_, _26936_, _02155_);
  nor (_26938_, _26937_, _26935_);
  nor (_26939_, _26810_, _09508_);
  nor (_26940_, _26939_, _09514_);
  and (_26941_, _26940_, _02155_);
  nor (_26942_, _26941_, _26938_);
  and (_26943_, _26942_, _02549_);
  nor (_26944_, _26922_, _02549_);
  or (_26945_, _26944_, _26943_);
  and (_26946_, _26945_, _03114_);
  nor (_26947_, _26819_, \oc8051_golden_model_1.SP [6]);
  nor (_26948_, _26947_, _09483_);
  and (_26949_, _26948_, _02052_);
  nor (_26951_, _26949_, _26946_);
  nor (_26952_, _26951_, _09488_);
  nor (_26953_, _26927_, _03311_);
  nor (_26954_, _26953_, _06188_);
  not (_26955_, _26954_);
  nor (_26956_, _26955_, _26952_);
  nor (_26957_, _26956_, _26916_);
  nor (_26958_, _26957_, _02031_);
  nor (_26959_, _26910_, _02032_);
  nand (_26960_, _05029_, _04182_);
  and (_26962_, _26960_, _26959_);
  or (_26963_, _26962_, _01765_);
  nor (_26964_, _26963_, _26958_);
  nor (_26965_, _12096_, _09478_);
  nor (_26966_, _26965_, _26910_);
  nor (_26967_, _26966_, _02037_);
  or (_26968_, _26967_, _01994_);
  or (_26969_, _26968_, _26964_);
  and (_26970_, _12103_, _03893_);
  nor (_26971_, _26970_, _26910_);
  nand (_26973_, _26971_, _01994_);
  and (_26974_, _26973_, _26969_);
  nor (_26975_, _26974_, _01718_);
  and (_26976_, _26927_, _01718_);
  nor (_26977_, _26976_, _26975_);
  and (_26978_, _26977_, _03059_);
  and (_26979_, _12112_, _03893_);
  nor (_26980_, _26979_, _26910_);
  nor (_26981_, _26980_, _03059_);
  or (_26982_, _26981_, _26978_);
  and (_26984_, _26982_, _03061_);
  nor (_26985_, _26984_, _26913_);
  nor (_26986_, _26985_, _02206_);
  nor (_26987_, _26910_, _04011_);
  not (_26988_, _26987_);
  nor (_26989_, _26971_, _02208_);
  and (_26990_, _26989_, _26988_);
  nor (_26991_, _26990_, _26986_);
  nor (_26992_, _26991_, _09562_);
  and (_26993_, _26926_, _01728_);
  or (_26995_, _26987_, _03065_);
  nor (_26996_, _26995_, _26922_);
  or (_26997_, _26996_, _26993_);
  or (_26998_, _26997_, _02202_);
  nor (_26999_, _26998_, _26992_);
  nor (_27000_, _12110_, _09478_);
  nor (_27001_, _27000_, _26910_);
  and (_27002_, _27001_, _02202_);
  nor (_27003_, _27002_, _26999_);
  and (_27004_, _27003_, _04958_);
  nor (_27006_, _12117_, _09478_);
  nor (_27007_, _27006_, _26910_);
  nor (_27008_, _27007_, _04958_);
  or (_27009_, _27008_, _27004_);
  and (_27010_, _27009_, _09472_);
  nor (_27011_, _09512_, _09508_);
  nor (_27012_, _27011_, _09513_);
  not (_27013_, _27012_);
  nor (_27014_, _27013_, _01726_);
  nor (_27015_, _27014_, _23146_);
  nor (_27017_, _27015_, _27010_);
  and (_27018_, _26927_, _01726_);
  or (_27019_, _27018_, _02083_);
  nor (_27020_, _27019_, _27017_);
  and (_27021_, _27013_, _02083_);
  or (_27022_, _27021_, _02366_);
  nor (_27023_, _27022_, _27020_);
  and (_27024_, _26919_, _02366_);
  nor (_27025_, _27024_, _03537_);
  not (_27026_, _27025_);
  nor (_27028_, _27026_, _27023_);
  nor (_27029_, _26927_, _01990_);
  nor (_27030_, _27029_, _02081_);
  not (_27031_, _27030_);
  nor (_27032_, _27031_, _27028_);
  and (_27033_, _12178_, _03893_);
  nor (_27034_, _27033_, _26910_);
  and (_27035_, _27034_, _02081_);
  nor (_27036_, _27035_, _27032_);
  or (_27037_, _27036_, _39633_);
  or (_27039_, _39632_, \oc8051_golden_model_1.SP [6]);
  and (_27040_, _27039_, _39026_);
  and (_41740_, _27040_, _27037_);
  nor (_27041_, _04257_, _09607_);
  not (_27042_, \oc8051_golden_model_1.TCON [0]);
  nor (_27043_, _03856_, _27042_);
  and (_27044_, _03856_, _04837_);
  nor (_27045_, _27044_, _27043_);
  nor (_27046_, _27045_, _02208_);
  not (_27047_, _27046_);
  nor (_27049_, _27047_, _27041_);
  and (_27050_, _10792_, _03856_);
  nor (_27051_, _27050_, _27043_);
  nor (_27052_, _27051_, _03061_);
  and (_27053_, _27045_, _01994_);
  and (_27054_, _03856_, _03002_);
  nor (_27055_, _27054_, _27043_);
  and (_27056_, _27055_, _06188_);
  and (_27057_, _03856_, \oc8051_golden_model_1.ACC [0]);
  nor (_27058_, _27057_, _27043_);
  nor (_27060_, _27058_, _02063_);
  nor (_27061_, _02062_, _27042_);
  or (_27062_, _27061_, _27060_);
  and (_27063_, _27062_, _03006_);
  nor (_27064_, _27043_, _27041_);
  nor (_27065_, _27064_, _03006_);
  or (_27066_, _27065_, _27063_);
  and (_27067_, _27066_, _02058_);
  nor (_27068_, _04487_, _27042_);
  and (_27069_, _10814_, _04487_);
  nor (_27071_, _27069_, _27068_);
  nor (_27072_, _27071_, _02058_);
  nor (_27073_, _27072_, _27067_);
  nor (_27074_, _27073_, _02155_);
  nor (_27075_, _27055_, _02519_);
  or (_27076_, _27075_, _27074_);
  and (_27077_, _27076_, _02549_);
  nor (_27078_, _27058_, _02549_);
  or (_27079_, _27078_, _27077_);
  and (_27080_, _27079_, _02054_);
  and (_27081_, _27043_, _02053_);
  or (_27082_, _27081_, _27080_);
  and (_27083_, _27082_, _02047_);
  nor (_27084_, _27064_, _02047_);
  or (_27085_, _27084_, _27083_);
  and (_27086_, _27085_, _02043_);
  nor (_27087_, _10798_, _09644_);
  nor (_27088_, _27087_, _27068_);
  nor (_27089_, _27088_, _02043_);
  or (_27090_, _27089_, _06188_);
  nor (_27092_, _27090_, _27086_);
  nor (_27093_, _27092_, _27056_);
  nor (_27094_, _27093_, _02031_);
  and (_27095_, _05120_, _03856_);
  nor (_27096_, _27043_, _02032_);
  not (_27097_, _27096_);
  nor (_27098_, _27097_, _27095_);
  or (_27099_, _27098_, _01765_);
  nor (_27100_, _27099_, _27094_);
  nor (_27101_, _10898_, _09607_);
  nor (_27103_, _27101_, _27043_);
  nor (_27104_, _27103_, _02037_);
  or (_27105_, _27104_, _01994_);
  nor (_27106_, _27105_, _27100_);
  nor (_27107_, _27106_, _27053_);
  or (_27108_, _27107_, _02210_);
  and (_27109_, _10914_, _03856_);
  or (_27110_, _27109_, _27043_);
  or (_27111_, _27110_, _03059_);
  and (_27112_, _27111_, _03061_);
  and (_27114_, _27112_, _27108_);
  nor (_27115_, _27114_, _27052_);
  nor (_27116_, _27115_, _02206_);
  nor (_27117_, _27116_, _27049_);
  nor (_27118_, _27117_, _02342_);
  nor (_27119_, _27043_, _04257_);
  or (_27120_, _27119_, _03065_);
  nor (_27121_, _27120_, _27058_);
  or (_27122_, _27121_, _02202_);
  nor (_27123_, _27122_, _27118_);
  nor (_27125_, _10913_, _09607_);
  or (_27126_, _27043_, _04953_);
  nor (_27127_, _27126_, _27125_);
  or (_27128_, _27127_, _02334_);
  nor (_27129_, _27128_, _27123_);
  nor (_27130_, _10789_, _09607_);
  nor (_27131_, _27130_, _27043_);
  nor (_27132_, _27131_, _04958_);
  or (_27133_, _27132_, _27129_);
  and (_27134_, _27133_, _02778_);
  nor (_27136_, _27064_, _02778_);
  or (_27137_, _27136_, _27134_);
  and (_27138_, _27137_, _01698_);
  and (_27139_, _27043_, _01697_);
  nor (_27140_, _27139_, _02081_);
  not (_27141_, _27140_);
  nor (_27142_, _27141_, _27138_);
  and (_27143_, _27064_, _02081_);
  or (_27144_, _27143_, _27142_);
  nand (_27145_, _27144_, _39632_);
  or (_27147_, _39632_, \oc8051_golden_model_1.TCON [0]);
  and (_27148_, _27147_, _39026_);
  and (_41742_, _27148_, _27145_);
  not (_27149_, \oc8051_golden_model_1.TCON [1]);
  nor (_27150_, _03856_, _27149_);
  nor (_27151_, _09607_, _03161_);
  or (_27152_, _27151_, _27150_);
  or (_27153_, _27152_, _02519_);
  or (_27154_, _03856_, \oc8051_golden_model_1.TCON [1]);
  and (_27155_, _11001_, _03856_);
  not (_27157_, _27155_);
  and (_27158_, _27157_, _27154_);
  or (_27159_, _27158_, _03006_);
  nand (_27160_, _03856_, _01804_);
  and (_27161_, _27160_, _27154_);
  and (_27162_, _27161_, _02062_);
  nor (_27163_, _02062_, _27149_);
  or (_27164_, _27163_, _02158_);
  or (_27165_, _27164_, _27162_);
  and (_27166_, _27165_, _02058_);
  and (_27168_, _27166_, _27159_);
  nor (_27169_, _04487_, _27149_);
  and (_27170_, _11005_, _04487_);
  or (_27171_, _27170_, _27169_);
  and (_27172_, _27171_, _02057_);
  or (_27173_, _27172_, _02155_);
  or (_27174_, _27173_, _27168_);
  and (_27175_, _27174_, _27153_);
  or (_27176_, _27175_, _02153_);
  or (_27177_, _27161_, _02549_);
  and (_27179_, _27177_, _02054_);
  and (_27180_, _27179_, _27176_);
  and (_27181_, _10992_, _04487_);
  or (_27182_, _27181_, _27169_);
  and (_27183_, _27182_, _02053_);
  or (_27184_, _27183_, _27180_);
  or (_27185_, _27184_, _02046_);
  or (_27186_, _27169_, _11020_);
  and (_27187_, _27186_, _27171_);
  or (_27188_, _27187_, _02047_);
  and (_27190_, _27188_, _02043_);
  and (_27191_, _27190_, _27185_);
  nor (_27192_, _11038_, _09644_);
  or (_27193_, _27192_, _27169_);
  and (_27194_, _27193_, _02042_);
  or (_27195_, _27194_, _06188_);
  or (_27196_, _27195_, _27191_);
  or (_27197_, _27152_, _05444_);
  and (_27198_, _27197_, _27196_);
  or (_27199_, _27198_, _02031_);
  and (_27201_, _05075_, _03856_);
  or (_27202_, _27150_, _02032_);
  or (_27203_, _27202_, _27201_);
  and (_27204_, _27203_, _02037_);
  and (_27205_, _27204_, _27199_);
  nor (_27206_, _11096_, _09607_);
  or (_27207_, _27206_, _27150_);
  and (_27208_, _27207_, _01765_);
  or (_27209_, _27208_, _27205_);
  and (_27210_, _27209_, _02212_);
  or (_27212_, _10989_, _09607_);
  and (_27213_, _27212_, _02210_);
  nand (_27214_, _03856_, _02893_);
  and (_27215_, _27214_, _01994_);
  or (_27216_, _27215_, _27213_);
  and (_27217_, _27216_, _27154_);
  or (_27218_, _27217_, _27210_);
  and (_27219_, _27218_, _03061_);
  or (_27220_, _11113_, _09607_);
  and (_27221_, _27154_, _02331_);
  and (_27223_, _27221_, _27220_);
  or (_27224_, _27223_, _27219_);
  and (_27225_, _27224_, _02208_);
  or (_27226_, _10988_, _09607_);
  and (_27227_, _27154_, _02206_);
  and (_27228_, _27227_, _27226_);
  or (_27229_, _27228_, _27225_);
  and (_27230_, _27229_, _03065_);
  or (_27231_, _27150_, _04209_);
  and (_27232_, _27161_, _02342_);
  and (_27233_, _27232_, _27231_);
  or (_27234_, _27233_, _27230_);
  and (_27235_, _27234_, _02335_);
  or (_27236_, _27160_, _04209_);
  and (_27237_, _27154_, _02334_);
  and (_27238_, _27237_, _27236_);
  or (_27239_, _27238_, _02366_);
  or (_27240_, _27214_, _04209_);
  and (_27241_, _27154_, _02202_);
  and (_27242_, _27241_, _27240_);
  or (_27244_, _27242_, _27239_);
  or (_27245_, _27244_, _27235_);
  or (_27246_, _27158_, _02778_);
  and (_27247_, _27246_, _01698_);
  and (_27248_, _27247_, _27245_);
  and (_27249_, _27182_, _01697_);
  or (_27250_, _27249_, _02081_);
  or (_27251_, _27250_, _27248_);
  or (_27252_, _27155_, _27150_);
  or (_27253_, _27252_, _02082_);
  and (_27255_, _27253_, _27251_);
  and (_27256_, _27255_, _39632_);
  nor (_27257_, _39632_, _27149_);
  or (_27258_, _27257_, rst);
  or (_41743_, _27258_, _27256_);
  not (_27259_, \oc8051_golden_model_1.TCON [2]);
  nor (_27260_, _03856_, _27259_);
  and (_27261_, _03856_, _04866_);
  nor (_27262_, _27261_, _27260_);
  and (_27263_, _27262_, _01994_);
  nor (_27265_, _09607_, _03624_);
  nor (_27266_, _27265_, _27260_);
  and (_27267_, _27266_, _06188_);
  and (_27268_, _03856_, \oc8051_golden_model_1.ACC [2]);
  nor (_27269_, _27268_, _27260_);
  nor (_27270_, _27269_, _02063_);
  nor (_27271_, _02062_, _27259_);
  or (_27272_, _27271_, _27270_);
  and (_27273_, _27272_, _03006_);
  nor (_27274_, _11199_, _09607_);
  nor (_27276_, _27274_, _27260_);
  nor (_27277_, _27276_, _03006_);
  or (_27278_, _27277_, _27273_);
  and (_27279_, _27278_, _02058_);
  nor (_27280_, _04487_, _27259_);
  and (_27281_, _11194_, _04487_);
  nor (_27282_, _27281_, _27280_);
  nor (_27283_, _27282_, _02058_);
  or (_27284_, _27283_, _02155_);
  or (_27285_, _27284_, _27279_);
  nand (_27287_, _27266_, _02155_);
  and (_27288_, _27287_, _27285_);
  and (_27289_, _27288_, _02549_);
  nor (_27290_, _27269_, _02549_);
  or (_27291_, _27290_, _27289_);
  and (_27292_, _27291_, _02054_);
  and (_27293_, _11192_, _04487_);
  nor (_27294_, _27293_, _27280_);
  nor (_27295_, _27294_, _02054_);
  or (_27296_, _27295_, _27292_);
  and (_27298_, _27296_, _02047_);
  nor (_27299_, _27280_, _11223_);
  nor (_27300_, _27299_, _27282_);
  and (_27301_, _27300_, _02046_);
  or (_27302_, _27301_, _27298_);
  and (_27303_, _27302_, _02043_);
  nor (_27304_, _11241_, _09644_);
  nor (_27305_, _27304_, _27280_);
  nor (_27306_, _27305_, _02043_);
  nor (_27307_, _27306_, _06188_);
  not (_27309_, _27307_);
  nor (_27310_, _27309_, _27303_);
  nor (_27311_, _27310_, _27267_);
  nor (_27312_, _27311_, _02031_);
  and (_27313_, _05211_, _03856_);
  nor (_27314_, _27260_, _02032_);
  not (_27315_, _27314_);
  nor (_27316_, _27315_, _27313_);
  or (_27317_, _27316_, _01765_);
  nor (_27318_, _27317_, _27312_);
  nor (_27320_, _11298_, _09607_);
  nor (_27321_, _27260_, _27320_);
  nor (_27322_, _27321_, _02037_);
  or (_27323_, _27322_, _01994_);
  nor (_27324_, _27323_, _27318_);
  nor (_27325_, _27324_, _27263_);
  or (_27326_, _27325_, _02210_);
  and (_27327_, _11189_, _03856_);
  or (_27328_, _27327_, _27260_);
  or (_27329_, _27328_, _03059_);
  and (_27331_, _27329_, _03061_);
  and (_27332_, _27331_, _27326_);
  and (_27333_, _11315_, _03856_);
  nor (_27334_, _27333_, _27260_);
  nor (_27335_, _27334_, _03061_);
  nor (_27336_, _27335_, _27332_);
  nor (_27337_, _27336_, _02206_);
  nor (_27338_, _27260_, _04309_);
  not (_27339_, _27338_);
  nor (_27340_, _27262_, _02208_);
  and (_27342_, _27340_, _27339_);
  nor (_27343_, _27342_, _27337_);
  nor (_27344_, _27343_, _02342_);
  or (_27345_, _27338_, _03065_);
  nor (_27346_, _27345_, _27269_);
  or (_27347_, _27346_, _02202_);
  nor (_27348_, _27347_, _27344_);
  nor (_27349_, _11187_, _09607_);
  or (_27350_, _27260_, _04953_);
  nor (_27351_, _27350_, _27349_);
  or (_27353_, _27351_, _02334_);
  nor (_27354_, _27353_, _27348_);
  nor (_27355_, _11314_, _09607_);
  nor (_27356_, _27355_, _27260_);
  nor (_27357_, _27356_, _04958_);
  or (_27358_, _27357_, _27354_);
  and (_27359_, _27358_, _02778_);
  nor (_27360_, _27276_, _02778_);
  or (_27361_, _27360_, _27359_);
  and (_27362_, _27361_, _01698_);
  nor (_27364_, _27294_, _01698_);
  or (_27365_, _27364_, _27362_);
  and (_27366_, _27365_, _02082_);
  and (_27367_, _11367_, _03856_);
  nor (_27368_, _27367_, _27260_);
  nor (_27369_, _27368_, _02082_);
  or (_27370_, _27369_, _27366_);
  or (_27371_, _27370_, _39633_);
  or (_27372_, _39632_, \oc8051_golden_model_1.TCON [2]);
  and (_27373_, _27372_, _39026_);
  and (_41744_, _27373_, _27371_);
  not (_27374_, \oc8051_golden_model_1.TCON [3]);
  nor (_27375_, _03856_, _27374_);
  and (_27376_, _03856_, _04719_);
  nor (_27377_, _27376_, _27375_);
  and (_27378_, _27377_, _01994_);
  nor (_27379_, _09607_, _03434_);
  nor (_27380_, _27379_, _27375_);
  and (_27381_, _27380_, _06188_);
  and (_27382_, _03856_, \oc8051_golden_model_1.ACC [3]);
  nor (_27384_, _27382_, _27375_);
  nor (_27385_, _27384_, _02063_);
  nor (_27386_, _02062_, _27374_);
  or (_27387_, _27386_, _27385_);
  and (_27388_, _27387_, _03006_);
  nor (_27389_, _11394_, _09607_);
  nor (_27390_, _27389_, _27375_);
  nor (_27391_, _27390_, _03006_);
  or (_27392_, _27391_, _27388_);
  and (_27393_, _27392_, _02058_);
  nor (_27395_, _04487_, _27374_);
  and (_27396_, _11398_, _04487_);
  nor (_27397_, _27396_, _27395_);
  nor (_27398_, _27397_, _02058_);
  or (_27399_, _27398_, _27393_);
  and (_27400_, _27399_, _02519_);
  nor (_27401_, _27380_, _02519_);
  or (_27402_, _27401_, _27400_);
  and (_27403_, _27402_, _02549_);
  nor (_27404_, _27384_, _02549_);
  or (_27406_, _27404_, _27403_);
  and (_27407_, _27406_, _02054_);
  and (_27408_, _11408_, _04487_);
  nor (_27409_, _27408_, _27395_);
  nor (_27410_, _27409_, _02054_);
  or (_27411_, _27410_, _27407_);
  and (_27412_, _27411_, _02047_);
  nor (_27413_, _27395_, _11415_);
  nor (_27414_, _27413_, _27397_);
  and (_27415_, _27414_, _02046_);
  or (_27417_, _27415_, _27412_);
  and (_27418_, _27417_, _02043_);
  nor (_27419_, _11433_, _09644_);
  nor (_27420_, _27419_, _27395_);
  nor (_27421_, _27420_, _02043_);
  nor (_27422_, _27421_, _06188_);
  not (_27423_, _27422_);
  nor (_27424_, _27423_, _27418_);
  nor (_27425_, _27424_, _27381_);
  nor (_27426_, _27425_, _02031_);
  and (_27428_, _05166_, _03856_);
  nor (_27429_, _27375_, _02032_);
  not (_27430_, _27429_);
  nor (_27431_, _27430_, _27428_);
  or (_27432_, _27431_, _01765_);
  nor (_27433_, _27432_, _27426_);
  nor (_27434_, _11490_, _09607_);
  nor (_27435_, _27375_, _27434_);
  nor (_27436_, _27435_, _02037_);
  or (_27437_, _27436_, _01994_);
  nor (_27439_, _27437_, _27433_);
  nor (_27440_, _27439_, _27378_);
  or (_27441_, _27440_, _02210_);
  and (_27442_, _11505_, _03856_);
  or (_27443_, _27442_, _27375_);
  or (_27444_, _27443_, _03059_);
  and (_27445_, _27444_, _03061_);
  and (_27446_, _27445_, _27441_);
  and (_27447_, _11511_, _03856_);
  nor (_27448_, _27447_, _27375_);
  nor (_27450_, _27448_, _03061_);
  nor (_27451_, _27450_, _27446_);
  nor (_27452_, _27451_, _02206_);
  nor (_27453_, _27375_, _04153_);
  not (_27454_, _27453_);
  nor (_27455_, _27377_, _02208_);
  and (_27456_, _27455_, _27454_);
  nor (_27457_, _27456_, _27452_);
  nor (_27458_, _27457_, _02342_);
  or (_27459_, _27453_, _03065_);
  nor (_27461_, _27459_, _27384_);
  or (_27462_, _27461_, _02202_);
  nor (_27463_, _27462_, _27458_);
  nor (_27464_, _11503_, _09607_);
  or (_27465_, _27375_, _04953_);
  nor (_27466_, _27465_, _27464_);
  or (_27467_, _27466_, _02334_);
  nor (_27468_, _27467_, _27463_);
  nor (_27469_, _11510_, _09607_);
  nor (_27470_, _27469_, _27375_);
  nor (_27472_, _27470_, _04958_);
  or (_27473_, _27472_, _27468_);
  and (_27474_, _27473_, _02778_);
  nor (_27475_, _27390_, _02778_);
  or (_27476_, _27475_, _27474_);
  and (_27477_, _27476_, _01698_);
  nor (_27478_, _27409_, _01698_);
  or (_27479_, _27478_, _27477_);
  and (_27480_, _27479_, _02082_);
  and (_27481_, _11567_, _03856_);
  nor (_27483_, _27481_, _27375_);
  nor (_27484_, _27483_, _02082_);
  or (_27485_, _27484_, _27480_);
  or (_27486_, _27485_, _39633_);
  or (_27487_, _39632_, \oc8051_golden_model_1.TCON [3]);
  and (_27488_, _27487_, _39026_);
  and (_41745_, _27488_, _27486_);
  not (_27489_, \oc8051_golden_model_1.TCON [4]);
  nor (_27490_, _03856_, _27489_);
  and (_27491_, _04831_, _03856_);
  nor (_27493_, _27491_, _27490_);
  and (_27494_, _27493_, _01994_);
  nor (_27495_, _04372_, _09607_);
  nor (_27496_, _27495_, _27490_);
  and (_27497_, _27496_, _06188_);
  and (_27498_, _03856_, \oc8051_golden_model_1.ACC [4]);
  nor (_27499_, _27498_, _27490_);
  nor (_27500_, _27499_, _02063_);
  nor (_27501_, _02062_, _27489_);
  or (_27502_, _27501_, _27500_);
  and (_27504_, _27502_, _03006_);
  nor (_27505_, _11611_, _09607_);
  nor (_27506_, _27505_, _27490_);
  nor (_27507_, _27506_, _03006_);
  or (_27508_, _27507_, _27504_);
  and (_27509_, _27508_, _02058_);
  nor (_27510_, _04487_, _27489_);
  and (_27511_, _11597_, _04487_);
  nor (_27512_, _27511_, _27510_);
  nor (_27513_, _27512_, _02058_);
  or (_27515_, _27513_, _27509_);
  and (_27516_, _27515_, _02519_);
  nor (_27517_, _27496_, _02519_);
  or (_27518_, _27517_, _27516_);
  and (_27519_, _27518_, _02549_);
  nor (_27520_, _27499_, _02549_);
  or (_27521_, _27520_, _27519_);
  and (_27522_, _27521_, _02054_);
  and (_27523_, _11595_, _04487_);
  nor (_27524_, _27523_, _27510_);
  nor (_27526_, _27524_, _02054_);
  or (_27527_, _27526_, _27522_);
  and (_27528_, _27527_, _02047_);
  nor (_27529_, _27510_, _11628_);
  nor (_27530_, _27529_, _27512_);
  and (_27531_, _27530_, _02046_);
  or (_27532_, _27531_, _27528_);
  and (_27533_, _27532_, _02043_);
  nor (_27534_, _11646_, _09644_);
  nor (_27535_, _27534_, _27510_);
  nor (_27537_, _27535_, _02043_);
  nor (_27538_, _27537_, _06188_);
  not (_27539_, _27538_);
  nor (_27540_, _27539_, _27533_);
  nor (_27541_, _27540_, _27497_);
  nor (_27542_, _27541_, _02031_);
  and (_27543_, _05303_, _03856_);
  nor (_27544_, _27490_, _02032_);
  not (_27545_, _27544_);
  nor (_27546_, _27545_, _27543_);
  or (_27547_, _27546_, _01765_);
  nor (_27548_, _27547_, _27542_);
  nor (_27549_, _11704_, _09607_);
  nor (_27550_, _27490_, _27549_);
  nor (_27551_, _27550_, _02037_);
  or (_27552_, _27551_, _01994_);
  nor (_27553_, _27552_, _27548_);
  nor (_27554_, _27553_, _27494_);
  or (_27555_, _27554_, _02210_);
  and (_27556_, _11592_, _03856_);
  or (_27558_, _27556_, _27490_);
  or (_27559_, _27558_, _03059_);
  and (_27560_, _27559_, _03061_);
  and (_27561_, _27560_, _27555_);
  and (_27562_, _11588_, _03856_);
  nor (_27563_, _27562_, _27490_);
  nor (_27564_, _27563_, _03061_);
  nor (_27565_, _27564_, _27561_);
  nor (_27566_, _27565_, _02206_);
  nor (_27567_, _27490_, _04420_);
  not (_27569_, _27567_);
  nor (_27570_, _27493_, _02208_);
  and (_27571_, _27570_, _27569_);
  nor (_27572_, _27571_, _27566_);
  nor (_27573_, _27572_, _02342_);
  or (_27574_, _27567_, _03065_);
  nor (_27575_, _27574_, _27499_);
  or (_27576_, _27575_, _02202_);
  nor (_27577_, _27576_, _27573_);
  nor (_27578_, _11590_, _09607_);
  or (_27580_, _27490_, _04953_);
  nor (_27581_, _27580_, _27578_);
  or (_27582_, _27581_, _02334_);
  nor (_27583_, _27582_, _27577_);
  nor (_27584_, _11587_, _09607_);
  nor (_27585_, _27584_, _27490_);
  nor (_27586_, _27585_, _04958_);
  or (_27587_, _27586_, _27583_);
  and (_27588_, _27587_, _02778_);
  nor (_27589_, _27506_, _02778_);
  or (_27591_, _27589_, _27588_);
  and (_27592_, _27591_, _01698_);
  nor (_27593_, _27524_, _01698_);
  or (_27594_, _27593_, _27592_);
  and (_27595_, _27594_, _02082_);
  and (_27596_, _11771_, _03856_);
  nor (_27597_, _27596_, _27490_);
  nor (_27598_, _27597_, _02082_);
  or (_27599_, _27598_, _27595_);
  or (_27600_, _27599_, _39633_);
  or (_27602_, _39632_, \oc8051_golden_model_1.TCON [4]);
  and (_27603_, _27602_, _39026_);
  and (_41746_, _27603_, _27600_);
  not (_27604_, \oc8051_golden_model_1.TCON [5]);
  nor (_27605_, _03856_, _27604_);
  and (_27606_, _04827_, _03856_);
  nor (_27607_, _27606_, _27605_);
  and (_27608_, _27607_, _01994_);
  nor (_27609_, _04057_, _09607_);
  nor (_27610_, _27609_, _27605_);
  and (_27612_, _27610_, _06188_);
  and (_27613_, _03856_, \oc8051_golden_model_1.ACC [5]);
  nor (_27614_, _27613_, _27605_);
  nor (_27615_, _27614_, _02063_);
  nor (_27616_, _02062_, _27604_);
  or (_27617_, _27616_, _27615_);
  and (_27618_, _27617_, _03006_);
  nor (_27619_, _11804_, _09607_);
  nor (_27620_, _27619_, _27605_);
  nor (_27621_, _27620_, _03006_);
  or (_27623_, _27621_, _27618_);
  and (_27624_, _27623_, _02058_);
  nor (_27625_, _04487_, _27604_);
  and (_27626_, _11789_, _04487_);
  nor (_27627_, _27626_, _27625_);
  nor (_27628_, _27627_, _02058_);
  or (_27629_, _27628_, _27624_);
  and (_27630_, _27629_, _02519_);
  nor (_27631_, _27610_, _02519_);
  or (_27632_, _27631_, _27630_);
  and (_27634_, _27632_, _02549_);
  nor (_27635_, _27614_, _02549_);
  or (_27636_, _27635_, _27634_);
  and (_27637_, _27636_, _02054_);
  and (_27638_, _11816_, _04487_);
  nor (_27639_, _27638_, _27625_);
  nor (_27640_, _27639_, _02054_);
  or (_27641_, _27640_, _27637_);
  and (_27642_, _27641_, _02047_);
  nor (_27643_, _27625_, _11823_);
  nor (_27645_, _27643_, _27627_);
  and (_27646_, _27645_, _02046_);
  or (_27647_, _27646_, _27642_);
  and (_27648_, _27647_, _02043_);
  nor (_27649_, _11841_, _09644_);
  nor (_27650_, _27649_, _27625_);
  nor (_27651_, _27650_, _02043_);
  nor (_27652_, _27651_, _06188_);
  not (_27653_, _27652_);
  nor (_27654_, _27653_, _27648_);
  nor (_27656_, _27654_, _27612_);
  nor (_27657_, _27656_, _02031_);
  and (_27658_, _05258_, _03856_);
  nor (_27659_, _27605_, _02032_);
  not (_27660_, _27659_);
  nor (_27661_, _27660_, _27658_);
  or (_27662_, _27661_, _01765_);
  nor (_27663_, _27662_, _27657_);
  nor (_27664_, _11900_, _09607_);
  nor (_27665_, _27664_, _27605_);
  nor (_27667_, _27665_, _02037_);
  or (_27668_, _27667_, _01994_);
  nor (_27669_, _27668_, _27663_);
  nor (_27670_, _27669_, _27608_);
  or (_27671_, _27670_, _02210_);
  and (_27672_, _11915_, _03856_);
  or (_27673_, _27672_, _27605_);
  or (_27674_, _27673_, _03059_);
  and (_27675_, _27674_, _03061_);
  and (_27676_, _27675_, _27671_);
  and (_27678_, _11786_, _03856_);
  nor (_27679_, _27678_, _27605_);
  nor (_27680_, _27679_, _03061_);
  nor (_27681_, _27680_, _27676_);
  nor (_27682_, _27681_, _02206_);
  nor (_27683_, _27605_, _04104_);
  not (_27684_, _27683_);
  nor (_27685_, _27607_, _02208_);
  and (_27686_, _27685_, _27684_);
  nor (_27687_, _27686_, _27682_);
  nor (_27689_, _27687_, _02342_);
  or (_27690_, _27683_, _03065_);
  nor (_27691_, _27690_, _27614_);
  or (_27692_, _27691_, _02202_);
  nor (_27693_, _27692_, _27689_);
  nor (_27694_, _11913_, _09607_);
  or (_27695_, _27605_, _04953_);
  nor (_27696_, _27695_, _27694_);
  or (_27697_, _27696_, _02334_);
  nor (_27698_, _27697_, _27693_);
  nor (_27700_, _11785_, _09607_);
  nor (_27701_, _27700_, _27605_);
  nor (_27702_, _27701_, _04958_);
  or (_27703_, _27702_, _27698_);
  and (_27704_, _27703_, _02778_);
  nor (_27705_, _27620_, _02778_);
  or (_27706_, _27705_, _27704_);
  and (_27707_, _27706_, _01698_);
  nor (_27708_, _27639_, _01698_);
  or (_27709_, _27708_, _27707_);
  and (_27711_, _27709_, _02082_);
  and (_27712_, _11974_, _03856_);
  nor (_27713_, _27712_, _27605_);
  nor (_27714_, _27713_, _02082_);
  or (_27715_, _27714_, _27711_);
  or (_27716_, _27715_, _39633_);
  or (_27717_, _39632_, \oc8051_golden_model_1.TCON [5]);
  and (_27718_, _27717_, _39026_);
  and (_41747_, _27718_, _27716_);
  not (_27719_, \oc8051_golden_model_1.TCON [6]);
  nor (_27720_, _03856_, _27719_);
  and (_27721_, _12103_, _03856_);
  nor (_27722_, _27721_, _27720_);
  and (_27723_, _27722_, _01994_);
  nor (_27724_, _03964_, _09607_);
  nor (_27725_, _27724_, _27720_);
  and (_27726_, _27725_, _06188_);
  and (_27727_, _03856_, \oc8051_golden_model_1.ACC [6]);
  nor (_27728_, _27727_, _27720_);
  nor (_27729_, _27728_, _02063_);
  nor (_27731_, _02062_, _27719_);
  or (_27732_, _27731_, _27729_);
  and (_27733_, _27732_, _03006_);
  nor (_27734_, _11993_, _09607_);
  nor (_27735_, _27734_, _27720_);
  nor (_27736_, _27735_, _03006_);
  or (_27737_, _27736_, _27733_);
  and (_27738_, _27737_, _02058_);
  nor (_27739_, _04487_, _27719_);
  and (_27740_, _11990_, _04487_);
  nor (_27742_, _27740_, _27739_);
  nor (_27743_, _27742_, _02058_);
  or (_27744_, _27743_, _27738_);
  and (_27745_, _27744_, _02519_);
  nor (_27746_, _27725_, _02519_);
  or (_27747_, _27746_, _27745_);
  and (_27748_, _27747_, _02549_);
  nor (_27749_, _27728_, _02549_);
  or (_27750_, _27749_, _27748_);
  and (_27751_, _27750_, _02054_);
  and (_27753_, _12017_, _04487_);
  nor (_27754_, _27753_, _27739_);
  nor (_27755_, _27754_, _02054_);
  or (_27756_, _27755_, _27751_);
  and (_27757_, _27756_, _02047_);
  nor (_27758_, _27739_, _12024_);
  nor (_27759_, _27758_, _27742_);
  and (_27760_, _27759_, _02046_);
  or (_27761_, _27760_, _27757_);
  and (_27762_, _27761_, _02043_);
  nor (_27764_, _12042_, _09644_);
  nor (_27765_, _27764_, _27739_);
  nor (_27766_, _27765_, _02043_);
  nor (_27767_, _27766_, _06188_);
  not (_27768_, _27767_);
  nor (_27769_, _27768_, _27762_);
  nor (_27770_, _27769_, _27726_);
  nor (_27771_, _27770_, _02031_);
  and (_27772_, _05029_, _03856_);
  nor (_27773_, _27720_, _02032_);
  not (_27775_, _27773_);
  nor (_27776_, _27775_, _27772_);
  or (_27777_, _27776_, _01765_);
  nor (_27778_, _27777_, _27771_);
  nor (_27779_, _12096_, _09607_);
  nor (_27780_, _27779_, _27720_);
  nor (_27781_, _27780_, _02037_);
  or (_27782_, _27781_, _01994_);
  nor (_27783_, _27782_, _27778_);
  nor (_27784_, _27783_, _27723_);
  or (_27786_, _27784_, _02210_);
  and (_27787_, _12112_, _03856_);
  or (_27788_, _27787_, _27720_);
  or (_27789_, _27788_, _03059_);
  and (_27790_, _27789_, _03061_);
  and (_27791_, _27790_, _27786_);
  and (_27792_, _12118_, _03856_);
  nor (_27793_, _27792_, _27720_);
  nor (_27794_, _27793_, _03061_);
  nor (_27795_, _27794_, _27791_);
  nor (_27797_, _27795_, _02206_);
  nor (_27798_, _27720_, _04011_);
  not (_27799_, _27798_);
  nor (_27800_, _27722_, _02208_);
  and (_27801_, _27800_, _27799_);
  nor (_27802_, _27801_, _27797_);
  nor (_27803_, _27802_, _02342_);
  or (_27804_, _27798_, _03065_);
  nor (_27805_, _27804_, _27728_);
  or (_27806_, _27805_, _02202_);
  nor (_27808_, _27806_, _27803_);
  nor (_27809_, _12110_, _09607_);
  or (_27810_, _27720_, _04953_);
  nor (_27811_, _27810_, _27809_);
  or (_27812_, _27811_, _02334_);
  nor (_27813_, _27812_, _27808_);
  nor (_27814_, _12117_, _09607_);
  nor (_27815_, _27814_, _27720_);
  nor (_27816_, _27815_, _04958_);
  or (_27817_, _27816_, _27813_);
  and (_27819_, _27817_, _02778_);
  nor (_27820_, _27735_, _02778_);
  or (_27821_, _27820_, _27819_);
  and (_27822_, _27821_, _01698_);
  nor (_27823_, _27754_, _01698_);
  or (_27824_, _27823_, _27822_);
  and (_27825_, _27824_, _02082_);
  and (_27826_, _12178_, _03856_);
  nor (_27827_, _27826_, _27720_);
  nor (_27828_, _27827_, _02082_);
  or (_27830_, _27828_, _27825_);
  or (_27831_, _27830_, _39633_);
  or (_27832_, _39632_, \oc8051_golden_model_1.TCON [6]);
  and (_27833_, _27832_, _39026_);
  and (_41748_, _27833_, _27831_);
  not (_27834_, \oc8051_golden_model_1.TH0 [0]);
  nor (_27835_, _03854_, _27834_);
  nor (_27836_, _04257_, _09714_);
  nor (_27837_, _27836_, _27835_);
  and (_27838_, _27837_, _15890_);
  and (_27840_, _03854_, _04837_);
  nor (_27841_, _27840_, _27835_);
  nor (_27842_, _27841_, _02208_);
  not (_27843_, _27842_);
  nor (_27844_, _27843_, _27836_);
  and (_27845_, _03854_, \oc8051_golden_model_1.ACC [0]);
  nor (_27846_, _27845_, _27835_);
  nor (_27847_, _27846_, _02549_);
  nor (_27848_, _27847_, _06188_);
  nor (_27849_, _27837_, _03006_);
  nor (_27851_, _02062_, _27834_);
  nor (_27852_, _27846_, _02063_);
  nor (_27853_, _27852_, _27851_);
  nor (_27854_, _27853_, _02158_);
  or (_27855_, _27854_, _02155_);
  nor (_27856_, _27855_, _27849_);
  or (_27857_, _27856_, _02153_);
  and (_27858_, _27857_, _27848_);
  and (_27859_, _03854_, _03002_);
  or (_27860_, _27835_, _24237_);
  nor (_27862_, _27860_, _27859_);
  nor (_27863_, _27862_, _27858_);
  nor (_27864_, _27863_, _02031_);
  and (_27865_, _05120_, _03854_);
  nor (_27866_, _27835_, _02032_);
  not (_27867_, _27866_);
  nor (_27868_, _27867_, _27865_);
  nor (_27869_, _27868_, _27864_);
  nor (_27870_, _27869_, _01765_);
  nor (_27871_, _10898_, _09714_);
  or (_27873_, _27835_, _02037_);
  nor (_27874_, _27873_, _27871_);
  or (_27875_, _27874_, _01994_);
  nor (_27876_, _27875_, _27870_);
  nand (_27877_, _27841_, _03059_);
  and (_27878_, _27877_, _07629_);
  nor (_27879_, _27878_, _27876_);
  and (_27880_, _10914_, _03854_);
  nor (_27881_, _27880_, _27835_);
  and (_27882_, _27881_, _02210_);
  nor (_27884_, _27882_, _27879_);
  and (_27885_, _27884_, _03061_);
  and (_27886_, _10792_, _03854_);
  nor (_27887_, _27886_, _27835_);
  nor (_27888_, _27887_, _03061_);
  or (_27889_, _27888_, _27885_);
  and (_27890_, _27889_, _02208_);
  nor (_27891_, _27890_, _27844_);
  nor (_27892_, _27891_, _02342_);
  and (_27893_, _10791_, _03854_);
  or (_27895_, _27893_, _27835_);
  and (_27896_, _27895_, _02342_);
  or (_27897_, _27896_, _27892_);
  and (_27898_, _27897_, _04953_);
  nor (_27899_, _10913_, _09714_);
  nor (_27900_, _27899_, _27835_);
  nor (_27901_, _27900_, _04953_);
  or (_27902_, _27901_, _27898_);
  and (_27903_, _27902_, _04958_);
  nor (_27904_, _10789_, _09714_);
  nor (_27906_, _27904_, _27835_);
  nor (_27907_, _27906_, _04958_);
  nor (_27908_, _27907_, _15890_);
  not (_27909_, _27908_);
  nor (_27910_, _27909_, _27903_);
  nor (_27911_, _27910_, _27838_);
  or (_27912_, _27911_, _39633_);
  or (_27913_, _39632_, \oc8051_golden_model_1.TH0 [0]);
  and (_27914_, _27913_, _39026_);
  and (_41750_, _27914_, _27912_);
  nor (_27915_, _03854_, \oc8051_golden_model_1.TH0 [1]);
  not (_27916_, _27915_);
  nor (_27917_, _10988_, _09714_);
  nor (_27918_, _27917_, _02208_);
  and (_27919_, _27918_, _27916_);
  nor (_27920_, _11113_, _09714_);
  nor (_27921_, _27920_, _03061_);
  and (_27922_, _27921_, _27916_);
  and (_27923_, _05075_, _03854_);
  not (_27924_, \oc8051_golden_model_1.TH0 [1]);
  nor (_27926_, _03854_, _27924_);
  nor (_27927_, _27926_, _02032_);
  not (_27928_, _27927_);
  nor (_27929_, _27928_, _27923_);
  not (_27930_, _27929_);
  and (_27931_, _03854_, _01804_);
  nor (_27932_, _27931_, _27915_);
  and (_27933_, _27932_, _02153_);
  and (_27934_, _27932_, _02062_);
  nor (_27935_, _02062_, _27924_);
  or (_27937_, _27935_, _27934_);
  and (_27938_, _27937_, _03006_);
  and (_27939_, _11001_, _03854_);
  nor (_27940_, _27939_, _27915_);
  and (_27941_, _27940_, _02158_);
  or (_27942_, _27941_, _27938_);
  and (_27943_, _27942_, _02519_);
  nor (_27944_, _09714_, _03161_);
  nor (_27945_, _27944_, _27926_);
  nor (_27946_, _27945_, _02519_);
  nor (_27948_, _27946_, _27943_);
  nor (_27949_, _27948_, _02153_);
  or (_27950_, _27949_, _06188_);
  nor (_27951_, _27950_, _27933_);
  and (_27952_, _27945_, _06188_);
  nor (_27953_, _27952_, _27951_);
  nor (_27954_, _27953_, _02031_);
  nor (_27955_, _27954_, _01765_);
  and (_27956_, _27955_, _27930_);
  and (_27957_, _11096_, _03854_);
  nor (_27959_, _27957_, _02037_);
  and (_27960_, _27959_, _27916_);
  nor (_27961_, _27960_, _27956_);
  nor (_27962_, _27961_, _07629_);
  nor (_27963_, _10989_, _09714_);
  nor (_27964_, _27963_, _03059_);
  and (_27965_, _03854_, _02893_);
  nor (_27966_, _27965_, _01995_);
  nor (_27967_, _27966_, _27964_);
  nor (_27968_, _27967_, _27915_);
  nor (_27970_, _27968_, _27962_);
  nor (_27971_, _27970_, _02331_);
  nor (_27972_, _27971_, _27922_);
  nor (_27973_, _27972_, _02206_);
  nor (_27974_, _27973_, _27919_);
  nor (_27975_, _27974_, _02342_);
  nor (_27976_, _27926_, _04209_);
  nor (_27977_, _27976_, _03065_);
  and (_27978_, _27977_, _27932_);
  nor (_27979_, _27978_, _27975_);
  or (_27981_, _27979_, _17216_);
  nand (_27982_, _27931_, _04208_);
  nor (_27983_, _27915_, _04958_);
  and (_27984_, _27983_, _27982_);
  nor (_27985_, _27984_, _02366_);
  and (_27986_, _27965_, _04208_);
  or (_27987_, _27915_, _04953_);
  or (_27988_, _27987_, _27986_);
  and (_27989_, _27988_, _27985_);
  and (_27990_, _27989_, _27981_);
  nor (_27992_, _27940_, _02778_);
  nor (_27993_, _27992_, _27990_);
  nor (_27994_, _27993_, _02081_);
  nor (_27995_, _27939_, _27926_);
  and (_27996_, _27995_, _02081_);
  nor (_27997_, _27996_, _27994_);
  or (_27998_, _27997_, _39633_);
  or (_27999_, _39632_, \oc8051_golden_model_1.TH0 [1]);
  and (_28000_, _27999_, _39026_);
  and (_41751_, _28000_, _27998_);
  not (_28002_, \oc8051_golden_model_1.TH0 [2]);
  nor (_28003_, _03854_, _28002_);
  nor (_28004_, _11314_, _09714_);
  nor (_28005_, _28004_, _28003_);
  nor (_28006_, _28005_, _04958_);
  nor (_28007_, _09714_, _03624_);
  nor (_28008_, _28007_, _28003_);
  and (_28009_, _28008_, _06188_);
  and (_28010_, _03854_, \oc8051_golden_model_1.ACC [2]);
  nor (_28011_, _28010_, _28003_);
  nor (_28013_, _28011_, _02063_);
  nor (_28014_, _02062_, _28002_);
  or (_28015_, _28014_, _28013_);
  and (_28016_, _28015_, _03006_);
  nor (_28017_, _11199_, _09714_);
  nor (_28018_, _28017_, _28003_);
  nor (_28019_, _28018_, _03006_);
  or (_28020_, _28019_, _28016_);
  and (_28021_, _28020_, _02519_);
  nor (_28022_, _28008_, _02519_);
  nor (_28024_, _28022_, _28021_);
  nor (_28025_, _28024_, _02153_);
  nor (_28026_, _28011_, _02549_);
  nor (_28027_, _28026_, _06188_);
  not (_28028_, _28027_);
  nor (_28029_, _28028_, _28025_);
  nor (_28030_, _28029_, _28009_);
  nor (_28031_, _28030_, _02031_);
  and (_28032_, _05211_, _03854_);
  nor (_28033_, _28003_, _02032_);
  not (_28035_, _28033_);
  nor (_28036_, _28035_, _28032_);
  nor (_28037_, _28036_, _28031_);
  nor (_28038_, _28037_, _01765_);
  nor (_28039_, _11298_, _09714_);
  or (_28040_, _28003_, _02037_);
  nor (_28041_, _28040_, _28039_);
  or (_28042_, _28041_, _01994_);
  nor (_28043_, _28042_, _28038_);
  and (_28044_, _03854_, _04866_);
  nor (_28046_, _28044_, _28003_);
  nand (_28047_, _28046_, _03059_);
  and (_28048_, _28047_, _07629_);
  nor (_28049_, _28048_, _28043_);
  and (_28050_, _11189_, _03854_);
  nor (_28051_, _28050_, _28003_);
  and (_28052_, _28051_, _02210_);
  nor (_28053_, _28052_, _28049_);
  and (_28054_, _28053_, _03061_);
  and (_28055_, _11315_, _03854_);
  nor (_28057_, _28055_, _28003_);
  nor (_28058_, _28057_, _03061_);
  or (_28059_, _28058_, _28054_);
  and (_28060_, _28059_, _02208_);
  nor (_28061_, _28003_, _04309_);
  not (_28062_, _28061_);
  nor (_28063_, _28046_, _02208_);
  and (_28064_, _28063_, _28062_);
  nor (_28065_, _28064_, _28060_);
  nor (_28066_, _28065_, _02342_);
  or (_28068_, _28061_, _03065_);
  nor (_28069_, _28068_, _28011_);
  or (_28070_, _28069_, _02202_);
  nor (_28071_, _28070_, _28066_);
  nor (_28072_, _11187_, _09714_);
  or (_28073_, _28003_, _04953_);
  nor (_28074_, _28073_, _28072_);
  or (_28075_, _28074_, _02334_);
  nor (_28076_, _28075_, _28071_);
  nor (_28077_, _28076_, _28006_);
  nor (_28079_, _28077_, _02366_);
  nor (_28080_, _28018_, _02778_);
  or (_28081_, _28080_, _02081_);
  nor (_28082_, _28081_, _28079_);
  and (_28083_, _11367_, _03854_);
  nor (_28084_, _28083_, _28003_);
  and (_28085_, _28084_, _02081_);
  nor (_28086_, _28085_, _28082_);
  or (_28087_, _28086_, _39633_);
  or (_28088_, _39632_, \oc8051_golden_model_1.TH0 [2]);
  and (_28090_, _28088_, _39026_);
  and (_41752_, _28090_, _28087_);
  not (_28091_, \oc8051_golden_model_1.TH0 [3]);
  nor (_28092_, _03854_, _28091_);
  nor (_28093_, _11510_, _09714_);
  nor (_28094_, _28093_, _28092_);
  nor (_28095_, _28094_, _04958_);
  and (_28096_, _11511_, _03854_);
  nor (_28097_, _28096_, _28092_);
  nor (_28098_, _28097_, _03061_);
  and (_28100_, _03854_, \oc8051_golden_model_1.ACC [3]);
  nor (_28101_, _28100_, _28092_);
  nor (_28102_, _28101_, _02549_);
  nor (_28103_, _28101_, _02063_);
  nor (_28104_, _02062_, _28091_);
  or (_28105_, _28104_, _28103_);
  and (_28106_, _28105_, _03006_);
  nor (_28107_, _11394_, _09714_);
  nor (_28108_, _28107_, _28092_);
  nor (_28109_, _28108_, _03006_);
  or (_28111_, _28109_, _28106_);
  and (_28112_, _28111_, _02519_);
  nor (_28113_, _09714_, _03434_);
  nor (_28114_, _28113_, _28092_);
  nor (_28115_, _28114_, _02519_);
  nor (_28116_, _28115_, _28112_);
  nor (_28117_, _28116_, _02153_);
  or (_28118_, _28117_, _06188_);
  nor (_28119_, _28118_, _28102_);
  and (_28120_, _28114_, _06188_);
  nor (_28122_, _28120_, _28119_);
  nor (_28123_, _28122_, _02031_);
  and (_28124_, _05166_, _03854_);
  nor (_28125_, _28092_, _02032_);
  not (_28126_, _28125_);
  nor (_28127_, _28126_, _28124_);
  nor (_28128_, _28127_, _01765_);
  not (_28129_, _28128_);
  nor (_28130_, _28129_, _28123_);
  nor (_28131_, _11490_, _09714_);
  nor (_28132_, _28131_, _28092_);
  nor (_28133_, _28132_, _02037_);
  or (_28134_, _28133_, _07629_);
  or (_28135_, _28134_, _28130_);
  and (_28136_, _11505_, _03854_);
  or (_28137_, _28092_, _03059_);
  or (_28138_, _28137_, _28136_);
  and (_28139_, _03854_, _04719_);
  nor (_28140_, _28139_, _28092_);
  and (_28141_, _28140_, _01994_);
  nor (_28143_, _28141_, _02331_);
  and (_28144_, _28143_, _28138_);
  and (_28145_, _28144_, _28135_);
  nor (_28146_, _28145_, _28098_);
  nor (_28147_, _28146_, _02206_);
  nor (_28148_, _28092_, _04153_);
  not (_28149_, _28148_);
  nor (_28150_, _28140_, _02208_);
  and (_28151_, _28150_, _28149_);
  nor (_28152_, _28151_, _28147_);
  nor (_28154_, _28152_, _02342_);
  or (_28155_, _28148_, _03065_);
  nor (_28156_, _28155_, _28101_);
  or (_28157_, _28156_, _02202_);
  nor (_28158_, _28157_, _28154_);
  nor (_28159_, _11503_, _09714_);
  or (_28160_, _28092_, _04953_);
  nor (_28161_, _28160_, _28159_);
  or (_28162_, _28161_, _02334_);
  nor (_28163_, _28162_, _28158_);
  nor (_28165_, _28163_, _28095_);
  nor (_28166_, _28165_, _02366_);
  nor (_28167_, _28108_, _02778_);
  or (_28168_, _28167_, _02081_);
  nor (_28169_, _28168_, _28166_);
  and (_28170_, _11567_, _03854_);
  nor (_28171_, _28170_, _28092_);
  and (_28172_, _28171_, _02081_);
  nor (_28173_, _28172_, _28169_);
  or (_28174_, _28173_, _39633_);
  or (_28176_, _39632_, \oc8051_golden_model_1.TH0 [3]);
  and (_28177_, _28176_, _39026_);
  and (_41753_, _28177_, _28174_);
  not (_28178_, \oc8051_golden_model_1.TH0 [4]);
  nor (_28179_, _03854_, _28178_);
  nor (_28180_, _11587_, _09714_);
  nor (_28181_, _28180_, _28179_);
  nor (_28182_, _28181_, _04958_);
  nor (_28183_, _28179_, _04420_);
  not (_28184_, _28183_);
  and (_28186_, _04831_, _03854_);
  nor (_28187_, _28186_, _28179_);
  nor (_28188_, _28187_, _02208_);
  and (_28189_, _28188_, _28184_);
  and (_28190_, _11588_, _03854_);
  nor (_28191_, _28190_, _28179_);
  nor (_28192_, _28191_, _03061_);
  and (_28193_, _05303_, _03854_);
  or (_28194_, _28193_, _28179_);
  and (_28195_, _28194_, _02031_);
  and (_28197_, _03854_, \oc8051_golden_model_1.ACC [4]);
  nor (_28198_, _28197_, _28179_);
  nor (_28199_, _28198_, _02549_);
  nor (_28200_, _28198_, _02063_);
  nor (_28201_, _02062_, _28178_);
  or (_28202_, _28201_, _28200_);
  and (_28203_, _28202_, _03006_);
  nor (_28204_, _11611_, _09714_);
  nor (_28205_, _28204_, _28179_);
  nor (_28206_, _28205_, _03006_);
  or (_28208_, _28206_, _28203_);
  and (_28209_, _28208_, _02519_);
  nor (_28210_, _04372_, _09714_);
  nor (_28211_, _28210_, _28179_);
  nor (_28212_, _28211_, _02519_);
  nor (_28213_, _28212_, _28209_);
  nor (_28214_, _28213_, _02153_);
  or (_28215_, _28214_, _06188_);
  nor (_28216_, _28215_, _28199_);
  and (_28217_, _28211_, _06188_);
  or (_28219_, _28217_, _02031_);
  nor (_28220_, _28219_, _28216_);
  or (_28221_, _28220_, _28195_);
  and (_28222_, _28221_, _02037_);
  nor (_28223_, _11704_, _09714_);
  nor (_28224_, _28223_, _28179_);
  nor (_28225_, _28224_, _02037_);
  or (_28226_, _28225_, _07629_);
  or (_28227_, _28226_, _28222_);
  and (_28228_, _11592_, _03854_);
  or (_28230_, _28179_, _03059_);
  or (_28231_, _28230_, _28228_);
  and (_28232_, _28187_, _01994_);
  nor (_28233_, _28232_, _02331_);
  and (_28234_, _28233_, _28231_);
  and (_28235_, _28234_, _28227_);
  nor (_28236_, _28235_, _28192_);
  nor (_28237_, _28236_, _02206_);
  nor (_28238_, _28237_, _28189_);
  nor (_28239_, _28238_, _02342_);
  or (_28241_, _28183_, _03065_);
  nor (_28242_, _28241_, _28198_);
  or (_28243_, _28242_, _02202_);
  nor (_28244_, _28243_, _28239_);
  nor (_28245_, _11590_, _09714_);
  or (_28246_, _28179_, _04953_);
  nor (_28247_, _28246_, _28245_);
  or (_28248_, _28247_, _02334_);
  nor (_28249_, _28248_, _28244_);
  nor (_28250_, _28249_, _28182_);
  nor (_28252_, _28250_, _02366_);
  nor (_28253_, _28205_, _02778_);
  or (_28254_, _28253_, _02081_);
  nor (_28255_, _28254_, _28252_);
  and (_28256_, _11771_, _03854_);
  nor (_28257_, _28256_, _28179_);
  and (_28258_, _28257_, _02081_);
  nor (_28259_, _28258_, _28255_);
  or (_28260_, _28259_, _39633_);
  or (_28261_, _39632_, \oc8051_golden_model_1.TH0 [4]);
  and (_28262_, _28261_, _39026_);
  and (_41754_, _28262_, _28260_);
  not (_28263_, \oc8051_golden_model_1.TH0 [5]);
  nor (_28264_, _03854_, _28263_);
  nor (_28265_, _11785_, _09714_);
  nor (_28266_, _28265_, _28264_);
  nor (_28267_, _28266_, _04958_);
  and (_28268_, _11786_, _03854_);
  nor (_28269_, _28268_, _28264_);
  nor (_28270_, _28269_, _03061_);
  and (_28272_, _04827_, _03854_);
  nor (_28273_, _28272_, _28264_);
  and (_28274_, _28273_, _01994_);
  and (_28275_, _03854_, \oc8051_golden_model_1.ACC [5]);
  nor (_28276_, _28275_, _28264_);
  nor (_28277_, _28276_, _02549_);
  nor (_28278_, _28276_, _02063_);
  nor (_28279_, _02062_, _28263_);
  or (_28280_, _28279_, _28278_);
  and (_28281_, _28280_, _03006_);
  nor (_28283_, _11804_, _09714_);
  nor (_28284_, _28283_, _28264_);
  nor (_28285_, _28284_, _03006_);
  or (_28286_, _28285_, _28281_);
  and (_28287_, _28286_, _02519_);
  nor (_28288_, _04057_, _09714_);
  nor (_28289_, _28288_, _28264_);
  nor (_28290_, _28289_, _02519_);
  nor (_28291_, _28290_, _28287_);
  nor (_28292_, _28291_, _02153_);
  or (_28294_, _28292_, _06188_);
  nor (_28295_, _28294_, _28277_);
  and (_28296_, _28289_, _06188_);
  nor (_28297_, _28296_, _28295_);
  nor (_28298_, _28297_, _02031_);
  and (_28299_, _05258_, _03854_);
  nor (_28300_, _28264_, _02032_);
  not (_28301_, _28300_);
  nor (_28302_, _28301_, _28299_);
  or (_28303_, _28302_, _01765_);
  nor (_28305_, _28303_, _28298_);
  nor (_28306_, _11900_, _09714_);
  nor (_28307_, _28306_, _28264_);
  nor (_28308_, _28307_, _02037_);
  or (_28309_, _28308_, _01994_);
  nor (_28310_, _28309_, _28305_);
  nor (_28311_, _28310_, _28274_);
  or (_28312_, _28311_, _02210_);
  and (_28313_, _11915_, _03854_);
  or (_28314_, _28313_, _28264_);
  or (_28316_, _28314_, _03059_);
  and (_28317_, _28316_, _03061_);
  and (_28318_, _28317_, _28312_);
  nor (_28319_, _28318_, _28270_);
  nor (_28320_, _28319_, _02206_);
  nor (_28321_, _28264_, _04104_);
  not (_28322_, _28321_);
  nor (_28323_, _28273_, _02208_);
  and (_28324_, _28323_, _28322_);
  nor (_28325_, _28324_, _28320_);
  nor (_28327_, _28325_, _02342_);
  or (_28328_, _28321_, _03065_);
  nor (_28329_, _28328_, _28276_);
  or (_28330_, _28329_, _02202_);
  nor (_28331_, _28330_, _28327_);
  nor (_28332_, _11913_, _09714_);
  or (_28333_, _28264_, _04953_);
  nor (_28334_, _28333_, _28332_);
  or (_28335_, _28334_, _02334_);
  nor (_28336_, _28335_, _28331_);
  nor (_28338_, _28336_, _28267_);
  nor (_28339_, _28338_, _02366_);
  nor (_28340_, _28284_, _02778_);
  or (_28341_, _28340_, _02081_);
  nor (_28342_, _28341_, _28339_);
  and (_28343_, _11974_, _03854_);
  nor (_28344_, _28343_, _28264_);
  and (_28345_, _28344_, _02081_);
  nor (_28346_, _28345_, _28342_);
  or (_28347_, _28346_, _39633_);
  or (_28349_, _39632_, \oc8051_golden_model_1.TH0 [5]);
  and (_28350_, _28349_, _39026_);
  and (_41755_, _28350_, _28347_);
  not (_28351_, \oc8051_golden_model_1.TH0 [6]);
  nor (_28352_, _03854_, _28351_);
  nor (_28353_, _12117_, _09714_);
  nor (_28354_, _28353_, _28352_);
  nor (_28355_, _28354_, _04958_);
  and (_28356_, _12118_, _03854_);
  nor (_28357_, _28356_, _28352_);
  nor (_28359_, _28357_, _03061_);
  and (_28360_, _12103_, _03854_);
  nor (_28361_, _28360_, _28352_);
  and (_28362_, _28361_, _01994_);
  nor (_28363_, _03964_, _09714_);
  nor (_28364_, _28363_, _28352_);
  and (_28365_, _28364_, _06188_);
  and (_28366_, _03854_, \oc8051_golden_model_1.ACC [6]);
  nor (_28367_, _28366_, _28352_);
  nor (_28368_, _28367_, _02063_);
  nor (_28370_, _02062_, _28351_);
  or (_28371_, _28370_, _28368_);
  and (_28372_, _28371_, _03006_);
  nor (_28373_, _11993_, _09714_);
  nor (_28374_, _28373_, _28352_);
  nor (_28375_, _28374_, _03006_);
  or (_28376_, _28375_, _28372_);
  and (_28377_, _28376_, _02519_);
  nor (_28378_, _28364_, _02519_);
  nor (_28379_, _28378_, _28377_);
  nor (_28381_, _28379_, _02153_);
  nor (_28382_, _28367_, _02549_);
  nor (_28383_, _28382_, _06188_);
  not (_28384_, _28383_);
  nor (_28385_, _28384_, _28381_);
  nor (_28386_, _28385_, _28365_);
  nor (_28387_, _28386_, _02031_);
  and (_28388_, _05029_, _03854_);
  nor (_28389_, _28352_, _02032_);
  not (_28390_, _28389_);
  nor (_28391_, _28390_, _28388_);
  or (_28392_, _28391_, _01765_);
  nor (_28393_, _28392_, _28387_);
  nor (_28394_, _12096_, _09714_);
  nor (_28395_, _28394_, _28352_);
  nor (_28396_, _28395_, _02037_);
  or (_28397_, _28396_, _01994_);
  nor (_28398_, _28397_, _28393_);
  nor (_28399_, _28398_, _28362_);
  or (_28400_, _28399_, _02210_);
  and (_28402_, _12112_, _03854_);
  or (_28403_, _28402_, _28352_);
  or (_28404_, _28403_, _03059_);
  and (_28405_, _28404_, _03061_);
  and (_28406_, _28405_, _28400_);
  nor (_28407_, _28406_, _28359_);
  nor (_28408_, _28407_, _02206_);
  nor (_28409_, _28352_, _04011_);
  not (_28410_, _28409_);
  nor (_28411_, _28361_, _02208_);
  and (_28413_, _28411_, _28410_);
  nor (_28414_, _28413_, _28408_);
  nor (_28415_, _28414_, _02342_);
  or (_28416_, _28409_, _03065_);
  nor (_28417_, _28416_, _28367_);
  or (_28418_, _28417_, _02202_);
  nor (_28419_, _28418_, _28415_);
  nor (_28420_, _12110_, _09714_);
  or (_28421_, _28352_, _04953_);
  nor (_28422_, _28421_, _28420_);
  or (_28424_, _28422_, _02334_);
  nor (_28425_, _28424_, _28419_);
  nor (_28426_, _28425_, _28355_);
  nor (_28427_, _28426_, _02366_);
  nor (_28428_, _28374_, _02778_);
  or (_28429_, _28428_, _02081_);
  nor (_28430_, _28429_, _28427_);
  and (_28431_, _12178_, _03854_);
  nor (_28432_, _28431_, _28352_);
  and (_28433_, _28432_, _02081_);
  nor (_28435_, _28433_, _28430_);
  or (_28436_, _28435_, _39633_);
  or (_28437_, _39632_, \oc8051_golden_model_1.TH0 [6]);
  and (_28438_, _28437_, _39026_);
  and (_41757_, _28438_, _28436_);
  not (_28439_, \oc8051_golden_model_1.TH1 [0]);
  nor (_28440_, _03871_, _28439_);
  nor (_28441_, _04257_, _09793_);
  nor (_28442_, _28441_, _28440_);
  and (_28443_, _28442_, _15890_);
  and (_28445_, _03871_, \oc8051_golden_model_1.ACC [0]);
  nor (_28446_, _28445_, _28440_);
  nor (_28447_, _28446_, _02549_);
  nor (_28448_, _28446_, _02063_);
  nor (_28449_, _02062_, _28439_);
  or (_28450_, _28449_, _28448_);
  and (_28451_, _28450_, _03006_);
  nor (_28452_, _28442_, _03006_);
  or (_28453_, _28452_, _28451_);
  and (_28454_, _28453_, _02519_);
  and (_28456_, _03871_, _03002_);
  nor (_28457_, _28456_, _28440_);
  nor (_28458_, _28457_, _02519_);
  nor (_28459_, _28458_, _28454_);
  nor (_28460_, _28459_, _02153_);
  or (_28461_, _28460_, _06188_);
  nor (_28462_, _28461_, _28447_);
  and (_28463_, _28457_, _06188_);
  nor (_28464_, _28463_, _28462_);
  nor (_28465_, _28464_, _02031_);
  and (_28467_, _05120_, _03871_);
  nor (_28468_, _28440_, _02032_);
  not (_28469_, _28468_);
  nor (_28470_, _28469_, _28467_);
  nor (_28471_, _28470_, _28465_);
  nor (_28472_, _28471_, _01765_);
  nor (_28473_, _10898_, _09793_);
  or (_28474_, _28440_, _02037_);
  nor (_28475_, _28474_, _28473_);
  or (_28476_, _28475_, _01994_);
  nor (_28478_, _28476_, _28472_);
  and (_28479_, _03871_, _04837_);
  nor (_28480_, _28479_, _28440_);
  nand (_28481_, _28480_, _03059_);
  and (_28482_, _28481_, _07629_);
  nor (_28483_, _28482_, _28478_);
  and (_28484_, _10914_, _03871_);
  nor (_28485_, _28484_, _28440_);
  and (_28486_, _28485_, _02210_);
  nor (_28487_, _28486_, _28483_);
  and (_28489_, _28487_, _03061_);
  and (_28490_, _10792_, _03871_);
  nor (_28491_, _28490_, _28440_);
  nor (_28492_, _28491_, _03061_);
  or (_28493_, _28492_, _28489_);
  and (_28494_, _28493_, _02208_);
  or (_28495_, _28480_, _02208_);
  nor (_28496_, _28495_, _28441_);
  nor (_28497_, _28496_, _28494_);
  nor (_28498_, _28497_, _02342_);
  and (_28500_, _10791_, _03871_);
  or (_28501_, _28500_, _28440_);
  and (_28502_, _28501_, _02342_);
  or (_28503_, _28502_, _28498_);
  and (_28504_, _28503_, _04953_);
  nor (_28505_, _10913_, _09793_);
  nor (_28506_, _28505_, _28440_);
  nor (_28507_, _28506_, _04953_);
  or (_28508_, _28507_, _28504_);
  and (_28509_, _28508_, _04958_);
  nor (_28511_, _10789_, _09793_);
  nor (_28512_, _28511_, _28440_);
  nor (_28513_, _28512_, _04958_);
  nor (_28514_, _28513_, _15890_);
  not (_28515_, _28514_);
  nor (_28516_, _28515_, _28509_);
  nor (_28517_, _28516_, _28443_);
  or (_28518_, _28517_, _39633_);
  or (_28519_, _39632_, \oc8051_golden_model_1.TH1 [0]);
  and (_28520_, _28519_, _39026_);
  and (_41758_, _28520_, _28518_);
  nor (_28522_, _03871_, \oc8051_golden_model_1.TH1 [1]);
  not (_28523_, _28522_);
  nor (_28524_, _11113_, _09793_);
  nor (_28525_, _28524_, _03061_);
  and (_28526_, _28525_, _28523_);
  and (_28527_, _05075_, _03871_);
  not (_28528_, \oc8051_golden_model_1.TH1 [1]);
  nor (_28529_, _03871_, _28528_);
  nor (_28530_, _28529_, _02032_);
  not (_28531_, _28530_);
  nor (_28532_, _28531_, _28527_);
  not (_28533_, _28532_);
  and (_28534_, _03871_, _01804_);
  nor (_28535_, _28534_, _28522_);
  and (_28536_, _28535_, _02153_);
  and (_28537_, _28535_, _02062_);
  nor (_28538_, _02062_, _28528_);
  or (_28539_, _28538_, _28537_);
  and (_28540_, _28539_, _03006_);
  and (_28542_, _11001_, _03871_);
  nor (_28543_, _28542_, _28522_);
  and (_28544_, _28543_, _02158_);
  or (_28545_, _28544_, _28540_);
  and (_28546_, _28545_, _02519_);
  nor (_28547_, _09793_, _03161_);
  nor (_28548_, _28547_, _28529_);
  nor (_28549_, _28548_, _02519_);
  nor (_28550_, _28549_, _28546_);
  nor (_28551_, _28550_, _02153_);
  or (_28553_, _28551_, _06188_);
  nor (_28554_, _28553_, _28536_);
  and (_28555_, _28548_, _06188_);
  nor (_28556_, _28555_, _28554_);
  nor (_28557_, _28556_, _02031_);
  nor (_28558_, _28557_, _01765_);
  and (_28559_, _28558_, _28533_);
  and (_28560_, _11096_, _03871_);
  nor (_28561_, _28560_, _02037_);
  and (_28562_, _28561_, _28523_);
  nor (_28564_, _28562_, _28559_);
  nor (_28565_, _28564_, _07629_);
  nor (_28566_, _10989_, _09793_);
  nor (_28567_, _28566_, _03059_);
  and (_28568_, _03871_, _02893_);
  nor (_28569_, _28568_, _01995_);
  nor (_28570_, _28569_, _28567_);
  nor (_28571_, _28570_, _28522_);
  nor (_28572_, _28571_, _28565_);
  nor (_28573_, _28572_, _02331_);
  nor (_28575_, _28573_, _28526_);
  nor (_28576_, _28575_, _02206_);
  nor (_28577_, _10988_, _09793_);
  nor (_28578_, _28577_, _02208_);
  and (_28579_, _28578_, _28523_);
  nor (_28580_, _28579_, _28576_);
  nor (_28581_, _28580_, _02342_);
  nor (_28582_, _28529_, _04209_);
  nor (_28583_, _28582_, _03065_);
  and (_28584_, _28583_, _28535_);
  nor (_28586_, _28584_, _28581_);
  or (_28587_, _28586_, _17216_);
  and (_28588_, _28534_, _04208_);
  nor (_28589_, _28588_, _04958_);
  and (_28590_, _28589_, _28523_);
  nor (_28591_, _28590_, _02366_);
  and (_28592_, _28568_, _04208_);
  or (_28593_, _28522_, _04953_);
  or (_28594_, _28593_, _28592_);
  and (_28595_, _28594_, _28591_);
  and (_28597_, _28595_, _28587_);
  nor (_28598_, _28543_, _02778_);
  nor (_28599_, _28598_, _28597_);
  nor (_28600_, _28599_, _02081_);
  nor (_28601_, _28542_, _28529_);
  and (_28602_, _28601_, _02081_);
  nor (_28603_, _28602_, _28600_);
  or (_28604_, _28603_, _39633_);
  or (_28605_, _39632_, \oc8051_golden_model_1.TH1 [1]);
  and (_28606_, _28605_, _39026_);
  and (_41759_, _28606_, _28604_);
  not (_28608_, \oc8051_golden_model_1.TH1 [2]);
  nor (_28609_, _03871_, _28608_);
  nor (_28610_, _11314_, _09793_);
  nor (_28611_, _28610_, _28609_);
  nor (_28612_, _28611_, _04958_);
  nor (_28613_, _28609_, _04309_);
  not (_28614_, _28613_);
  and (_28615_, _03871_, _04866_);
  nor (_28616_, _28615_, _28609_);
  nor (_28618_, _28616_, _02208_);
  and (_28619_, _28618_, _28614_);
  and (_28620_, _11315_, _03871_);
  nor (_28621_, _28620_, _28609_);
  nor (_28622_, _28621_, _03061_);
  and (_28623_, _28616_, _01994_);
  and (_28624_, _03871_, \oc8051_golden_model_1.ACC [2]);
  nor (_28625_, _28624_, _28609_);
  nor (_28626_, _28625_, _02549_);
  nor (_28627_, _28625_, _02063_);
  nor (_28629_, _02062_, _28608_);
  or (_28630_, _28629_, _28627_);
  and (_28631_, _28630_, _03006_);
  nor (_28632_, _11199_, _09793_);
  nor (_28633_, _28632_, _28609_);
  nor (_28634_, _28633_, _03006_);
  or (_28635_, _28634_, _28631_);
  and (_28636_, _28635_, _02519_);
  nor (_28637_, _09793_, _03624_);
  nor (_28638_, _28637_, _28609_);
  nor (_28640_, _28638_, _02519_);
  nor (_28641_, _28640_, _28636_);
  nor (_28642_, _28641_, _02153_);
  or (_28643_, _28642_, _06188_);
  nor (_28644_, _28643_, _28626_);
  and (_28645_, _28638_, _06188_);
  nor (_28646_, _28645_, _28644_);
  nor (_28647_, _28646_, _02031_);
  and (_28648_, _05211_, _03871_);
  nor (_28649_, _28609_, _02032_);
  not (_28651_, _28649_);
  nor (_28652_, _28651_, _28648_);
  or (_28653_, _28652_, _01765_);
  nor (_28654_, _28653_, _28647_);
  nor (_28655_, _11298_, _09793_);
  nor (_28656_, _28655_, _28609_);
  nor (_28657_, _28656_, _02037_);
  or (_28658_, _28657_, _01994_);
  nor (_28659_, _28658_, _28654_);
  nor (_28660_, _28659_, _28623_);
  or (_28662_, _28660_, _02210_);
  and (_28663_, _11189_, _03871_);
  or (_28664_, _28663_, _28609_);
  or (_28665_, _28664_, _03059_);
  and (_28666_, _28665_, _03061_);
  and (_28667_, _28666_, _28662_);
  nor (_28668_, _28667_, _28622_);
  nor (_28669_, _28668_, _02206_);
  nor (_28670_, _28669_, _28619_);
  nor (_28671_, _28670_, _02342_);
  or (_28672_, _28613_, _03065_);
  nor (_28673_, _28672_, _28625_);
  or (_28674_, _28673_, _02202_);
  nor (_28675_, _28674_, _28671_);
  nor (_28676_, _11187_, _09793_);
  or (_28677_, _28609_, _04953_);
  nor (_28678_, _28677_, _28676_);
  or (_28679_, _28678_, _02334_);
  nor (_28680_, _28679_, _28675_);
  nor (_28681_, _28680_, _28612_);
  nor (_28683_, _28681_, _02366_);
  nor (_28684_, _28633_, _02778_);
  or (_28685_, _28684_, _02081_);
  nor (_28686_, _28685_, _28683_);
  and (_28687_, _11367_, _03871_);
  nor (_28688_, _28687_, _28609_);
  and (_28689_, _28688_, _02081_);
  nor (_28690_, _28689_, _28686_);
  or (_28691_, _28690_, _39633_);
  or (_28692_, _39632_, \oc8051_golden_model_1.TH1 [2]);
  and (_28694_, _28692_, _39026_);
  and (_41761_, _28694_, _28691_);
  not (_28695_, \oc8051_golden_model_1.TH1 [3]);
  nor (_28696_, _03871_, _28695_);
  nor (_28697_, _11510_, _09793_);
  nor (_28698_, _28697_, _28696_);
  nor (_28699_, _28698_, _04958_);
  nor (_28700_, _28696_, _04153_);
  not (_28701_, _28700_);
  and (_28702_, _03871_, _04719_);
  nor (_28704_, _28702_, _28696_);
  nor (_28705_, _28704_, _02208_);
  and (_28706_, _28705_, _28701_);
  and (_28707_, _11511_, _03871_);
  nor (_28708_, _28707_, _28696_);
  nor (_28709_, _28708_, _03061_);
  and (_28710_, _03871_, \oc8051_golden_model_1.ACC [3]);
  nor (_28711_, _28710_, _28696_);
  nor (_28712_, _28711_, _02549_);
  nor (_28713_, _28711_, _02063_);
  nor (_28715_, _02062_, _28695_);
  or (_28716_, _28715_, _28713_);
  and (_28717_, _28716_, _03006_);
  nor (_28718_, _11394_, _09793_);
  nor (_28719_, _28718_, _28696_);
  nor (_28720_, _28719_, _03006_);
  or (_28721_, _28720_, _28717_);
  and (_28722_, _28721_, _02519_);
  nor (_28723_, _09793_, _03434_);
  nor (_28724_, _28723_, _28696_);
  nor (_28726_, _28724_, _02519_);
  nor (_28727_, _28726_, _28722_);
  nor (_28728_, _28727_, _02153_);
  or (_28729_, _28728_, _06188_);
  nor (_28730_, _28729_, _28712_);
  and (_28731_, _28724_, _06188_);
  nor (_28732_, _28731_, _28730_);
  nor (_28733_, _28732_, _02031_);
  and (_28734_, _05166_, _03871_);
  nor (_28735_, _28696_, _02032_);
  not (_28737_, _28735_);
  nor (_28738_, _28737_, _28734_);
  nor (_28739_, _28738_, _01765_);
  not (_28740_, _28739_);
  nor (_28741_, _28740_, _28733_);
  nor (_28742_, _11490_, _09793_);
  nor (_28743_, _28742_, _28696_);
  nor (_28744_, _28743_, _02037_);
  or (_28745_, _28744_, _07629_);
  or (_28746_, _28745_, _28741_);
  and (_28748_, _11505_, _03871_);
  or (_28749_, _28696_, _03059_);
  or (_28750_, _28749_, _28748_);
  and (_28751_, _28704_, _01994_);
  nor (_28752_, _28751_, _02331_);
  and (_28753_, _28752_, _28750_);
  and (_28754_, _28753_, _28746_);
  nor (_28755_, _28754_, _28709_);
  nor (_28756_, _28755_, _02206_);
  nor (_28757_, _28756_, _28706_);
  nor (_28759_, _28757_, _02342_);
  or (_28760_, _28700_, _03065_);
  nor (_28761_, _28760_, _28711_);
  or (_28762_, _28761_, _02202_);
  nor (_28763_, _28762_, _28759_);
  nor (_28764_, _11503_, _09793_);
  or (_28765_, _28696_, _04953_);
  nor (_28766_, _28765_, _28764_);
  or (_28767_, _28766_, _02334_);
  nor (_28768_, _28767_, _28763_);
  nor (_28770_, _28768_, _28699_);
  nor (_28771_, _28770_, _02366_);
  nor (_28772_, _28719_, _02778_);
  or (_28773_, _28772_, _02081_);
  nor (_28774_, _28773_, _28771_);
  and (_28775_, _11567_, _03871_);
  nor (_28776_, _28775_, _28696_);
  and (_28777_, _28776_, _02081_);
  nor (_28778_, _28777_, _28774_);
  or (_28779_, _28778_, _39633_);
  or (_28781_, _39632_, \oc8051_golden_model_1.TH1 [3]);
  and (_28782_, _28781_, _39026_);
  and (_41762_, _28782_, _28779_);
  not (_28783_, \oc8051_golden_model_1.TH1 [4]);
  nor (_28784_, _03871_, _28783_);
  nor (_28785_, _11587_, _09793_);
  nor (_28786_, _28785_, _28784_);
  nor (_28787_, _28786_, _04958_);
  and (_28788_, _11588_, _03871_);
  nor (_28789_, _28788_, _28784_);
  nor (_28791_, _28789_, _03061_);
  and (_28792_, _05303_, _03871_);
  or (_28793_, _28792_, _28784_);
  and (_28794_, _28793_, _02031_);
  and (_28795_, _03871_, \oc8051_golden_model_1.ACC [4]);
  nor (_28796_, _28795_, _28784_);
  nor (_28797_, _28796_, _02063_);
  nor (_28798_, _02062_, _28783_);
  or (_28799_, _28798_, _28797_);
  and (_28800_, _28799_, _03006_);
  nor (_28802_, _11611_, _09793_);
  nor (_28803_, _28802_, _28784_);
  nor (_28804_, _28803_, _03006_);
  or (_28805_, _28804_, _28800_);
  and (_28806_, _28805_, _02519_);
  nor (_28807_, _04372_, _09793_);
  nor (_28808_, _28807_, _28784_);
  nor (_28809_, _28808_, _02519_);
  nor (_28810_, _28809_, _28806_);
  nor (_28811_, _28810_, _02153_);
  nor (_28813_, _28796_, _02549_);
  nor (_28814_, _28813_, _06188_);
  not (_28815_, _28814_);
  nor (_28816_, _28815_, _28811_);
  and (_28817_, _28808_, _06188_);
  or (_28818_, _28817_, _02031_);
  nor (_28819_, _28818_, _28816_);
  or (_28820_, _28819_, _28794_);
  and (_28821_, _28820_, _02037_);
  nor (_28822_, _11704_, _09793_);
  nor (_28823_, _28822_, _28784_);
  nor (_28824_, _28823_, _02037_);
  or (_28825_, _28824_, _07629_);
  or (_28826_, _28825_, _28821_);
  and (_28827_, _11592_, _03871_);
  or (_28828_, _28784_, _03059_);
  or (_28829_, _28828_, _28827_);
  and (_28830_, _04831_, _03871_);
  nor (_28831_, _28830_, _28784_);
  and (_28832_, _28831_, _01994_);
  nor (_28834_, _28832_, _02331_);
  and (_28835_, _28834_, _28829_);
  and (_28836_, _28835_, _28826_);
  nor (_28837_, _28836_, _28791_);
  nor (_28838_, _28837_, _02206_);
  nor (_28839_, _28784_, _04420_);
  not (_28840_, _28839_);
  nor (_28841_, _28831_, _02208_);
  and (_28842_, _28841_, _28840_);
  nor (_28843_, _28842_, _28838_);
  nor (_28845_, _28843_, _02342_);
  or (_28846_, _28839_, _03065_);
  nor (_28847_, _28846_, _28796_);
  or (_28848_, _28847_, _02202_);
  nor (_28849_, _28848_, _28845_);
  nor (_28850_, _11590_, _09793_);
  or (_28851_, _28784_, _04953_);
  nor (_28852_, _28851_, _28850_);
  or (_28853_, _28852_, _02334_);
  nor (_28854_, _28853_, _28849_);
  nor (_28856_, _28854_, _28787_);
  nor (_28857_, _28856_, _02366_);
  nor (_28858_, _28803_, _02778_);
  or (_28859_, _28858_, _02081_);
  nor (_28860_, _28859_, _28857_);
  and (_28861_, _11771_, _03871_);
  nor (_28862_, _28861_, _28784_);
  and (_28863_, _28862_, _02081_);
  nor (_28864_, _28863_, _28860_);
  or (_28865_, _28864_, _39633_);
  or (_28867_, _39632_, \oc8051_golden_model_1.TH1 [4]);
  and (_28868_, _28867_, _39026_);
  and (_41763_, _28868_, _28865_);
  not (_28869_, \oc8051_golden_model_1.TH1 [5]);
  nor (_28870_, _03871_, _28869_);
  nor (_28871_, _11785_, _09793_);
  nor (_28872_, _28871_, _28870_);
  nor (_28873_, _28872_, _04958_);
  and (_28874_, _11786_, _03871_);
  nor (_28875_, _28874_, _28870_);
  nor (_28877_, _28875_, _03061_);
  and (_28878_, _04827_, _03871_);
  nor (_28879_, _28878_, _28870_);
  and (_28880_, _28879_, _01994_);
  and (_28881_, _03871_, \oc8051_golden_model_1.ACC [5]);
  nor (_28882_, _28881_, _28870_);
  nor (_28883_, _28882_, _02549_);
  nor (_28884_, _28882_, _02063_);
  nor (_28885_, _02062_, _28869_);
  or (_28886_, _28885_, _28884_);
  and (_28888_, _28886_, _03006_);
  nor (_28889_, _11804_, _09793_);
  nor (_28890_, _28889_, _28870_);
  nor (_28891_, _28890_, _03006_);
  or (_28892_, _28891_, _28888_);
  and (_28893_, _28892_, _02519_);
  nor (_28894_, _04057_, _09793_);
  nor (_28895_, _28894_, _28870_);
  nor (_28896_, _28895_, _02519_);
  nor (_28897_, _28896_, _28893_);
  nor (_28899_, _28897_, _02153_);
  or (_28900_, _28899_, _06188_);
  nor (_28901_, _28900_, _28883_);
  and (_28902_, _28895_, _06188_);
  nor (_28903_, _28902_, _28901_);
  nor (_28904_, _28903_, _02031_);
  and (_28905_, _05258_, _03871_);
  nor (_28906_, _28870_, _02032_);
  not (_28907_, _28906_);
  nor (_28908_, _28907_, _28905_);
  or (_28910_, _28908_, _01765_);
  nor (_28911_, _28910_, _28904_);
  nor (_28912_, _11900_, _09793_);
  nor (_28913_, _28912_, _28870_);
  nor (_28914_, _28913_, _02037_);
  or (_28915_, _28914_, _01994_);
  nor (_28916_, _28915_, _28911_);
  nor (_28917_, _28916_, _28880_);
  or (_28918_, _28917_, _02210_);
  and (_28919_, _11915_, _03871_);
  or (_28921_, _28919_, _28870_);
  or (_28922_, _28921_, _03059_);
  and (_28923_, _28922_, _03061_);
  and (_28924_, _28923_, _28918_);
  nor (_28925_, _28924_, _28877_);
  nor (_28926_, _28925_, _02206_);
  nor (_28927_, _28870_, _04104_);
  not (_28928_, _28927_);
  nor (_28929_, _28879_, _02208_);
  and (_28930_, _28929_, _28928_);
  nor (_28932_, _28930_, _28926_);
  nor (_28933_, _28932_, _02342_);
  or (_28934_, _28927_, _03065_);
  nor (_28935_, _28934_, _28882_);
  or (_28936_, _28935_, _02202_);
  nor (_28937_, _28936_, _28933_);
  nor (_28938_, _11913_, _09793_);
  or (_28939_, _28870_, _04953_);
  nor (_28940_, _28939_, _28938_);
  or (_28941_, _28940_, _02334_);
  nor (_28943_, _28941_, _28937_);
  nor (_28944_, _28943_, _28873_);
  nor (_28945_, _28944_, _02366_);
  nor (_28946_, _28890_, _02778_);
  or (_28947_, _28946_, _02081_);
  nor (_28948_, _28947_, _28945_);
  and (_28949_, _11974_, _03871_);
  nor (_28950_, _28949_, _28870_);
  and (_28951_, _28950_, _02081_);
  nor (_28952_, _28951_, _28948_);
  or (_28954_, _28952_, _39633_);
  or (_28955_, _39632_, \oc8051_golden_model_1.TH1 [5]);
  and (_28956_, _28955_, _39026_);
  and (_41764_, _28956_, _28954_);
  not (_28957_, \oc8051_golden_model_1.TH1 [6]);
  nor (_28958_, _03871_, _28957_);
  nor (_28959_, _12117_, _09793_);
  nor (_28960_, _28959_, _28958_);
  nor (_28961_, _28960_, _04958_);
  and (_28962_, _12118_, _03871_);
  nor (_28964_, _28962_, _28958_);
  nor (_28965_, _28964_, _03061_);
  and (_28966_, _12103_, _03871_);
  nor (_28967_, _28966_, _28958_);
  and (_28968_, _28967_, _01994_);
  and (_28969_, _03871_, \oc8051_golden_model_1.ACC [6]);
  nor (_28970_, _28969_, _28958_);
  nor (_28971_, _28970_, _02549_);
  nor (_28972_, _28970_, _02063_);
  nor (_28973_, _02062_, _28957_);
  or (_28974_, _28973_, _28972_);
  and (_28975_, _28974_, _03006_);
  nor (_28976_, _11993_, _09793_);
  nor (_28977_, _28976_, _28958_);
  nor (_28978_, _28977_, _03006_);
  or (_28979_, _28978_, _28975_);
  and (_28980_, _28979_, _02519_);
  nor (_28981_, _03964_, _09793_);
  nor (_28982_, _28981_, _28958_);
  nor (_28983_, _28982_, _02519_);
  nor (_28985_, _28983_, _28980_);
  nor (_28986_, _28985_, _02153_);
  or (_28987_, _28986_, _06188_);
  nor (_28988_, _28987_, _28971_);
  and (_28989_, _28982_, _06188_);
  nor (_28990_, _28989_, _28988_);
  nor (_28991_, _28990_, _02031_);
  and (_28992_, _05029_, _03871_);
  nor (_28993_, _28958_, _02032_);
  not (_28994_, _28993_);
  nor (_28996_, _28994_, _28992_);
  or (_28997_, _28996_, _01765_);
  nor (_28998_, _28997_, _28991_);
  nor (_28999_, _12096_, _09793_);
  nor (_29000_, _28999_, _28958_);
  nor (_29001_, _29000_, _02037_);
  or (_29002_, _29001_, _01994_);
  nor (_29003_, _29002_, _28998_);
  nor (_29004_, _29003_, _28968_);
  or (_29005_, _29004_, _02210_);
  and (_29007_, _12112_, _03871_);
  or (_29008_, _29007_, _28958_);
  or (_29009_, _29008_, _03059_);
  and (_29010_, _29009_, _03061_);
  and (_29011_, _29010_, _29005_);
  nor (_29012_, _29011_, _28965_);
  nor (_29013_, _29012_, _02206_);
  nor (_29014_, _28958_, _04011_);
  not (_29015_, _29014_);
  nor (_29016_, _28967_, _02208_);
  and (_29018_, _29016_, _29015_);
  nor (_29019_, _29018_, _29013_);
  nor (_29020_, _29019_, _02342_);
  or (_29021_, _29014_, _03065_);
  nor (_29022_, _29021_, _28970_);
  or (_29023_, _29022_, _02202_);
  nor (_29024_, _29023_, _29020_);
  nor (_29025_, _12110_, _09793_);
  or (_29026_, _28958_, _04953_);
  nor (_29027_, _29026_, _29025_);
  or (_29029_, _29027_, _02334_);
  nor (_29030_, _29029_, _29024_);
  nor (_29031_, _29030_, _28961_);
  nor (_29032_, _29031_, _02366_);
  nor (_29033_, _28977_, _02778_);
  or (_29034_, _29033_, _02081_);
  nor (_29035_, _29034_, _29032_);
  and (_29036_, _12178_, _03871_);
  nor (_29037_, _29036_, _28958_);
  and (_29038_, _29037_, _02081_);
  nor (_29040_, _29038_, _29035_);
  or (_29041_, _29040_, _39633_);
  or (_29042_, _39632_, \oc8051_golden_model_1.TH1 [6]);
  and (_29043_, _29042_, _39026_);
  and (_41765_, _29043_, _29041_);
  not (_29044_, \oc8051_golden_model_1.TL0 [0]);
  nor (_29045_, _03876_, _29044_);
  nor (_29046_, _04257_, _09872_);
  nor (_29047_, _29046_, _29045_);
  and (_29048_, _29047_, _15890_);
  and (_29050_, _03876_, \oc8051_golden_model_1.ACC [0]);
  nor (_29051_, _29050_, _29045_);
  nor (_29052_, _29051_, _02549_);
  nor (_29053_, _29051_, _02063_);
  nor (_29054_, _02062_, _29044_);
  or (_29055_, _29054_, _29053_);
  and (_29056_, _29055_, _03006_);
  nor (_29057_, _29047_, _03006_);
  or (_29058_, _29057_, _29056_);
  and (_29059_, _29058_, _02519_);
  and (_29061_, _03876_, _03002_);
  nor (_29062_, _29061_, _29045_);
  nor (_29063_, _29062_, _02519_);
  nor (_29064_, _29063_, _29059_);
  nor (_29065_, _29064_, _02153_);
  or (_29066_, _29065_, _06188_);
  nor (_29067_, _29066_, _29052_);
  and (_29068_, _29062_, _06188_);
  nor (_29069_, _29068_, _29067_);
  nor (_29070_, _29069_, _02031_);
  and (_29073_, _05120_, _03876_);
  nor (_29074_, _29045_, _02032_);
  not (_29075_, _29074_);
  nor (_29076_, _29075_, _29073_);
  nor (_29077_, _29076_, _29070_);
  nor (_29078_, _29077_, _01765_);
  nor (_29079_, _10898_, _09872_);
  or (_29080_, _29045_, _02037_);
  nor (_29081_, _29080_, _29079_);
  or (_29082_, _29081_, _01994_);
  nor (_29084_, _29082_, _29078_);
  and (_29085_, _03876_, _04837_);
  nor (_29086_, _29085_, _29045_);
  nor (_29087_, _29086_, _01995_);
  or (_29088_, _29087_, _29084_);
  and (_29089_, _29088_, _03059_);
  and (_29090_, _10914_, _03876_);
  nor (_29091_, _29090_, _29045_);
  nor (_29092_, _29091_, _03059_);
  or (_29093_, _29092_, _29089_);
  and (_29095_, _29093_, _03061_);
  and (_29096_, _10792_, _03876_);
  nor (_29097_, _29096_, _29045_);
  nor (_29098_, _29097_, _03061_);
  or (_29099_, _29098_, _29095_);
  and (_29100_, _29099_, _02208_);
  or (_29101_, _29086_, _02208_);
  nor (_29102_, _29101_, _29046_);
  nor (_29103_, _29102_, _29100_);
  nor (_29104_, _29103_, _02342_);
  and (_29106_, _10791_, _03876_);
  or (_29107_, _29106_, _29045_);
  and (_29108_, _29107_, _02342_);
  or (_29109_, _29108_, _29104_);
  and (_29110_, _29109_, _04953_);
  nor (_29111_, _10913_, _09872_);
  nor (_29112_, _29111_, _29045_);
  nor (_29113_, _29112_, _04953_);
  or (_29114_, _29113_, _29110_);
  and (_29115_, _29114_, _04958_);
  nor (_29117_, _10789_, _09872_);
  nor (_29118_, _29117_, _29045_);
  nor (_29119_, _29118_, _04958_);
  nor (_29120_, _29119_, _15890_);
  not (_29121_, _29120_);
  nor (_29122_, _29121_, _29115_);
  nor (_29123_, _29122_, _29048_);
  or (_29124_, _29123_, _39633_);
  or (_29125_, _39632_, \oc8051_golden_model_1.TL0 [0]);
  and (_29126_, _29125_, _39026_);
  and (_41767_, _29126_, _29124_);
  nor (_29127_, _03876_, \oc8051_golden_model_1.TL0 [1]);
  not (_29128_, _29127_);
  nor (_29129_, _11113_, _09872_);
  nor (_29130_, _29129_, _03061_);
  and (_29131_, _29130_, _29128_);
  and (_29132_, _05075_, _03876_);
  not (_29133_, \oc8051_golden_model_1.TL0 [1]);
  nor (_29134_, _03876_, _29133_);
  nor (_29135_, _29134_, _02032_);
  not (_29137_, _29135_);
  nor (_29138_, _29137_, _29132_);
  not (_29139_, _29138_);
  and (_29140_, _03876_, _01804_);
  nor (_29141_, _29140_, _29127_);
  and (_29142_, _29141_, _02153_);
  and (_29143_, _29141_, _02062_);
  nor (_29144_, _02062_, _29133_);
  or (_29145_, _29144_, _29143_);
  and (_29146_, _29145_, _03006_);
  and (_29148_, _11001_, _03876_);
  nor (_29149_, _29148_, _29127_);
  and (_29150_, _29149_, _02158_);
  or (_29151_, _29150_, _29146_);
  and (_29152_, _29151_, _02519_);
  nor (_29153_, _09872_, _03161_);
  nor (_29154_, _29153_, _29134_);
  nor (_29155_, _29154_, _02519_);
  nor (_29156_, _29155_, _29152_);
  nor (_29157_, _29156_, _02153_);
  or (_29159_, _29157_, _06188_);
  nor (_29160_, _29159_, _29142_);
  and (_29161_, _29154_, _06188_);
  nor (_29162_, _29161_, _29160_);
  nor (_29163_, _29162_, _02031_);
  nor (_29164_, _29163_, _01765_);
  and (_29165_, _29164_, _29139_);
  and (_29166_, _11096_, _03876_);
  nor (_29167_, _29166_, _02037_);
  and (_29168_, _29167_, _29128_);
  nor (_29170_, _29168_, _29165_);
  nor (_29171_, _29170_, _07629_);
  nor (_29172_, _10989_, _09872_);
  nor (_29173_, _29172_, _03059_);
  and (_29174_, _03876_, _02893_);
  nor (_29175_, _29174_, _01995_);
  nor (_29176_, _29175_, _29173_);
  nor (_29177_, _29176_, _29127_);
  nor (_29178_, _29177_, _29171_);
  nor (_29179_, _29178_, _02331_);
  nor (_29182_, _29179_, _29131_);
  nor (_29183_, _29182_, _02206_);
  nor (_29184_, _10988_, _09872_);
  nor (_29185_, _29184_, _02208_);
  and (_29186_, _29185_, _29128_);
  nor (_29187_, _29186_, _29183_);
  nor (_29188_, _29187_, _02342_);
  nor (_29189_, _29134_, _04209_);
  nor (_29190_, _29189_, _03065_);
  and (_29191_, _29190_, _29141_);
  nor (_29193_, _29191_, _29188_);
  or (_29194_, _29193_, _17216_);
  nand (_29195_, _29140_, _04208_);
  nor (_29196_, _29127_, _04958_);
  and (_29197_, _29196_, _29195_);
  nor (_29198_, _29197_, _02366_);
  and (_29199_, _29174_, _04208_);
  or (_29200_, _29127_, _04953_);
  or (_29201_, _29200_, _29199_);
  and (_29202_, _29201_, _29198_);
  and (_29204_, _29202_, _29194_);
  nor (_29205_, _29149_, _02778_);
  nor (_29206_, _29205_, _29204_);
  nor (_29207_, _29206_, _02081_);
  nor (_29208_, _29148_, _29134_);
  and (_29209_, _29208_, _02081_);
  nor (_29210_, _29209_, _29207_);
  or (_29211_, _29210_, _39633_);
  or (_29212_, _39632_, \oc8051_golden_model_1.TL0 [1]);
  and (_29213_, _29212_, _39026_);
  and (_41768_, _29213_, _29211_);
  not (_29215_, \oc8051_golden_model_1.TL0 [2]);
  nor (_29216_, _03876_, _29215_);
  nor (_29217_, _11314_, _09872_);
  nor (_29218_, _29217_, _29216_);
  nor (_29219_, _29218_, _04958_);
  and (_29220_, _11315_, _03876_);
  nor (_29221_, _29220_, _29216_);
  nor (_29222_, _29221_, _03061_);
  and (_29223_, _03876_, _04866_);
  nor (_29225_, _29223_, _29216_);
  and (_29226_, _29225_, _01994_);
  and (_29227_, _03876_, \oc8051_golden_model_1.ACC [2]);
  nor (_29228_, _29227_, _29216_);
  nor (_29229_, _29228_, _02549_);
  nor (_29230_, _29228_, _02063_);
  nor (_29231_, _02062_, _29215_);
  or (_29232_, _29231_, _29230_);
  and (_29233_, _29232_, _03006_);
  nor (_29234_, _11199_, _09872_);
  nor (_29236_, _29234_, _29216_);
  nor (_29237_, _29236_, _03006_);
  or (_29238_, _29237_, _29233_);
  and (_29239_, _29238_, _02519_);
  nor (_29240_, _09872_, _03624_);
  nor (_29241_, _29240_, _29216_);
  nor (_29242_, _29241_, _02519_);
  nor (_29243_, _29242_, _29239_);
  nor (_29244_, _29243_, _02153_);
  or (_29245_, _29244_, _06188_);
  nor (_29246_, _29245_, _29229_);
  and (_29247_, _29241_, _06188_);
  nor (_29248_, _29247_, _29246_);
  nor (_29249_, _29248_, _02031_);
  and (_29250_, _05211_, _03876_);
  nor (_29251_, _29216_, _02032_);
  not (_29252_, _29251_);
  nor (_29253_, _29252_, _29250_);
  or (_29254_, _29253_, _01765_);
  nor (_29255_, _29254_, _29249_);
  nor (_29257_, _11298_, _09872_);
  nor (_29258_, _29257_, _29216_);
  nor (_29259_, _29258_, _02037_);
  or (_29260_, _29259_, _01994_);
  nor (_29261_, _29260_, _29255_);
  nor (_29262_, _29261_, _29226_);
  or (_29263_, _29262_, _02210_);
  and (_29264_, _11189_, _03876_);
  or (_29265_, _29264_, _29216_);
  or (_29266_, _29265_, _03059_);
  and (_29268_, _29266_, _03061_);
  and (_29269_, _29268_, _29263_);
  nor (_29270_, _29269_, _29222_);
  nor (_29271_, _29270_, _02206_);
  nor (_29272_, _29216_, _04309_);
  not (_29273_, _29272_);
  nor (_29274_, _29225_, _02208_);
  and (_29275_, _29274_, _29273_);
  nor (_29276_, _29275_, _29271_);
  nor (_29277_, _29276_, _02342_);
  or (_29279_, _29272_, _03065_);
  nor (_29280_, _29279_, _29228_);
  or (_29281_, _29280_, _02202_);
  nor (_29282_, _29281_, _29277_);
  nor (_29283_, _11187_, _09872_);
  or (_29284_, _29216_, _04953_);
  nor (_29285_, _29284_, _29283_);
  or (_29286_, _29285_, _02334_);
  nor (_29287_, _29286_, _29282_);
  nor (_29288_, _29287_, _29219_);
  nor (_29291_, _29288_, _02366_);
  nor (_29292_, _29236_, _02778_);
  or (_29293_, _29292_, _02081_);
  nor (_29294_, _29293_, _29291_);
  and (_29295_, _11367_, _03876_);
  nor (_29296_, _29295_, _29216_);
  and (_29297_, _29296_, _02081_);
  nor (_29298_, _29297_, _29294_);
  or (_29299_, _29298_, _39633_);
  or (_29300_, _39632_, \oc8051_golden_model_1.TL0 [2]);
  and (_29302_, _29300_, _39026_);
  and (_41769_, _29302_, _29299_);
  not (_29303_, \oc8051_golden_model_1.TL0 [3]);
  nor (_29304_, _03876_, _29303_);
  nor (_29305_, _11510_, _09872_);
  nor (_29306_, _29305_, _29304_);
  nor (_29307_, _29306_, _04958_);
  nor (_29308_, _29304_, _04153_);
  not (_29309_, _29308_);
  and (_29310_, _03876_, _04719_);
  nor (_29312_, _29310_, _29304_);
  nor (_29313_, _29312_, _02208_);
  and (_29314_, _29313_, _29309_);
  and (_29315_, _11511_, _03876_);
  nor (_29316_, _29315_, _29304_);
  nor (_29317_, _29316_, _03061_);
  nor (_29318_, _09872_, _03434_);
  nor (_29319_, _29318_, _29304_);
  and (_29320_, _29319_, _06188_);
  and (_29321_, _03876_, \oc8051_golden_model_1.ACC [3]);
  nor (_29323_, _29321_, _29304_);
  nor (_29324_, _29323_, _02063_);
  nor (_29325_, _02062_, _29303_);
  or (_29326_, _29325_, _29324_);
  and (_29327_, _29326_, _03006_);
  nor (_29328_, _11394_, _09872_);
  nor (_29329_, _29328_, _29304_);
  nor (_29330_, _29329_, _03006_);
  or (_29331_, _29330_, _29327_);
  and (_29332_, _29331_, _02519_);
  nor (_29334_, _29319_, _02519_);
  nor (_29335_, _29334_, _29332_);
  nor (_29336_, _29335_, _02153_);
  nor (_29337_, _29323_, _02549_);
  nor (_29338_, _29337_, _06188_);
  not (_29339_, _29338_);
  nor (_29340_, _29339_, _29336_);
  nor (_29341_, _29340_, _29320_);
  nor (_29342_, _29341_, _02031_);
  and (_29343_, _05166_, _03876_);
  nor (_29345_, _29304_, _02032_);
  not (_29346_, _29345_);
  nor (_29347_, _29346_, _29343_);
  nor (_29348_, _29347_, _01765_);
  not (_29349_, _29348_);
  nor (_29350_, _29349_, _29342_);
  nor (_29351_, _11490_, _09872_);
  nor (_29352_, _29351_, _29304_);
  nor (_29353_, _29352_, _02037_);
  or (_29354_, _29353_, _07629_);
  or (_29356_, _29354_, _29350_);
  and (_29357_, _11505_, _03876_);
  or (_29358_, _29304_, _03059_);
  or (_29359_, _29358_, _29357_);
  and (_29360_, _29312_, _01994_);
  nor (_29361_, _29360_, _02331_);
  and (_29362_, _29361_, _29359_);
  and (_29363_, _29362_, _29356_);
  nor (_29364_, _29363_, _29317_);
  nor (_29365_, _29364_, _02206_);
  nor (_29367_, _29365_, _29314_);
  nor (_29368_, _29367_, _02342_);
  or (_29369_, _29308_, _03065_);
  nor (_29370_, _29369_, _29323_);
  or (_29371_, _29370_, _02202_);
  nor (_29372_, _29371_, _29368_);
  nor (_29373_, _11503_, _09872_);
  or (_29374_, _29304_, _04953_);
  nor (_29375_, _29374_, _29373_);
  or (_29376_, _29375_, _02334_);
  nor (_29378_, _29376_, _29372_);
  nor (_29379_, _29378_, _29307_);
  nor (_29380_, _29379_, _02366_);
  nor (_29381_, _29329_, _02778_);
  or (_29382_, _29381_, _02081_);
  nor (_29383_, _29382_, _29380_);
  and (_29384_, _11567_, _03876_);
  nor (_29385_, _29384_, _29304_);
  and (_29386_, _29385_, _02081_);
  nor (_29387_, _29386_, _29383_);
  or (_29389_, _29387_, _39633_);
  or (_29390_, _39632_, \oc8051_golden_model_1.TL0 [3]);
  and (_29391_, _29390_, _39026_);
  and (_41770_, _29391_, _29389_);
  not (_29392_, \oc8051_golden_model_1.TL0 [4]);
  nor (_29393_, _03876_, _29392_);
  nor (_29394_, _11587_, _09872_);
  nor (_29395_, _29394_, _29393_);
  nor (_29396_, _29395_, _04958_);
  nor (_29397_, _29393_, _04420_);
  not (_29399_, _29397_);
  and (_29400_, _04831_, _03876_);
  nor (_29401_, _29400_, _29393_);
  nor (_29402_, _29401_, _02208_);
  and (_29403_, _29402_, _29399_);
  and (_29404_, _11588_, _03876_);
  nor (_29405_, _29404_, _29393_);
  nor (_29406_, _29405_, _03061_);
  and (_29407_, _05303_, _03876_);
  or (_29408_, _29407_, _29393_);
  and (_29410_, _29408_, _02031_);
  and (_29411_, _03876_, \oc8051_golden_model_1.ACC [4]);
  nor (_29412_, _29411_, _29393_);
  nor (_29413_, _29412_, _02549_);
  nor (_29414_, _29412_, _02063_);
  nor (_29415_, _02062_, _29392_);
  or (_29416_, _29415_, _29414_);
  and (_29417_, _29416_, _03006_);
  nor (_29418_, _11611_, _09872_);
  nor (_29419_, _29418_, _29393_);
  nor (_29421_, _29419_, _03006_);
  or (_29422_, _29421_, _29417_);
  and (_29423_, _29422_, _02519_);
  nor (_29424_, _04372_, _09872_);
  nor (_29425_, _29424_, _29393_);
  nor (_29426_, _29425_, _02519_);
  nor (_29427_, _29426_, _29423_);
  nor (_29428_, _29427_, _02153_);
  or (_29429_, _29428_, _06188_);
  nor (_29430_, _29429_, _29413_);
  and (_29432_, _29425_, _06188_);
  or (_29433_, _29432_, _02031_);
  nor (_29434_, _29433_, _29430_);
  or (_29435_, _29434_, _29410_);
  and (_29436_, _29435_, _02037_);
  nor (_29437_, _11704_, _09872_);
  nor (_29438_, _29437_, _29393_);
  nor (_29439_, _29438_, _02037_);
  or (_29440_, _29439_, _07629_);
  or (_29441_, _29440_, _29436_);
  and (_29443_, _11592_, _03876_);
  or (_29444_, _29393_, _03059_);
  or (_29445_, _29444_, _29443_);
  and (_29446_, _29401_, _01994_);
  nor (_29447_, _29446_, _02331_);
  and (_29448_, _29447_, _29445_);
  and (_29449_, _29448_, _29441_);
  nor (_29450_, _29449_, _29406_);
  nor (_29451_, _29450_, _02206_);
  nor (_29452_, _29451_, _29403_);
  nor (_29454_, _29452_, _02342_);
  or (_29455_, _29397_, _03065_);
  nor (_29456_, _29455_, _29412_);
  or (_29457_, _29456_, _02202_);
  nor (_29458_, _29457_, _29454_);
  nor (_29459_, _11590_, _09872_);
  or (_29460_, _29393_, _04953_);
  nor (_29461_, _29460_, _29459_);
  or (_29462_, _29461_, _02334_);
  nor (_29463_, _29462_, _29458_);
  nor (_29465_, _29463_, _29396_);
  nor (_29466_, _29465_, _02366_);
  nor (_29467_, _29419_, _02778_);
  or (_29468_, _29467_, _02081_);
  nor (_29469_, _29468_, _29466_);
  and (_29470_, _11771_, _03876_);
  nor (_29471_, _29470_, _29393_);
  and (_29472_, _29471_, _02081_);
  nor (_29473_, _29472_, _29469_);
  or (_29474_, _29473_, _39633_);
  or (_29476_, _39632_, \oc8051_golden_model_1.TL0 [4]);
  and (_29477_, _29476_, _39026_);
  and (_41771_, _29477_, _29474_);
  not (_29478_, \oc8051_golden_model_1.TL0 [5]);
  nor (_29479_, _03876_, _29478_);
  nor (_29480_, _11785_, _09872_);
  nor (_29481_, _29480_, _29479_);
  nor (_29482_, _29481_, _04958_);
  and (_29483_, _11786_, _03876_);
  nor (_29484_, _29483_, _29479_);
  nor (_29486_, _29484_, _03061_);
  and (_29487_, _04827_, _03876_);
  nor (_29488_, _29487_, _29479_);
  and (_29489_, _29488_, _01994_);
  nor (_29490_, _04057_, _09872_);
  nor (_29491_, _29490_, _29479_);
  and (_29492_, _29491_, _06188_);
  and (_29493_, _03876_, \oc8051_golden_model_1.ACC [5]);
  nor (_29494_, _29493_, _29479_);
  nor (_29495_, _29494_, _02063_);
  nor (_29497_, _02062_, _29478_);
  or (_29498_, _29497_, _29495_);
  and (_29499_, _29498_, _03006_);
  nor (_29500_, _11804_, _09872_);
  nor (_29501_, _29500_, _29479_);
  nor (_29502_, _29501_, _03006_);
  or (_29503_, _29502_, _29499_);
  and (_29504_, _29503_, _02519_);
  nor (_29505_, _29491_, _02519_);
  nor (_29506_, _29505_, _29504_);
  nor (_29509_, _29506_, _02153_);
  nor (_29510_, _29494_, _02549_);
  nor (_29511_, _29510_, _06188_);
  not (_29512_, _29511_);
  nor (_29513_, _29512_, _29509_);
  nor (_29514_, _29513_, _29492_);
  nor (_29515_, _29514_, _02031_);
  and (_29516_, _05258_, _03876_);
  nor (_29517_, _29479_, _02032_);
  not (_29518_, _29517_);
  nor (_29520_, _29518_, _29516_);
  or (_29521_, _29520_, _01765_);
  nor (_29522_, _29521_, _29515_);
  nor (_29523_, _11900_, _09872_);
  nor (_29524_, _29523_, _29479_);
  nor (_29525_, _29524_, _02037_);
  or (_29526_, _29525_, _01994_);
  nor (_29527_, _29526_, _29522_);
  nor (_29528_, _29527_, _29489_);
  or (_29529_, _29528_, _02210_);
  and (_29531_, _11915_, _03876_);
  or (_29532_, _29531_, _29479_);
  or (_29533_, _29532_, _03059_);
  and (_29534_, _29533_, _03061_);
  and (_29535_, _29534_, _29529_);
  nor (_29536_, _29535_, _29486_);
  nor (_29537_, _29536_, _02206_);
  nor (_29538_, _29479_, _04104_);
  not (_29539_, _29538_);
  nor (_29540_, _29488_, _02208_);
  and (_29542_, _29540_, _29539_);
  nor (_29543_, _29542_, _29537_);
  nor (_29544_, _29543_, _02342_);
  or (_29545_, _29538_, _03065_);
  nor (_29546_, _29545_, _29494_);
  or (_29547_, _29546_, _02202_);
  nor (_29548_, _29547_, _29544_);
  nor (_29549_, _11913_, _09872_);
  or (_29550_, _29479_, _04953_);
  nor (_29551_, _29550_, _29549_);
  or (_29552_, _29551_, _02334_);
  nor (_29553_, _29552_, _29548_);
  nor (_29554_, _29553_, _29482_);
  nor (_29555_, _29554_, _02366_);
  nor (_29556_, _29501_, _02778_);
  or (_29557_, _29556_, _02081_);
  nor (_29558_, _29557_, _29555_);
  and (_29559_, _11974_, _03876_);
  nor (_29560_, _29559_, _29479_);
  and (_29561_, _29560_, _02081_);
  nor (_29563_, _29561_, _29558_);
  or (_29564_, _29563_, _39633_);
  or (_29565_, _39632_, \oc8051_golden_model_1.TL0 [5]);
  and (_29566_, _29565_, _39026_);
  and (_41772_, _29566_, _29564_);
  not (_29567_, \oc8051_golden_model_1.TL0 [6]);
  nor (_29568_, _03876_, _29567_);
  nor (_29569_, _12117_, _09872_);
  nor (_29570_, _29569_, _29568_);
  nor (_29571_, _29570_, _04958_);
  and (_29573_, _12118_, _03876_);
  nor (_29574_, _29573_, _29568_);
  nor (_29575_, _29574_, _03061_);
  and (_29576_, _12103_, _03876_);
  nor (_29577_, _29576_, _29568_);
  and (_29578_, _29577_, _01994_);
  and (_29579_, _03876_, \oc8051_golden_model_1.ACC [6]);
  nor (_29580_, _29579_, _29568_);
  nor (_29581_, _29580_, _02549_);
  nor (_29582_, _29580_, _02063_);
  nor (_29584_, _02062_, _29567_);
  or (_29585_, _29584_, _29582_);
  and (_29586_, _29585_, _03006_);
  nor (_29587_, _11993_, _09872_);
  nor (_29588_, _29587_, _29568_);
  nor (_29589_, _29588_, _03006_);
  or (_29590_, _29589_, _29586_);
  and (_29591_, _29590_, _02519_);
  nor (_29592_, _03964_, _09872_);
  nor (_29593_, _29592_, _29568_);
  nor (_29595_, _29593_, _02519_);
  nor (_29596_, _29595_, _29591_);
  nor (_29597_, _29596_, _02153_);
  or (_29598_, _29597_, _06188_);
  nor (_29599_, _29598_, _29581_);
  and (_29600_, _29593_, _06188_);
  nor (_29601_, _29600_, _29599_);
  nor (_29602_, _29601_, _02031_);
  and (_29603_, _05029_, _03876_);
  nor (_29604_, _29568_, _02032_);
  not (_29606_, _29604_);
  nor (_29607_, _29606_, _29603_);
  or (_29608_, _29607_, _01765_);
  nor (_29609_, _29608_, _29602_);
  nor (_29610_, _12096_, _09872_);
  nor (_29611_, _29610_, _29568_);
  nor (_29612_, _29611_, _02037_);
  or (_29613_, _29612_, _01994_);
  nor (_29614_, _29613_, _29609_);
  nor (_29615_, _29614_, _29578_);
  or (_29618_, _29615_, _02210_);
  and (_29619_, _12112_, _03876_);
  or (_29620_, _29619_, _29568_);
  or (_29621_, _29620_, _03059_);
  and (_29622_, _29621_, _03061_);
  and (_29623_, _29622_, _29618_);
  nor (_29624_, _29623_, _29575_);
  nor (_29625_, _29624_, _02206_);
  nor (_29626_, _29568_, _04011_);
  not (_29627_, _29626_);
  nor (_29629_, _29577_, _02208_);
  and (_29630_, _29629_, _29627_);
  nor (_29631_, _29630_, _29625_);
  nor (_29632_, _29631_, _02342_);
  or (_29633_, _29626_, _03065_);
  nor (_29634_, _29633_, _29580_);
  or (_29635_, _29634_, _02202_);
  nor (_29636_, _29635_, _29632_);
  nor (_29637_, _12110_, _09872_);
  or (_29638_, _29568_, _04953_);
  nor (_29640_, _29638_, _29637_);
  or (_29641_, _29640_, _02334_);
  nor (_29642_, _29641_, _29636_);
  nor (_29643_, _29642_, _29571_);
  nor (_29644_, _29643_, _02366_);
  nor (_29645_, _29588_, _02778_);
  or (_29646_, _29645_, _02081_);
  nor (_29647_, _29646_, _29644_);
  and (_29648_, _12178_, _03876_);
  nor (_29649_, _29648_, _29568_);
  and (_29651_, _29649_, _02081_);
  nor (_29652_, _29651_, _29647_);
  or (_29653_, _29652_, _39633_);
  or (_29654_, _39632_, \oc8051_golden_model_1.TL0 [6]);
  and (_29655_, _29654_, _39026_);
  and (_41773_, _29655_, _29653_);
  not (_29656_, \oc8051_golden_model_1.TL1 [0]);
  nor (_29657_, _03864_, _29656_);
  nor (_29658_, _04257_, _09951_);
  nor (_29659_, _29658_, _29657_);
  and (_29661_, _29659_, _15890_);
  and (_29662_, _03864_, _04837_);
  nor (_29663_, _29662_, _29657_);
  nor (_29664_, _29663_, _02208_);
  not (_29665_, _29664_);
  nor (_29666_, _29665_, _29658_);
  and (_29667_, _03864_, \oc8051_golden_model_1.ACC [0]);
  nor (_29668_, _29667_, _29657_);
  nor (_29669_, _29668_, _02549_);
  nor (_29670_, _29668_, _02063_);
  nor (_29672_, _02062_, _29656_);
  or (_29673_, _29672_, _29670_);
  and (_29674_, _29673_, _03006_);
  nor (_29675_, _29659_, _03006_);
  or (_29676_, _29675_, _29674_);
  and (_29677_, _29676_, _02519_);
  and (_29678_, _04197_, _03002_);
  nor (_29679_, _29678_, _29657_);
  nor (_29680_, _29679_, _02519_);
  nor (_29681_, _29680_, _29677_);
  nor (_29683_, _29681_, _02153_);
  or (_29684_, _29683_, _06188_);
  nor (_29685_, _29684_, _29669_);
  and (_29686_, _29679_, _06188_);
  nor (_29687_, _29686_, _29685_);
  nor (_29688_, _29687_, _02031_);
  nor (_29689_, _29657_, _02032_);
  nand (_29690_, _05120_, _04197_);
  and (_29691_, _29690_, _29689_);
  nor (_29692_, _29691_, _29688_);
  nor (_29693_, _29692_, _01765_);
  or (_29694_, _10898_, _09951_);
  nor (_29695_, _29657_, _02037_);
  and (_29696_, _29695_, _29694_);
  or (_29697_, _29696_, _01994_);
  nor (_29698_, _29697_, _29693_);
  nor (_29699_, _29663_, _01995_);
  or (_29700_, _29699_, _29698_);
  and (_29701_, _29700_, _03059_);
  and (_29702_, _10914_, _03864_);
  nor (_29704_, _29702_, _29657_);
  nor (_29705_, _29704_, _03059_);
  or (_29706_, _29705_, _29701_);
  and (_29707_, _29706_, _03061_);
  and (_29708_, _10792_, _03864_);
  nor (_29709_, _29708_, _29657_);
  nor (_29710_, _29709_, _03061_);
  or (_29711_, _29710_, _29707_);
  and (_29712_, _29711_, _02208_);
  nor (_29713_, _29712_, _29666_);
  nor (_29715_, _29713_, _02342_);
  and (_29716_, _10791_, _03864_);
  or (_29717_, _29716_, _29657_);
  and (_29718_, _29717_, _02342_);
  or (_29719_, _29718_, _29715_);
  and (_29720_, _29719_, _04953_);
  not (_29721_, _03864_);
  nor (_29722_, _10913_, _29721_);
  nor (_29723_, _29722_, _29657_);
  nor (_29724_, _29723_, _04953_);
  or (_29727_, _29724_, _29720_);
  and (_29728_, _29727_, _04958_);
  nor (_29729_, _10789_, _09951_);
  nor (_29730_, _29729_, _29657_);
  nor (_29731_, _29730_, _04958_);
  nor (_29732_, _29731_, _15890_);
  not (_29733_, _29732_);
  nor (_29734_, _29733_, _29728_);
  nor (_29735_, _29734_, _29661_);
  or (_29736_, _29735_, _39633_);
  or (_29738_, _39632_, \oc8051_golden_model_1.TL1 [0]);
  and (_29739_, _29738_, _39026_);
  and (_41775_, _29739_, _29736_);
  nor (_29740_, _03864_, \oc8051_golden_model_1.TL1 [1]);
  not (_29741_, _29740_);
  or (_29742_, _10988_, _29721_);
  and (_29743_, _29742_, _02206_);
  and (_29744_, _29743_, _29741_);
  or (_29745_, _11113_, _29721_);
  and (_29746_, _29745_, _02331_);
  and (_29748_, _29746_, _29741_);
  not (_29749_, \oc8051_golden_model_1.TL1 [1]);
  nor (_29750_, _03864_, _29749_);
  nor (_29751_, _09951_, _03161_);
  nor (_29752_, _29751_, _29750_);
  and (_29753_, _29752_, _06188_);
  and (_29754_, _03864_, \oc8051_golden_model_1.ACC [1]);
  or (_29755_, _29754_, _29750_);
  and (_29756_, _29755_, _02062_);
  nor (_29757_, _02062_, _29749_);
  or (_29759_, _29757_, _29756_);
  and (_29760_, _29759_, _03006_);
  and (_29761_, _11001_, _03864_);
  nor (_29762_, _29761_, _29740_);
  and (_29763_, _29762_, _02158_);
  or (_29764_, _29763_, _29760_);
  and (_29765_, _29764_, _02519_);
  nor (_29766_, _29752_, _02519_);
  nor (_29767_, _29766_, _29765_);
  nor (_29768_, _29767_, _02153_);
  and (_29770_, _29755_, _02153_);
  nor (_29771_, _29770_, _06188_);
  not (_29772_, _29771_);
  nor (_29773_, _29772_, _29768_);
  nor (_29774_, _29773_, _29753_);
  nor (_29775_, _29774_, _02031_);
  nor (_29776_, _29775_, _01765_);
  nor (_29777_, _29750_, _02032_);
  nand (_29778_, _05075_, _04197_);
  nand (_29779_, _29778_, _29777_);
  and (_29781_, _29779_, _29776_);
  nand (_29782_, _11096_, _03864_);
  and (_29783_, _29782_, _01765_);
  and (_29784_, _29783_, _29741_);
  nor (_29785_, _29784_, _29781_);
  nor (_29786_, _29785_, _07629_);
  nor (_29787_, _10989_, _09951_);
  nor (_29788_, _29787_, _03059_);
  and (_29789_, _04197_, _02893_);
  nor (_29790_, _29789_, _01995_);
  nor (_29792_, _29790_, _29788_);
  nor (_29793_, _29792_, _29740_);
  nor (_29794_, _29793_, _29786_);
  nor (_29795_, _29794_, _02331_);
  nor (_29796_, _29795_, _29748_);
  nor (_29797_, _29796_, _02206_);
  nor (_29798_, _29797_, _29744_);
  nor (_29799_, _29798_, _02342_);
  nor (_29800_, _29750_, _04209_);
  nor (_29801_, _29800_, _03065_);
  and (_29803_, _29801_, _29755_);
  nor (_29804_, _29803_, _29799_);
  or (_29805_, _29804_, _17216_);
  and (_29806_, _11112_, _03864_);
  nor (_29807_, _29806_, _04958_);
  and (_29808_, _29807_, _29741_);
  nor (_29809_, _29808_, _02366_);
  and (_29810_, _29789_, _04208_);
  or (_29811_, _29740_, _04953_);
  or (_29812_, _29811_, _29810_);
  and (_29814_, _29812_, _29809_);
  and (_29815_, _29814_, _29805_);
  nor (_29816_, _29762_, _02778_);
  nor (_29817_, _29816_, _29815_);
  nor (_29818_, _29817_, _02081_);
  nor (_29819_, _29761_, _29750_);
  and (_29820_, _29819_, _02081_);
  nor (_29821_, _29820_, _29818_);
  or (_29822_, _29821_, _39633_);
  or (_29823_, _39632_, \oc8051_golden_model_1.TL1 [1]);
  and (_29825_, _29823_, _39026_);
  and (_41776_, _29825_, _29822_);
  not (_29826_, \oc8051_golden_model_1.TL1 [2]);
  nor (_29827_, _03864_, _29826_);
  nor (_29828_, _11314_, _09951_);
  nor (_29829_, _29828_, _29827_);
  nor (_29830_, _29829_, _04958_);
  and (_29831_, _11315_, _04197_);
  nor (_29832_, _29831_, _29827_);
  nor (_29833_, _29832_, _03061_);
  and (_29835_, _03864_, _04866_);
  nor (_29836_, _29835_, _29827_);
  and (_29837_, _29836_, _01994_);
  and (_29838_, _03864_, \oc8051_golden_model_1.ACC [2]);
  nor (_29839_, _29838_, _29827_);
  nor (_29840_, _29839_, _02549_);
  nor (_29841_, _29839_, _02063_);
  nor (_29842_, _02062_, _29826_);
  or (_29843_, _29842_, _29841_);
  and (_29844_, _29843_, _03006_);
  nor (_29845_, _11199_, _09951_);
  nor (_29846_, _29845_, _29827_);
  nor (_29847_, _29846_, _03006_);
  or (_29848_, _29847_, _29844_);
  and (_29849_, _29848_, _02519_);
  nor (_29850_, _09951_, _03624_);
  nor (_29851_, _29850_, _29827_);
  nor (_29852_, _29851_, _02519_);
  nor (_29853_, _29852_, _29849_);
  nor (_29854_, _29853_, _02153_);
  or (_29856_, _29854_, _06188_);
  nor (_29857_, _29856_, _29840_);
  and (_29858_, _29851_, _06188_);
  nor (_29859_, _29858_, _29857_);
  nor (_29860_, _29859_, _02031_);
  nor (_29861_, _29827_, _02032_);
  nand (_29862_, _05211_, _04197_);
  and (_29863_, _29862_, _29861_);
  or (_29864_, _29863_, _01765_);
  nor (_29865_, _29864_, _29860_);
  nor (_29867_, _11298_, _29721_);
  nor (_29868_, _29867_, _29827_);
  nor (_29869_, _29868_, _02037_);
  or (_29870_, _29869_, _01994_);
  nor (_29871_, _29870_, _29865_);
  nor (_29872_, _29871_, _29837_);
  or (_29873_, _29872_, _02210_);
  and (_29874_, _11189_, _03864_);
  or (_29875_, _29874_, _29827_);
  or (_29876_, _29875_, _03059_);
  and (_29878_, _29876_, _03061_);
  and (_29879_, _29878_, _29873_);
  nor (_29880_, _29879_, _29833_);
  nor (_29881_, _29880_, _02206_);
  nor (_29882_, _29827_, _04309_);
  not (_29883_, _29882_);
  nor (_29884_, _29836_, _02208_);
  and (_29885_, _29884_, _29883_);
  nor (_29886_, _29885_, _29881_);
  nor (_29887_, _29886_, _02342_);
  or (_29889_, _29882_, _03065_);
  nor (_29890_, _29889_, _29839_);
  or (_29891_, _29890_, _02202_);
  nor (_29892_, _29891_, _29887_);
  or (_29893_, _11187_, _09951_);
  nor (_29894_, _29827_, _04953_);
  and (_29895_, _29894_, _29893_);
  or (_29896_, _29895_, _02334_);
  nor (_29897_, _29896_, _29892_);
  nor (_29898_, _29897_, _29830_);
  nor (_29900_, _29898_, _02366_);
  nor (_29901_, _29846_, _02778_);
  or (_29902_, _29901_, _02081_);
  nor (_29903_, _29902_, _29900_);
  and (_29904_, _11367_, _03864_);
  nor (_29905_, _29904_, _29827_);
  and (_29906_, _29905_, _02081_);
  nor (_29907_, _29906_, _29903_);
  or (_29908_, _29907_, _39633_);
  or (_29909_, _39632_, \oc8051_golden_model_1.TL1 [2]);
  and (_29911_, _29909_, _39026_);
  and (_41777_, _29911_, _29908_);
  not (_29912_, \oc8051_golden_model_1.TL1 [3]);
  nor (_29913_, _03864_, _29912_);
  nor (_29914_, _11510_, _09951_);
  nor (_29915_, _29914_, _29913_);
  nor (_29916_, _29915_, _04958_);
  and (_29917_, _11511_, _04197_);
  nor (_29918_, _29917_, _29913_);
  nor (_29919_, _29918_, _03061_);
  nor (_29921_, _09951_, _03434_);
  nor (_29922_, _29921_, _29913_);
  and (_29923_, _29922_, _06188_);
  and (_29924_, _03864_, \oc8051_golden_model_1.ACC [3]);
  nor (_29925_, _29924_, _29913_);
  nor (_29926_, _29925_, _02063_);
  nor (_29927_, _02062_, _29912_);
  or (_29928_, _29927_, _29926_);
  and (_29929_, _29928_, _03006_);
  nor (_29930_, _11394_, _09951_);
  nor (_29932_, _29930_, _29913_);
  nor (_29933_, _29932_, _03006_);
  or (_29934_, _29933_, _29929_);
  and (_29935_, _29934_, _02519_);
  nor (_29936_, _29922_, _02519_);
  nor (_29937_, _29936_, _29935_);
  nor (_29938_, _29937_, _02153_);
  nor (_29939_, _29925_, _02549_);
  nor (_29940_, _29939_, _06188_);
  not (_29941_, _29940_);
  nor (_29943_, _29941_, _29938_);
  nor (_29944_, _29943_, _29923_);
  nor (_29945_, _29944_, _02031_);
  nor (_29946_, _29913_, _02032_);
  nand (_29947_, _05166_, _04197_);
  and (_29948_, _29947_, _29946_);
  or (_29949_, _29948_, _01765_);
  nor (_29950_, _29949_, _29945_);
  nor (_29951_, _11490_, _09951_);
  nor (_29952_, _29951_, _29913_);
  nor (_29954_, _29952_, _02037_);
  or (_29955_, _29954_, _07629_);
  or (_29956_, _29955_, _29950_);
  and (_29957_, _11505_, _04197_);
  or (_29958_, _29913_, _03059_);
  or (_29959_, _29958_, _29957_);
  and (_29960_, _03864_, _04719_);
  nor (_29961_, _29960_, _29913_);
  and (_29962_, _29961_, _01994_);
  nor (_29963_, _29962_, _02331_);
  and (_29965_, _29963_, _29959_);
  and (_29966_, _29965_, _29956_);
  nor (_29967_, _29966_, _29919_);
  nor (_29968_, _29967_, _02206_);
  nor (_29969_, _29913_, _04153_);
  not (_29970_, _29969_);
  nor (_29971_, _29961_, _02208_);
  and (_29972_, _29971_, _29970_);
  nor (_29973_, _29972_, _29968_);
  nor (_29974_, _29973_, _02342_);
  or (_29976_, _29969_, _03065_);
  nor (_29977_, _29976_, _29925_);
  or (_29978_, _29977_, _02202_);
  nor (_29979_, _29978_, _29974_);
  or (_29980_, _11503_, _09951_);
  nor (_29981_, _29913_, _04953_);
  and (_29982_, _29981_, _29980_);
  or (_29983_, _29982_, _02334_);
  nor (_29984_, _29983_, _29979_);
  nor (_29985_, _29984_, _29916_);
  nor (_29987_, _29985_, _02366_);
  nor (_29988_, _29932_, _02778_);
  or (_29989_, _29988_, _02081_);
  nor (_29990_, _29989_, _29987_);
  and (_29991_, _11567_, _03864_);
  nor (_29992_, _29991_, _29913_);
  and (_29993_, _29992_, _02081_);
  nor (_29994_, _29993_, _29990_);
  or (_29995_, _29994_, _39633_);
  or (_29996_, _39632_, \oc8051_golden_model_1.TL1 [3]);
  and (_29997_, _29996_, _39026_);
  and (_41778_, _29997_, _29995_);
  not (_29998_, \oc8051_golden_model_1.TL1 [4]);
  nor (_29999_, _03864_, _29998_);
  nor (_30000_, _11587_, _09951_);
  nor (_30001_, _30000_, _29999_);
  nor (_30002_, _30001_, _04958_);
  and (_30003_, _11588_, _04197_);
  nor (_30004_, _30003_, _29999_);
  nor (_30005_, _30004_, _03061_);
  and (_30007_, _05303_, _03864_);
  or (_30008_, _30007_, _29999_);
  and (_30009_, _30008_, _02031_);
  and (_30010_, _03864_, \oc8051_golden_model_1.ACC [4]);
  nor (_30011_, _30010_, _29999_);
  nor (_30012_, _30011_, _02549_);
  nor (_30013_, _30011_, _02063_);
  nor (_30014_, _02062_, _29998_);
  or (_30015_, _30014_, _30013_);
  and (_30016_, _30015_, _03006_);
  nor (_30018_, _11611_, _09951_);
  nor (_30019_, _30018_, _29999_);
  nor (_30020_, _30019_, _03006_);
  or (_30021_, _30020_, _30016_);
  and (_30022_, _30021_, _02519_);
  nor (_30023_, _04372_, _09951_);
  nor (_30024_, _30023_, _29999_);
  nor (_30025_, _30024_, _02519_);
  nor (_30026_, _30025_, _30022_);
  nor (_30027_, _30026_, _02153_);
  or (_30029_, _30027_, _06188_);
  nor (_30030_, _30029_, _30012_);
  and (_30031_, _30024_, _06188_);
  or (_30032_, _30031_, _02031_);
  nor (_30033_, _30032_, _30030_);
  or (_30034_, _30033_, _30009_);
  and (_30035_, _30034_, _02037_);
  nor (_30036_, _11704_, _09951_);
  nor (_30037_, _30036_, _29999_);
  nor (_30038_, _30037_, _02037_);
  or (_30040_, _30038_, _07629_);
  or (_30041_, _30040_, _30035_);
  and (_30042_, _11592_, _04197_);
  or (_30043_, _29999_, _03059_);
  or (_30044_, _30043_, _30042_);
  and (_30045_, _04831_, _03864_);
  nor (_30046_, _30045_, _29999_);
  and (_30047_, _30046_, _01994_);
  nor (_30048_, _30047_, _02331_);
  and (_30049_, _30048_, _30044_);
  and (_30051_, _30049_, _30041_);
  nor (_30052_, _30051_, _30005_);
  nor (_30053_, _30052_, _02206_);
  nor (_30054_, _29999_, _04420_);
  not (_30055_, _30054_);
  nor (_30056_, _30046_, _02208_);
  and (_30057_, _30056_, _30055_);
  nor (_30058_, _30057_, _30053_);
  nor (_30059_, _30058_, _02342_);
  or (_30060_, _30054_, _03065_);
  nor (_30062_, _30060_, _30011_);
  or (_30063_, _30062_, _02202_);
  nor (_30064_, _30063_, _30059_);
  or (_30065_, _11590_, _09951_);
  nor (_30066_, _29999_, _04953_);
  and (_30067_, _30066_, _30065_);
  or (_30068_, _30067_, _02334_);
  nor (_30069_, _30068_, _30064_);
  nor (_30070_, _30069_, _30002_);
  nor (_30071_, _30070_, _02366_);
  nor (_30073_, _30019_, _02778_);
  or (_30074_, _30073_, _02081_);
  nor (_30075_, _30074_, _30071_);
  and (_30076_, _11771_, _03864_);
  nor (_30077_, _30076_, _29999_);
  and (_30078_, _30077_, _02081_);
  nor (_30079_, _30078_, _30075_);
  or (_30080_, _30079_, _39633_);
  or (_30081_, _39632_, \oc8051_golden_model_1.TL1 [4]);
  and (_30082_, _30081_, _39026_);
  and (_41780_, _30082_, _30080_);
  not (_30084_, \oc8051_golden_model_1.TL1 [5]);
  nor (_30085_, _03864_, _30084_);
  nor (_30086_, _11785_, _09951_);
  nor (_30087_, _30086_, _30085_);
  nor (_30088_, _30087_, _04958_);
  and (_30089_, _11786_, _04197_);
  nor (_30090_, _30089_, _30085_);
  nor (_30091_, _30090_, _03061_);
  and (_30092_, _04827_, _03864_);
  nor (_30094_, _30092_, _30085_);
  and (_30095_, _30094_, _01994_);
  and (_30096_, _03864_, \oc8051_golden_model_1.ACC [5]);
  nor (_30097_, _30096_, _30085_);
  nor (_30098_, _30097_, _02549_);
  nor (_30099_, _30097_, _02063_);
  nor (_30100_, _02062_, _30084_);
  or (_30101_, _30100_, _30099_);
  and (_30102_, _30101_, _03006_);
  nor (_30103_, _11804_, _09951_);
  nor (_30105_, _30103_, _30085_);
  nor (_30106_, _30105_, _03006_);
  or (_30107_, _30106_, _30102_);
  and (_30108_, _30107_, _02519_);
  nor (_30109_, _04057_, _09951_);
  nor (_30110_, _30109_, _30085_);
  nor (_30111_, _30110_, _02519_);
  nor (_30112_, _30111_, _30108_);
  nor (_30113_, _30112_, _02153_);
  or (_30114_, _30113_, _06188_);
  nor (_30116_, _30114_, _30098_);
  and (_30117_, _30110_, _06188_);
  nor (_30118_, _30117_, _30116_);
  nor (_30119_, _30118_, _02031_);
  nor (_30120_, _30085_, _02032_);
  nand (_30121_, _05258_, _04197_);
  and (_30122_, _30121_, _30120_);
  or (_30123_, _30122_, _01765_);
  nor (_30124_, _30123_, _30119_);
  nor (_30125_, _11900_, _29721_);
  nor (_30127_, _30125_, _30085_);
  nor (_30128_, _30127_, _02037_);
  or (_30129_, _30128_, _01994_);
  nor (_30130_, _30129_, _30124_);
  nor (_30131_, _30130_, _30095_);
  or (_30132_, _30131_, _02210_);
  and (_30133_, _11915_, _03864_);
  or (_30134_, _30133_, _30085_);
  or (_30135_, _30134_, _03059_);
  and (_30136_, _30135_, _03061_);
  and (_30138_, _30136_, _30132_);
  nor (_30139_, _30138_, _30091_);
  nor (_30140_, _30139_, _02206_);
  nor (_30141_, _30085_, _04104_);
  not (_30142_, _30141_);
  nor (_30143_, _30094_, _02208_);
  and (_30144_, _30143_, _30142_);
  nor (_30145_, _30144_, _30140_);
  nor (_30146_, _30145_, _02342_);
  or (_30147_, _30141_, _03065_);
  nor (_30148_, _30147_, _30097_);
  or (_30149_, _30148_, _02202_);
  nor (_30150_, _30149_, _30146_);
  or (_30151_, _11913_, _09951_);
  nor (_30152_, _30085_, _04953_);
  and (_30153_, _30152_, _30151_);
  or (_30154_, _30153_, _02334_);
  nor (_30155_, _30154_, _30150_);
  nor (_30156_, _30155_, _30088_);
  nor (_30157_, _30156_, _02366_);
  nor (_30159_, _30105_, _02778_);
  or (_30160_, _30159_, _02081_);
  nor (_30161_, _30160_, _30157_);
  and (_30162_, _11974_, _03864_);
  nor (_30163_, _30162_, _30085_);
  and (_30164_, _30163_, _02081_);
  nor (_30165_, _30164_, _30161_);
  or (_30166_, _30165_, _39633_);
  or (_30167_, _39632_, \oc8051_golden_model_1.TL1 [5]);
  and (_30168_, _30167_, _39026_);
  and (_41781_, _30168_, _30166_);
  not (_30170_, \oc8051_golden_model_1.TL1 [6]);
  nor (_30171_, _03864_, _30170_);
  nor (_30172_, _12117_, _09951_);
  nor (_30173_, _30172_, _30171_);
  nor (_30174_, _30173_, _04958_);
  and (_30175_, _12118_, _04197_);
  nor (_30176_, _30175_, _30171_);
  nor (_30177_, _30176_, _03061_);
  and (_30178_, _12103_, _03864_);
  nor (_30180_, _30178_, _30171_);
  and (_30181_, _30180_, _01994_);
  and (_30182_, _03864_, \oc8051_golden_model_1.ACC [6]);
  nor (_30183_, _30182_, _30171_);
  nor (_30184_, _30183_, _02549_);
  nor (_30185_, _30183_, _02063_);
  nor (_30186_, _02062_, _30170_);
  or (_30187_, _30186_, _30185_);
  and (_30188_, _30187_, _03006_);
  nor (_30189_, _11993_, _09951_);
  nor (_30191_, _30189_, _30171_);
  nor (_30192_, _30191_, _03006_);
  or (_30193_, _30192_, _30188_);
  and (_30194_, _30193_, _02519_);
  nor (_30195_, _03964_, _09951_);
  nor (_30196_, _30195_, _30171_);
  nor (_30197_, _30196_, _02519_);
  nor (_30198_, _30197_, _30194_);
  nor (_30199_, _30198_, _02153_);
  or (_30200_, _30199_, _06188_);
  nor (_30202_, _30200_, _30184_);
  and (_30203_, _30196_, _06188_);
  nor (_30204_, _30203_, _30202_);
  nor (_30205_, _30204_, _02031_);
  nor (_30206_, _30171_, _02032_);
  nand (_30207_, _05029_, _04197_);
  and (_30208_, _30207_, _30206_);
  or (_30209_, _30208_, _01765_);
  nor (_30210_, _30209_, _30205_);
  nor (_30211_, _12096_, _29721_);
  nor (_30213_, _30211_, _30171_);
  nor (_30214_, _30213_, _02037_);
  or (_30215_, _30214_, _01994_);
  nor (_30216_, _30215_, _30210_);
  nor (_30217_, _30216_, _30181_);
  or (_30218_, _30217_, _02210_);
  and (_30219_, _12112_, _03864_);
  or (_30220_, _30219_, _30171_);
  or (_30221_, _30220_, _03059_);
  and (_30222_, _30221_, _03061_);
  and (_30224_, _30222_, _30218_);
  nor (_30225_, _30224_, _30177_);
  nor (_30226_, _30225_, _02206_);
  nor (_30227_, _30171_, _04011_);
  not (_30228_, _30227_);
  nor (_30229_, _30180_, _02208_);
  and (_30230_, _30229_, _30228_);
  nor (_30231_, _30230_, _30226_);
  nor (_30232_, _30231_, _02342_);
  or (_30233_, _30227_, _03065_);
  nor (_30235_, _30233_, _30183_);
  or (_30236_, _30235_, _02202_);
  nor (_30237_, _30236_, _30232_);
  or (_30238_, _12110_, _09951_);
  nor (_30239_, _30171_, _04953_);
  and (_30240_, _30239_, _30238_);
  or (_30241_, _30240_, _02334_);
  nor (_30242_, _30241_, _30237_);
  nor (_30243_, _30242_, _30174_);
  nor (_30244_, _30243_, _02366_);
  nor (_30246_, _30191_, _02778_);
  or (_30247_, _30246_, _02081_);
  nor (_30248_, _30247_, _30244_);
  and (_30249_, _12178_, _03864_);
  nor (_30250_, _30249_, _30171_);
  and (_30251_, _30250_, _02081_);
  nor (_30252_, _30251_, _30248_);
  or (_30253_, _30252_, _39633_);
  or (_30254_, _39632_, \oc8051_golden_model_1.TL1 [6]);
  and (_30255_, _30254_, _39026_);
  and (_41782_, _30255_, _30253_);
  not (_30257_, \oc8051_golden_model_1.TMOD [0]);
  nor (_30258_, _03878_, _30257_);
  nor (_30259_, _04257_, _10030_);
  nor (_30260_, _30259_, _30258_);
  and (_30261_, _30260_, _15890_);
  and (_30262_, _03878_, \oc8051_golden_model_1.ACC [0]);
  nor (_30263_, _30262_, _30258_);
  nor (_30264_, _30263_, _02549_);
  nor (_30265_, _30264_, _06188_);
  nor (_30267_, _30260_, _03006_);
  nor (_30268_, _02062_, _30257_);
  nor (_30269_, _30263_, _02063_);
  nor (_30270_, _30269_, _30268_);
  nor (_30271_, _30270_, _02158_);
  or (_30272_, _30271_, _02155_);
  nor (_30273_, _30272_, _30267_);
  or (_30274_, _30273_, _02153_);
  and (_30275_, _30274_, _30265_);
  and (_30276_, _03878_, _03002_);
  or (_30278_, _30258_, _24237_);
  nor (_30279_, _30278_, _30276_);
  nor (_30280_, _30279_, _30275_);
  nor (_30281_, _30280_, _02031_);
  and (_30282_, _05120_, _03878_);
  nor (_30283_, _30258_, _02032_);
  not (_30284_, _30283_);
  nor (_30285_, _30284_, _30282_);
  nor (_30286_, _30285_, _30281_);
  nor (_30287_, _30286_, _01765_);
  nor (_30289_, _10898_, _10030_);
  or (_30290_, _30258_, _02037_);
  nor (_30291_, _30290_, _30289_);
  or (_30292_, _30291_, _01994_);
  nor (_30293_, _30292_, _30287_);
  and (_30294_, _03878_, _04837_);
  nor (_30295_, _30294_, _30258_);
  nor (_30296_, _30295_, _01995_);
  or (_30297_, _30296_, _30293_);
  and (_30298_, _30297_, _03059_);
  and (_30300_, _10914_, _03878_);
  nor (_30301_, _30300_, _30258_);
  nor (_30302_, _30301_, _03059_);
  or (_30303_, _30302_, _30298_);
  and (_30304_, _30303_, _03061_);
  and (_30305_, _10792_, _03878_);
  nor (_30306_, _30305_, _30258_);
  nor (_30307_, _30306_, _03061_);
  or (_30308_, _30307_, _30304_);
  and (_30309_, _30308_, _02208_);
  or (_30310_, _30295_, _02208_);
  nor (_30311_, _30310_, _30259_);
  nor (_30312_, _30311_, _30309_);
  nor (_30313_, _30312_, _02342_);
  and (_30314_, _10791_, _03878_);
  or (_30315_, _30314_, _30258_);
  and (_30316_, _30315_, _02342_);
  or (_30317_, _30316_, _30313_);
  and (_30318_, _30317_, _04953_);
  nor (_30319_, _10913_, _10030_);
  nor (_30321_, _30319_, _30258_);
  nor (_30322_, _30321_, _04953_);
  or (_30323_, _30322_, _30318_);
  and (_30324_, _30323_, _04958_);
  nor (_30325_, _10789_, _10030_);
  nor (_30326_, _30325_, _30258_);
  nor (_30327_, _30326_, _04958_);
  nor (_30328_, _30327_, _15890_);
  not (_30329_, _30328_);
  nor (_30330_, _30329_, _30324_);
  nor (_30332_, _30330_, _30261_);
  or (_30333_, _30332_, _39633_);
  or (_30334_, _39632_, \oc8051_golden_model_1.TMOD [0]);
  and (_30335_, _30334_, _39026_);
  and (_41784_, _30335_, _30333_);
  nor (_30336_, _03878_, \oc8051_golden_model_1.TMOD [1]);
  not (_30337_, _30336_);
  nor (_30338_, _11113_, _10030_);
  nor (_30339_, _30338_, _03061_);
  and (_30340_, _30339_, _30337_);
  and (_30342_, _05075_, _03878_);
  not (_30343_, \oc8051_golden_model_1.TMOD [1]);
  nor (_30344_, _03878_, _30343_);
  nor (_30345_, _30344_, _02032_);
  not (_30346_, _30345_);
  nor (_30347_, _30346_, _30342_);
  not (_30348_, _30347_);
  nor (_30349_, _10030_, _03161_);
  nor (_30350_, _30349_, _30344_);
  and (_30351_, _30350_, _06188_);
  and (_30353_, _03878_, _01804_);
  nor (_30354_, _30353_, _30336_);
  and (_30355_, _30354_, _02062_);
  nor (_30356_, _02062_, _30343_);
  or (_30357_, _30356_, _30355_);
  and (_30358_, _30357_, _03006_);
  and (_30359_, _11001_, _03878_);
  nor (_30360_, _30359_, _30336_);
  and (_30361_, _30360_, _02158_);
  or (_30362_, _30361_, _30358_);
  and (_30364_, _30362_, _02519_);
  nor (_30365_, _30350_, _02519_);
  nor (_30366_, _30365_, _30364_);
  nor (_30367_, _30366_, _02153_);
  and (_30368_, _30354_, _02153_);
  nor (_30369_, _30368_, _06188_);
  not (_30370_, _30369_);
  nor (_30371_, _30370_, _30367_);
  nor (_30372_, _30371_, _30351_);
  nor (_30373_, _30372_, _02031_);
  nor (_30375_, _30373_, _01765_);
  and (_30376_, _30375_, _30348_);
  and (_30377_, _11096_, _03878_);
  nor (_30378_, _30377_, _02037_);
  and (_30379_, _30378_, _30337_);
  nor (_30380_, _30379_, _30376_);
  nor (_30381_, _30380_, _07629_);
  nor (_30382_, _10989_, _10030_);
  nor (_30383_, _30382_, _03059_);
  and (_30384_, _03878_, _02893_);
  nor (_30386_, _30384_, _01995_);
  or (_30387_, _30386_, _30383_);
  and (_30388_, _30387_, _30337_);
  nor (_30389_, _30388_, _30381_);
  nor (_30390_, _30389_, _02331_);
  nor (_30391_, _30390_, _30340_);
  nor (_30392_, _30391_, _02206_);
  nor (_30393_, _10988_, _10030_);
  nor (_30394_, _30393_, _02208_);
  and (_30395_, _30394_, _30337_);
  nor (_30397_, _30395_, _30392_);
  nor (_30398_, _30397_, _02342_);
  nor (_30399_, _30344_, _04209_);
  nor (_30400_, _30399_, _03065_);
  and (_30401_, _30400_, _30354_);
  nor (_30402_, _30401_, _30398_);
  or (_30403_, _30402_, _17216_);
  nand (_30404_, _30353_, _04208_);
  nor (_30405_, _30336_, _04958_);
  and (_30406_, _30405_, _30404_);
  nor (_30408_, _30406_, _02366_);
  and (_30409_, _30384_, _04208_);
  or (_30410_, _30336_, _04953_);
  or (_30411_, _30410_, _30409_);
  and (_30412_, _30411_, _30408_);
  and (_30413_, _30412_, _30403_);
  nor (_30414_, _30360_, _02778_);
  nor (_30415_, _30414_, _30413_);
  nor (_30416_, _30415_, _02081_);
  nor (_30417_, _30359_, _30344_);
  and (_30419_, _30417_, _02081_);
  nor (_30420_, _30419_, _30416_);
  or (_30421_, _30420_, _39633_);
  or (_30422_, _39632_, \oc8051_golden_model_1.TMOD [1]);
  and (_30423_, _30422_, _39026_);
  and (_41785_, _30423_, _30421_);
  not (_30424_, \oc8051_golden_model_1.TMOD [2]);
  nor (_30425_, _03878_, _30424_);
  nor (_30426_, _11314_, _10030_);
  nor (_30427_, _30426_, _30425_);
  nor (_30429_, _30427_, _04958_);
  and (_30430_, _05211_, _03878_);
  nor (_30431_, _30425_, _02032_);
  not (_30432_, _30431_);
  nor (_30433_, _30432_, _30430_);
  nor (_30434_, _10030_, _03624_);
  nor (_30435_, _30434_, _30425_);
  and (_30436_, _30435_, _06188_);
  nor (_30437_, _11199_, _10030_);
  nor (_30438_, _30437_, _30425_);
  nor (_30440_, _30438_, _03006_);
  nor (_30441_, _02062_, _30424_);
  and (_30442_, _03878_, \oc8051_golden_model_1.ACC [2]);
  nor (_30443_, _30442_, _30425_);
  nor (_30444_, _30443_, _02063_);
  nor (_30445_, _30444_, _30441_);
  nor (_30446_, _30445_, _02158_);
  or (_30447_, _30446_, _30440_);
  and (_30448_, _30447_, _02519_);
  nor (_30449_, _30435_, _02519_);
  or (_30451_, _30449_, _30448_);
  and (_30452_, _30451_, _02549_);
  nor (_30453_, _30443_, _02549_);
  nor (_30454_, _30453_, _06188_);
  not (_30455_, _30454_);
  nor (_30456_, _30455_, _30452_);
  nor (_30457_, _30456_, _30436_);
  nor (_30458_, _30457_, _02031_);
  nor (_30459_, _30458_, _30433_);
  nor (_30460_, _30459_, _01765_);
  nor (_30462_, _11298_, _10030_);
  or (_30463_, _30425_, _02037_);
  nor (_30464_, _30463_, _30462_);
  or (_30465_, _30464_, _01994_);
  nor (_30466_, _30465_, _30460_);
  and (_30467_, _03878_, _04866_);
  nor (_30468_, _30467_, _30425_);
  nor (_30469_, _30468_, _01995_);
  or (_30470_, _30469_, _30466_);
  and (_30471_, _30470_, _03059_);
  and (_30472_, _11189_, _03878_);
  nor (_30473_, _30472_, _30425_);
  nor (_30474_, _30473_, _03059_);
  or (_30475_, _30474_, _30471_);
  and (_30476_, _30475_, _03061_);
  and (_30477_, _11315_, _03878_);
  nor (_30478_, _30477_, _30425_);
  nor (_30479_, _30478_, _03061_);
  or (_30480_, _30479_, _30476_);
  and (_30481_, _30480_, _02208_);
  nor (_30483_, _30425_, _04309_);
  or (_30484_, _30468_, _02208_);
  nor (_30485_, _30484_, _30483_);
  nor (_30486_, _30485_, _30481_);
  nor (_30487_, _30486_, _02342_);
  or (_30488_, _30483_, _03065_);
  nor (_30489_, _30488_, _30443_);
  or (_30490_, _30489_, _02202_);
  nor (_30491_, _30490_, _30487_);
  nor (_30492_, _11187_, _10030_);
  or (_30494_, _30425_, _04953_);
  nor (_30495_, _30494_, _30492_);
  or (_30496_, _30495_, _02334_);
  nor (_30497_, _30496_, _30491_);
  nor (_30498_, _30497_, _30429_);
  nor (_30499_, _30498_, _02366_);
  nor (_30500_, _30438_, _02778_);
  or (_30501_, _30500_, _02081_);
  nor (_30502_, _30501_, _30499_);
  and (_30503_, _11367_, _03878_);
  nor (_30505_, _30503_, _30425_);
  and (_30506_, _30505_, _02081_);
  nor (_30507_, _30506_, _30502_);
  or (_30508_, _30507_, _39633_);
  or (_30509_, _39632_, \oc8051_golden_model_1.TMOD [2]);
  and (_30510_, _30509_, _39026_);
  and (_41786_, _30510_, _30508_);
  not (_30511_, \oc8051_golden_model_1.TMOD [3]);
  nor (_30512_, _03878_, _30511_);
  nor (_30513_, _11510_, _10030_);
  nor (_30515_, _30513_, _30512_);
  nor (_30516_, _30515_, _04958_);
  and (_30517_, _11511_, _03878_);
  nor (_30518_, _30517_, _30512_);
  nor (_30519_, _30518_, _03061_);
  nor (_30520_, _10030_, _03434_);
  nor (_30521_, _30520_, _30512_);
  and (_30522_, _30521_, _06188_);
  and (_30523_, _03878_, \oc8051_golden_model_1.ACC [3]);
  nor (_30524_, _30523_, _30512_);
  nor (_30526_, _30524_, _02063_);
  nor (_30527_, _02062_, _30511_);
  or (_30528_, _30527_, _30526_);
  and (_30529_, _30528_, _03006_);
  nor (_30530_, _11394_, _10030_);
  nor (_30531_, _30530_, _30512_);
  nor (_30532_, _30531_, _03006_);
  or (_30533_, _30532_, _30529_);
  and (_30534_, _30533_, _02519_);
  nor (_30535_, _30521_, _02519_);
  nor (_30537_, _30535_, _30534_);
  nor (_30538_, _30537_, _02153_);
  nor (_30539_, _30524_, _02549_);
  nor (_30540_, _30539_, _06188_);
  not (_30541_, _30540_);
  nor (_30542_, _30541_, _30538_);
  nor (_30543_, _30542_, _30522_);
  nor (_30544_, _30543_, _02031_);
  and (_30545_, _05166_, _03878_);
  nor (_30546_, _30512_, _02032_);
  not (_30548_, _30546_);
  nor (_30549_, _30548_, _30545_);
  nor (_30550_, _30549_, _01765_);
  not (_30551_, _30550_);
  nor (_30552_, _30551_, _30544_);
  nor (_30553_, _11490_, _10030_);
  nor (_30554_, _30553_, _30512_);
  nor (_30555_, _30554_, _02037_);
  or (_30556_, _30555_, _07629_);
  or (_30557_, _30556_, _30552_);
  and (_30559_, _11505_, _03878_);
  or (_30560_, _30512_, _03059_);
  or (_30561_, _30560_, _30559_);
  and (_30562_, _03878_, _04719_);
  nor (_30563_, _30562_, _30512_);
  and (_30564_, _30563_, _01994_);
  nor (_30565_, _30564_, _02331_);
  and (_30566_, _30565_, _30561_);
  and (_30567_, _30566_, _30557_);
  nor (_30568_, _30567_, _30519_);
  nor (_30570_, _30568_, _02206_);
  nor (_30571_, _30512_, _04153_);
  not (_30572_, _30571_);
  nor (_30573_, _30563_, _02208_);
  and (_30574_, _30573_, _30572_);
  nor (_30575_, _30574_, _30570_);
  nor (_30576_, _30575_, _02342_);
  or (_30577_, _30571_, _03065_);
  nor (_30578_, _30577_, _30524_);
  or (_30579_, _30578_, _02202_);
  nor (_30581_, _30579_, _30576_);
  nor (_30582_, _11503_, _10030_);
  or (_30583_, _30512_, _04953_);
  nor (_30584_, _30583_, _30582_);
  or (_30585_, _30584_, _02334_);
  nor (_30586_, _30585_, _30581_);
  nor (_30587_, _30586_, _30516_);
  nor (_30588_, _30587_, _02366_);
  nor (_30589_, _30531_, _02778_);
  or (_30590_, _30589_, _02081_);
  nor (_30592_, _30590_, _30588_);
  and (_30593_, _11567_, _03878_);
  nor (_30594_, _30593_, _30512_);
  and (_30595_, _30594_, _02081_);
  nor (_30596_, _30595_, _30592_);
  or (_30597_, _30596_, _39633_);
  or (_30598_, _39632_, \oc8051_golden_model_1.TMOD [3]);
  and (_30599_, _30598_, _39026_);
  and (_41787_, _30599_, _30597_);
  not (_30600_, \oc8051_golden_model_1.TMOD [4]);
  nor (_30602_, _03878_, _30600_);
  nor (_30603_, _11587_, _10030_);
  nor (_30604_, _30603_, _30602_);
  nor (_30605_, _30604_, _04958_);
  and (_30606_, _11588_, _03878_);
  nor (_30607_, _30606_, _30602_);
  nor (_30608_, _30607_, _03061_);
  and (_30609_, _05303_, _03878_);
  or (_30610_, _30609_, _30602_);
  and (_30611_, _30610_, _02031_);
  and (_30613_, _03878_, \oc8051_golden_model_1.ACC [4]);
  nor (_30614_, _30613_, _30602_);
  nor (_30615_, _30614_, _02063_);
  nor (_30616_, _02062_, _30600_);
  or (_30617_, _30616_, _30615_);
  and (_30618_, _30617_, _03006_);
  nor (_30619_, _11611_, _10030_);
  nor (_30620_, _30619_, _30602_);
  nor (_30621_, _30620_, _03006_);
  or (_30622_, _30621_, _30618_);
  and (_30624_, _30622_, _02519_);
  nor (_30625_, _04372_, _10030_);
  nor (_30626_, _30625_, _30602_);
  nor (_30627_, _30626_, _02519_);
  nor (_30628_, _30627_, _30624_);
  nor (_30629_, _30628_, _02153_);
  nor (_30630_, _30614_, _02549_);
  nor (_30631_, _30630_, _06188_);
  not (_30632_, _30631_);
  nor (_30633_, _30632_, _30629_);
  and (_30634_, _30626_, _06188_);
  or (_30635_, _30634_, _02031_);
  nor (_30636_, _30635_, _30633_);
  or (_30637_, _30636_, _30611_);
  and (_30638_, _30637_, _02037_);
  nor (_30639_, _11704_, _10030_);
  nor (_30640_, _30639_, _30602_);
  nor (_30641_, _30640_, _02037_);
  or (_30642_, _30641_, _07629_);
  or (_30643_, _30642_, _30638_);
  and (_30645_, _11592_, _03878_);
  or (_30646_, _30602_, _03059_);
  or (_30647_, _30646_, _30645_);
  and (_30648_, _04831_, _03878_);
  nor (_30649_, _30648_, _30602_);
  and (_30650_, _30649_, _01994_);
  nor (_30651_, _30650_, _02331_);
  and (_30652_, _30651_, _30647_);
  and (_30653_, _30652_, _30643_);
  nor (_30654_, _30653_, _30608_);
  nor (_30656_, _30654_, _02206_);
  nor (_30657_, _30602_, _04420_);
  not (_30658_, _30657_);
  nor (_30659_, _30649_, _02208_);
  and (_30660_, _30659_, _30658_);
  nor (_30661_, _30660_, _30656_);
  nor (_30662_, _30661_, _02342_);
  or (_30663_, _30657_, _03065_);
  nor (_30664_, _30663_, _30614_);
  or (_30665_, _30664_, _02202_);
  nor (_30667_, _30665_, _30662_);
  nor (_30668_, _11590_, _10030_);
  or (_30669_, _30602_, _04953_);
  nor (_30670_, _30669_, _30668_);
  or (_30671_, _30670_, _02334_);
  nor (_30672_, _30671_, _30667_);
  nor (_30673_, _30672_, _30605_);
  nor (_30674_, _30673_, _02366_);
  nor (_30675_, _30620_, _02778_);
  or (_30676_, _30675_, _02081_);
  nor (_30678_, _30676_, _30674_);
  and (_30679_, _11771_, _03878_);
  nor (_30680_, _30679_, _30602_);
  and (_30681_, _30680_, _02081_);
  nor (_30682_, _30681_, _30678_);
  or (_30683_, _30682_, _39633_);
  or (_30684_, _39632_, \oc8051_golden_model_1.TMOD [4]);
  and (_30685_, _30684_, _39026_);
  and (_41788_, _30685_, _30683_);
  not (_30686_, \oc8051_golden_model_1.TMOD [5]);
  nor (_30688_, _03878_, _30686_);
  nor (_30689_, _11785_, _10030_);
  nor (_30690_, _30689_, _30688_);
  nor (_30691_, _30690_, _04958_);
  and (_30692_, _11786_, _03878_);
  nor (_30693_, _30692_, _30688_);
  nor (_30694_, _30693_, _03061_);
  and (_30695_, _04827_, _03878_);
  nor (_30696_, _30695_, _30688_);
  and (_30697_, _30696_, _01994_);
  nor (_30699_, _04057_, _10030_);
  nor (_30700_, _30699_, _30688_);
  and (_30701_, _30700_, _06188_);
  and (_30702_, _03878_, \oc8051_golden_model_1.ACC [5]);
  nor (_30703_, _30702_, _30688_);
  nor (_30704_, _30703_, _02063_);
  nor (_30705_, _02062_, _30686_);
  or (_30706_, _30705_, _30704_);
  and (_30707_, _30706_, _03006_);
  nor (_30708_, _11804_, _10030_);
  nor (_30710_, _30708_, _30688_);
  nor (_30711_, _30710_, _03006_);
  or (_30712_, _30711_, _30707_);
  and (_30713_, _30712_, _02519_);
  nor (_30714_, _30700_, _02519_);
  nor (_30715_, _30714_, _30713_);
  nor (_30716_, _30715_, _02153_);
  nor (_30717_, _30703_, _02549_);
  nor (_30718_, _30717_, _06188_);
  not (_30719_, _30718_);
  nor (_30721_, _30719_, _30716_);
  nor (_30722_, _30721_, _30701_);
  nor (_30723_, _30722_, _02031_);
  and (_30724_, _05258_, _03878_);
  nor (_30725_, _30688_, _02032_);
  not (_30726_, _30725_);
  nor (_30727_, _30726_, _30724_);
  or (_30728_, _30727_, _01765_);
  nor (_30729_, _30728_, _30723_);
  nor (_30730_, _11900_, _10030_);
  nor (_30732_, _30730_, _30688_);
  nor (_30733_, _30732_, _02037_);
  or (_30734_, _30733_, _01994_);
  nor (_30735_, _30734_, _30729_);
  nor (_30736_, _30735_, _30697_);
  or (_30737_, _30736_, _02210_);
  and (_30738_, _11915_, _03878_);
  or (_30739_, _30738_, _30688_);
  or (_30740_, _30739_, _03059_);
  and (_30741_, _30740_, _03061_);
  and (_30743_, _30741_, _30737_);
  nor (_30744_, _30743_, _30694_);
  nor (_30745_, _30744_, _02206_);
  nor (_30746_, _30688_, _04104_);
  not (_30747_, _30746_);
  nor (_30748_, _30696_, _02208_);
  and (_30749_, _30748_, _30747_);
  nor (_30750_, _30749_, _30745_);
  nor (_30751_, _30750_, _02342_);
  or (_30752_, _30746_, _03065_);
  nor (_30754_, _30752_, _30703_);
  or (_30755_, _30754_, _02202_);
  nor (_30756_, _30755_, _30751_);
  nor (_30757_, _11913_, _10030_);
  or (_30758_, _30688_, _04953_);
  nor (_30759_, _30758_, _30757_);
  or (_30760_, _30759_, _02334_);
  nor (_30761_, _30760_, _30756_);
  nor (_30762_, _30761_, _30691_);
  nor (_30763_, _30762_, _02366_);
  nor (_30765_, _30710_, _02778_);
  or (_30766_, _30765_, _02081_);
  nor (_30767_, _30766_, _30763_);
  and (_30768_, _11974_, _03878_);
  nor (_30769_, _30768_, _30688_);
  and (_30770_, _30769_, _02081_);
  nor (_30771_, _30770_, _30767_);
  or (_30772_, _30771_, _39633_);
  or (_30773_, _39632_, \oc8051_golden_model_1.TMOD [5]);
  and (_30774_, _30773_, _39026_);
  and (_41789_, _30774_, _30772_);
  not (_30776_, \oc8051_golden_model_1.TMOD [6]);
  nor (_30777_, _03878_, _30776_);
  nor (_30778_, _12117_, _10030_);
  nor (_30779_, _30778_, _30777_);
  nor (_30780_, _30779_, _04958_);
  and (_30781_, _12118_, _03878_);
  nor (_30782_, _30781_, _30777_);
  nor (_30783_, _30782_, _03061_);
  and (_30784_, _12103_, _03878_);
  nor (_30786_, _30784_, _30777_);
  and (_30787_, _30786_, _01994_);
  and (_30788_, _03878_, \oc8051_golden_model_1.ACC [6]);
  nor (_30789_, _30788_, _30777_);
  nor (_30790_, _30789_, _02549_);
  nor (_30791_, _30789_, _02063_);
  nor (_30792_, _02062_, _30776_);
  or (_30793_, _30792_, _30791_);
  and (_30794_, _30793_, _03006_);
  nor (_30795_, _11993_, _10030_);
  nor (_30796_, _30795_, _30777_);
  nor (_30797_, _30796_, _03006_);
  or (_30798_, _30797_, _30794_);
  and (_30799_, _30798_, _02519_);
  nor (_30800_, _03964_, _10030_);
  nor (_30801_, _30800_, _30777_);
  nor (_30802_, _30801_, _02519_);
  nor (_30803_, _30802_, _30799_);
  nor (_30804_, _30803_, _02153_);
  or (_30805_, _30804_, _06188_);
  nor (_30807_, _30805_, _30790_);
  and (_30808_, _30801_, _06188_);
  nor (_30809_, _30808_, _30807_);
  nor (_30810_, _30809_, _02031_);
  and (_30811_, _05029_, _03878_);
  nor (_30812_, _30777_, _02032_);
  not (_30813_, _30812_);
  nor (_30814_, _30813_, _30811_);
  or (_30815_, _30814_, _01765_);
  nor (_30816_, _30815_, _30810_);
  nor (_30818_, _12096_, _10030_);
  nor (_30819_, _30818_, _30777_);
  nor (_30820_, _30819_, _02037_);
  or (_30821_, _30820_, _01994_);
  nor (_30822_, _30821_, _30816_);
  nor (_30823_, _30822_, _30787_);
  or (_30824_, _30823_, _02210_);
  and (_30825_, _12112_, _03878_);
  or (_30826_, _30825_, _30777_);
  or (_30827_, _30826_, _03059_);
  and (_30829_, _30827_, _03061_);
  and (_30830_, _30829_, _30824_);
  nor (_30831_, _30830_, _30783_);
  nor (_30832_, _30831_, _02206_);
  nor (_30833_, _30777_, _04011_);
  not (_30834_, _30833_);
  nor (_30835_, _30786_, _02208_);
  and (_30836_, _30835_, _30834_);
  nor (_30837_, _30836_, _30832_);
  nor (_30838_, _30837_, _02342_);
  or (_30840_, _30833_, _03065_);
  nor (_30841_, _30840_, _30789_);
  or (_30842_, _30841_, _02202_);
  nor (_30843_, _30842_, _30838_);
  nor (_30844_, _12110_, _10030_);
  or (_30845_, _30777_, _04953_);
  nor (_30846_, _30845_, _30844_);
  or (_30847_, _30846_, _02334_);
  nor (_30848_, _30847_, _30843_);
  nor (_30849_, _30848_, _30780_);
  nor (_30851_, _30849_, _02366_);
  nor (_30852_, _30796_, _02778_);
  or (_30853_, _30852_, _02081_);
  nor (_30854_, _30853_, _30851_);
  and (_30855_, _12178_, _03878_);
  nor (_30856_, _30855_, _30777_);
  and (_30857_, _30856_, _02081_);
  nor (_30858_, _30857_, _30854_);
  or (_30859_, _30858_, _39633_);
  or (_30860_, _39632_, \oc8051_golden_model_1.TMOD [6]);
  and (_30862_, _30860_, _39026_);
  and (_41790_, _30862_, _30859_);
  not (_30863_, _23330_);
  and (_30864_, _30863_, _02679_);
  and (_30865_, _10747_, _10751_);
  nor (_30866_, _30865_, _01439_);
  and (_30867_, _10722_, _07581_);
  nor (_30868_, _30867_, _01439_);
  and (_30869_, _10118_, _07534_);
  nor (_30870_, _30869_, _01439_);
  and (_30872_, _06781_, \oc8051_golden_model_1.PC [0]);
  nor (_30873_, _06781_, \oc8051_golden_model_1.PC [0]);
  nor (_30874_, _30873_, _30872_);
  and (_30875_, _30874_, _10122_);
  not (_30876_, _01736_);
  and (_30877_, _10133_, _04953_);
  nor (_30878_, _30877_, _01439_);
  not (_30879_, _01728_);
  and (_30880_, _10139_, _02208_);
  nor (_30881_, _30880_, _01439_);
  not (_30883_, _01722_);
  and (_30884_, _10147_, _03059_);
  nor (_30885_, _30884_, _01439_);
  and (_30886_, _01994_, _01439_);
  nor (_30887_, _02218_, _01765_);
  and (_30888_, _30887_, _10542_);
  nor (_30889_, _30888_, _01439_);
  nor (_30890_, _02679_, _01755_);
  nor (_30891_, _10158_, _01439_);
  nor (_30892_, _02679_, _01750_);
  nor (_30894_, _02679_, _01757_);
  and (_30895_, _01752_, _01747_);
  or (_30896_, _30895_, _02679_);
  and (_30897_, _10299_, _06859_);
  nor (_30898_, _30897_, _01439_);
  or (_30899_, _30898_, _10323_);
  nor (_30900_, _10312_, _01439_);
  and (_30901_, _10312_, _01439_);
  nor (_30902_, _30901_, _30900_);
  and (_30903_, _30902_, _01747_);
  not (_30905_, _30903_);
  and (_30906_, _30905_, _30897_);
  or (_30907_, _30906_, _30899_);
  and (_30908_, _30907_, _04534_);
  and (_30909_, _30908_, _30896_);
  and (_30910_, _10435_, \oc8051_golden_model_1.PC [0]);
  and (_30911_, _02027_, _01439_);
  nor (_30912_, _30911_, _10380_);
  and (_30913_, _30912_, _10437_);
  or (_30914_, _30913_, _30910_);
  nor (_30916_, _30914_, _04534_);
  nor (_30917_, _30916_, _30909_);
  nor (_30918_, _30917_, _02079_);
  and (_30919_, _02079_, \oc8051_golden_model_1.PC [0]);
  nor (_30920_, _30919_, _30918_);
  and (_30921_, _30920_, _03006_);
  not (_30922_, _30921_);
  and (_30923_, _02679_, \oc8051_golden_model_1.PC [0]);
  nor (_30924_, _30923_, _10228_);
  not (_30925_, _30924_);
  and (_30927_, _30925_, _10295_);
  and (_30928_, _04257_, _04152_);
  and (_30929_, _30928_, _10292_);
  nand (_30930_, _30929_, _11196_);
  nor (_30931_, _30930_, _01439_);
  or (_30932_, _30931_, _03006_);
  or (_30933_, _30932_, _30927_);
  and (_30934_, _30933_, _10287_);
  and (_30935_, _30934_, _30922_);
  nor (_30936_, _10287_, _01439_);
  nor (_30938_, _30936_, _03446_);
  not (_30939_, _30938_);
  nor (_30940_, _30939_, _30935_);
  nor (_30941_, _02679_, _01745_);
  and (_30942_, _10460_, _10452_);
  not (_30943_, _30942_);
  nor (_30944_, _30943_, _30941_);
  not (_30945_, _30944_);
  nor (_30946_, _30945_, _30940_);
  nor (_30947_, _30942_, _01439_);
  nor (_30949_, _30947_, _10464_);
  not (_30950_, _30949_);
  nor (_30951_, _30950_, _30946_);
  or (_30952_, _30951_, _10475_);
  nor (_30953_, _30952_, _30894_);
  and (_30954_, _08770_, _01439_);
  nor (_30955_, _30925_, _08770_);
  or (_30956_, _30955_, _10471_);
  nor (_30957_, _30956_, _30954_);
  or (_30958_, _30957_, _08790_);
  nor (_30959_, _30958_, _30953_);
  or (_30960_, _10482_, _01439_);
  or (_30961_, _30924_, _08842_);
  and (_30962_, _30961_, _08790_);
  and (_30963_, _30962_, _30960_);
  or (_30964_, _30963_, _30959_);
  and (_30965_, _30964_, _02547_);
  and (_30966_, _08877_, _01439_);
  nor (_30967_, _30925_, _08877_);
  nor (_30968_, _30967_, _30966_);
  nor (_30970_, _30968_, _02547_);
  nor (_30971_, _30970_, _30965_);
  nor (_30972_, _30971_, _02246_);
  and (_30973_, _08922_, _01439_);
  nor (_30974_, _30925_, _08922_);
  or (_30975_, _30974_, _30973_);
  and (_30976_, _30975_, _02246_);
  or (_30977_, _30976_, _30972_);
  and (_30978_, _30977_, _08882_);
  and (_30979_, _08881_, _01439_);
  or (_30981_, _30979_, _30978_);
  and (_30982_, _30981_, _01750_);
  or (_30983_, _30982_, _10159_);
  nor (_30984_, _30983_, _30892_);
  or (_30985_, _30984_, _10513_);
  nor (_30986_, _30985_, _30891_);
  and (_30987_, _10153_, _01778_);
  not (_30988_, _30987_);
  or (_30989_, _30988_, _30986_);
  nor (_30990_, _30989_, _30890_);
  nor (_30992_, _30987_, _01439_);
  nor (_30993_, _30992_, _01767_);
  not (_30994_, _30993_);
  nor (_30995_, _30994_, _30990_);
  nor (_30996_, _02679_, _04460_);
  not (_30997_, _30888_);
  nor (_30998_, _30997_, _30996_);
  not (_30999_, _30998_);
  nor (_31000_, _30999_, _30995_);
  or (_31001_, _31000_, _01711_);
  nor (_31003_, _31001_, _30889_);
  nor (_31004_, _02679_, _01712_);
  or (_31005_, _31004_, _10550_);
  nor (_31006_, _31005_, _31003_);
  nor (_31007_, _30912_, _10551_);
  nor (_31008_, _31007_, _31006_);
  and (_31009_, _31008_, _01995_);
  or (_31010_, _31009_, _30886_);
  and (_31011_, _31010_, _10150_);
  and (_31012_, _10149_, _01878_);
  or (_31014_, _31012_, _31011_);
  and (_31015_, _31014_, _03308_);
  nor (_31016_, _02679_, _03308_);
  or (_31017_, _31016_, _31015_);
  and (_31018_, _31017_, _10605_);
  not (_31019_, _30884_);
  nor (_31020_, _30912_, _07587_);
  and (_31021_, _07587_, _01439_);
  nor (_31022_, _31021_, _10605_);
  not (_31023_, _31022_);
  nor (_31025_, _31023_, _31020_);
  nor (_31026_, _31025_, _31019_);
  not (_31027_, _31026_);
  nor (_31028_, _31027_, _31018_);
  nor (_31029_, _31028_, _30885_);
  and (_31030_, _31029_, _30883_);
  nor (_31031_, _02679_, _30883_);
  or (_31032_, _31031_, _31030_);
  and (_31033_, _31032_, _10630_);
  not (_31034_, _30880_);
  nor (_31036_, _07587_, _01439_);
  and (_31037_, _30912_, _07587_);
  or (_31038_, _31037_, _31036_);
  and (_31039_, _31038_, _10629_);
  nor (_31040_, _31039_, _31034_);
  not (_31041_, _31040_);
  nor (_31042_, _31041_, _31033_);
  nor (_31043_, _31042_, _30881_);
  and (_31044_, _31043_, _30879_);
  nor (_31045_, _02679_, _30879_);
  or (_31047_, _31045_, _31044_);
  and (_31048_, _31047_, _10650_);
  and (_31049_, _06787_, \oc8051_golden_model_1.PC [0]);
  nor (_31050_, _06787_, \oc8051_golden_model_1.PC [0]);
  or (_31051_, _31050_, _10650_);
  or (_31052_, _31051_, _31049_);
  and (_31053_, _31052_, _30877_);
  not (_31054_, _31053_);
  nor (_31055_, _31054_, _31048_);
  nor (_31056_, _31055_, _30878_);
  and (_31058_, _31056_, _30876_);
  nor (_31059_, _02679_, _30876_);
  or (_31060_, _31059_, _31058_);
  and (_31061_, _31060_, _10123_);
  and (_31062_, _10120_, _07416_);
  not (_31063_, _31062_);
  or (_31064_, _31063_, _31061_);
  nor (_31065_, _31064_, _30875_);
  nor (_31066_, _31062_, _01439_);
  nor (_31067_, _31066_, _02350_);
  not (_31069_, _31067_);
  nor (_31070_, _31069_, _31065_);
  and (_31071_, _05120_, _02350_);
  or (_31072_, _31071_, _31070_);
  and (_31073_, _31072_, _04964_);
  nor (_31074_, _02679_, _04964_);
  or (_31075_, _31074_, _31073_);
  and (_31076_, _31075_, _10689_);
  not (_31077_, _30869_);
  and (_31078_, _30925_, _08690_);
  nor (_31080_, _08690_, _01439_);
  or (_31081_, _31080_, _10689_);
  nor (_31082_, _31081_, _31078_);
  nor (_31083_, _31082_, _31077_);
  not (_31084_, _31083_);
  nor (_31085_, _31084_, _31076_);
  nor (_31086_, _31085_, _30870_);
  and (_31087_, _31086_, _02084_);
  and (_31088_, _05120_, _02083_);
  or (_31089_, _31088_, _31087_);
  and (_31091_, _31089_, _10712_);
  nor (_31092_, _02679_, _10712_);
  nor (_31093_, _31092_, _31091_);
  nor (_31094_, _31093_, _02243_);
  not (_31095_, _30867_);
  and (_31096_, _08690_, \oc8051_golden_model_1.PC [0]);
  nor (_31097_, _30924_, _08690_);
  nor (_31098_, _31097_, _31096_);
  and (_31099_, _31098_, _02243_);
  nor (_31100_, _31099_, _31095_);
  not (_31102_, _31100_);
  nor (_31103_, _31102_, _31094_);
  nor (_31104_, _31103_, _30868_);
  nor (_31105_, _31104_, _03537_);
  and (_31106_, _03537_, _02679_);
  nor (_31107_, _31106_, _01697_);
  not (_31108_, _31107_);
  nor (_31109_, _31108_, _31105_);
  not (_31110_, _30865_);
  and (_31111_, _31098_, _01697_);
  nor (_31113_, _31111_, _31110_);
  not (_31114_, _31113_);
  nor (_31115_, _31114_, _31109_);
  nor (_31116_, _31115_, _30866_);
  nor (_31117_, _31116_, _30863_);
  or (_31118_, _31117_, _10762_);
  nor (_31119_, _31118_, _30864_);
  and (_31120_, _10762_, _01439_);
  nor (_31121_, _31120_, _31119_);
  nand (_31122_, _31121_, _39632_);
  or (_31123_, _39632_, \oc8051_golden_model_1.PC [0]);
  and (_31124_, _31123_, _39026_);
  and (_41793_, _31124_, _31122_);
  and (_31125_, _02366_, _01412_);
  nor (_31126_, _23257_, _03084_);
  nor (_31127_, _10133_, _10226_);
  nor (_31128_, _10139_, _10226_);
  nor (_31129_, _10147_, _10226_);
  nor (_31130_, _04919_, _01412_);
  and (_31131_, _08881_, _01805_);
  and (_31133_, _08770_, _01805_);
  nor (_31134_, _10230_, _10228_);
  nor (_31135_, _31134_, _10231_);
  not (_31136_, _31135_);
  nor (_31137_, _31136_, _08770_);
  or (_31138_, _31137_, _31133_);
  nor (_31139_, _31138_, _10471_);
  nor (_31140_, _10460_, _10226_);
  and (_31141_, _02079_, _01805_);
  or (_31142_, _10437_, _01412_);
  nor (_31144_, _10382_, _10380_);
  nor (_31145_, _31144_, _10383_);
  or (_31146_, _31145_, _10435_);
  and (_31147_, _31146_, _04535_);
  nand (_31148_, _31147_, _31142_);
  and (_31149_, _02893_, _10323_);
  nor (_31150_, _02560_, _02552_);
  nor (_31151_, _31150_, _10226_);
  and (_31152_, _02893_, _02060_);
  nor (_31153_, _30900_, _02062_);
  nor (_31155_, _31153_, _01412_);
  and (_31156_, _31153_, _01412_);
  nor (_31157_, _31156_, _31155_);
  nor (_31158_, _31157_, _02060_);
  nor (_31159_, _31158_, _06851_);
  not (_31160_, _31159_);
  nor (_31161_, _31160_, _31152_);
  not (_31162_, _31150_);
  and (_31163_, _06851_, _10226_);
  nor (_31164_, _31163_, _31162_);
  not (_31166_, _31164_);
  nor (_31167_, _31166_, _31161_);
  or (_31168_, _31167_, _02160_);
  nor (_31169_, _31168_, _31151_);
  and (_31170_, _02160_, _01412_);
  or (_31171_, _31170_, _06845_);
  or (_31172_, _31171_, _31169_);
  nand (_31173_, _06845_, _01805_);
  and (_31174_, _31173_, _31172_);
  nor (_31175_, _31174_, _10323_);
  or (_31177_, _31175_, _04535_);
  nor (_31178_, _31177_, _31149_);
  nor (_31179_, _31178_, _02079_);
  and (_31180_, _31179_, _31148_);
  or (_31181_, _31180_, _31141_);
  nand (_31182_, _31181_, _03006_);
  and (_31183_, _31135_, _10295_);
  and (_31184_, _10293_, _01805_);
  nor (_31185_, _31184_, _31183_);
  nand (_31186_, _31185_, _02158_);
  nand (_31188_, _31186_, _31182_);
  nand (_31189_, _31188_, _10287_);
  nor (_31190_, _10287_, _10226_);
  nor (_31191_, _31190_, _02057_);
  nand (_31192_, _31191_, _31189_);
  and (_31193_, _02057_, _01412_);
  nor (_31194_, _31193_, _03446_);
  nand (_31195_, _31194_, _31192_);
  and (_31196_, _02893_, _03446_);
  nor (_31197_, _31196_, _02155_);
  nand (_31199_, _31197_, _31195_);
  and (_31200_, _02155_, _01412_);
  nor (_31201_, _31200_, _22169_);
  nand (_31202_, _31201_, _31199_);
  nor (_31203_, _10452_, _10226_);
  nor (_31204_, _31203_, _02153_);
  nand (_31205_, _31204_, _31202_);
  and (_31206_, _02153_, _01412_);
  nor (_31207_, _31206_, _10462_);
  and (_31208_, _31207_, _31205_);
  or (_31210_, _31208_, _31140_);
  nand (_31211_, _31210_, _02054_);
  and (_31212_, _02053_, \oc8051_golden_model_1.PC [1]);
  nor (_31213_, _31212_, _10464_);
  and (_31214_, _31213_, _31211_);
  nor (_31215_, _02893_, _01757_);
  or (_31216_, _31215_, _31214_);
  nand (_31217_, _31216_, _03114_);
  and (_31218_, _02052_, _01412_);
  nor (_31219_, _31218_, _10475_);
  and (_31221_, _31219_, _31217_);
  or (_31222_, _31221_, _31139_);
  nand (_31223_, _31222_, _08836_);
  or (_31224_, _31136_, _08842_);
  or (_31225_, _10482_, _10226_);
  and (_31226_, _31225_, _08790_);
  nand (_31227_, _31226_, _31224_);
  nand (_31228_, _31227_, _31223_);
  nand (_31229_, _31228_, _02547_);
  nor (_31230_, _31136_, _08877_);
  not (_31232_, _31230_);
  and (_31233_, _08877_, _01805_);
  nor (_31234_, _31233_, _02547_);
  and (_31235_, _31234_, _31232_);
  nor (_31236_, _31235_, _02246_);
  nand (_31237_, _31236_, _31229_);
  nor (_31238_, _31135_, _08922_);
  and (_31239_, _08922_, _10226_);
  or (_31240_, _31239_, _08917_);
  or (_31241_, _31240_, _31238_);
  and (_31243_, _31241_, _08882_);
  and (_31244_, _31243_, _31237_);
  or (_31245_, _31244_, _31131_);
  nand (_31246_, _31245_, _02047_);
  and (_31247_, _02046_, \oc8051_golden_model_1.PC [1]);
  nor (_31248_, _31247_, _03310_);
  nand (_31249_, _31248_, _31246_);
  nor (_31250_, _02893_, _01750_);
  not (_31251_, _02147_);
  not (_31252_, _22232_);
  and (_31254_, _31252_, _22229_);
  and (_31255_, _31254_, _31251_);
  not (_31256_, _31255_);
  nor (_31257_, _31256_, _31250_);
  nand (_31258_, _31257_, _31249_);
  nor (_31259_, _31255_, _01412_);
  nor (_31260_, _31259_, _10155_);
  nand (_31261_, _31260_, _31258_);
  and (_31262_, _10157_, _01805_);
  or (_31263_, _31262_, _10158_);
  nand (_31265_, _31263_, _31261_);
  nor (_31266_, _10157_, _10226_);
  nor (_31267_, _31266_, _02182_);
  nand (_31268_, _31267_, _31265_);
  and (_31269_, _02182_, _01412_);
  nor (_31270_, _31269_, _10513_);
  nand (_31271_, _31270_, _31268_);
  and (_31272_, _02893_, _10513_);
  nor (_31273_, _31272_, _02181_);
  and (_31274_, _31273_, _31271_);
  and (_31276_, _02181_, _01412_);
  or (_31277_, _31276_, _31274_);
  nand (_31278_, _31277_, _09041_);
  nor (_31279_, _04916_, _01777_);
  nor (_31280_, _09041_, _01805_);
  nor (_31281_, _31280_, _31279_);
  nand (_31282_, _31281_, _31278_);
  and (_31283_, _31279_, _01805_);
  nor (_31284_, _31283_, _02623_);
  nand (_31285_, _31284_, _31282_);
  and (_31286_, _02623_, _10226_);
  nor (_31287_, _31286_, _07017_);
  nand (_31288_, _31287_, _31285_);
  nor (_31289_, _07016_, _01412_);
  nor (_31290_, _31289_, _01876_);
  nand (_31291_, _31290_, _31288_);
  nor (_31292_, _01805_, _01778_);
  nor (_31293_, _31292_, _02042_);
  and (_31294_, _31293_, _31291_);
  and (_31295_, _02042_, \oc8051_golden_model_1.PC [1]);
  or (_31297_, _31295_, _31294_);
  nand (_31298_, _31297_, _04460_);
  and (_31299_, _02893_, _01767_);
  nor (_31300_, _31299_, _02218_);
  nand (_31301_, _31300_, _31298_);
  and (_31302_, _02218_, _01805_);
  not (_31303_, _31302_);
  and (_31304_, _31303_, _10534_);
  nand (_31305_, _31304_, _31301_);
  nor (_31306_, _10534_, _01412_);
  nor (_31308_, _31306_, _01765_);
  nand (_31309_, _31308_, _31305_);
  and (_31310_, _01805_, _01765_);
  nor (_31311_, _31310_, _10546_);
  nand (_31312_, _31311_, _31309_);
  nor (_31313_, _10542_, _10226_);
  nor (_31314_, _31313_, _02124_);
  nand (_31315_, _31314_, _31312_);
  and (_31316_, _02124_, _01412_);
  nor (_31317_, _31316_, _01711_);
  nand (_31319_, _31317_, _31315_);
  and (_31320_, _02893_, _01711_);
  nor (_31321_, _31320_, _10550_);
  nand (_31322_, _31321_, _31319_);
  and (_31323_, _31145_, _10550_);
  nor (_31324_, _31323_, _04920_);
  and (_31325_, _31324_, _31322_);
  or (_31326_, _31325_, _31130_);
  nand (_31327_, _31326_, _01995_);
  and (_31328_, _01994_, _10226_);
  nor (_31330_, _31328_, _07239_);
  nand (_31331_, _31330_, _31327_);
  and (_31332_, _07239_, _01412_);
  nor (_31333_, _31332_, _10149_);
  nand (_31334_, _31333_, _31331_);
  and (_31335_, _10149_, _01863_);
  nor (_31336_, _31335_, _02123_);
  nand (_31337_, _31336_, _31334_);
  and (_31338_, _02123_, _01412_);
  nor (_31339_, _31338_, _01718_);
  nand (_31341_, _31339_, _31337_);
  and (_31342_, _02893_, _01718_);
  nor (_31343_, _31342_, _10604_);
  nand (_31344_, _31343_, _31341_);
  nor (_31345_, _31145_, _07587_);
  and (_31346_, _07587_, \oc8051_golden_model_1.PC [1]);
  nor (_31347_, _31346_, _10605_);
  not (_31348_, _31347_);
  nor (_31349_, _31348_, _31345_);
  nor (_31350_, _31349_, _10609_);
  and (_31352_, _31350_, _31344_);
  or (_31353_, _31352_, _31129_);
  nand (_31354_, _31353_, _10618_);
  nor (_31355_, _10618_, _01412_);
  nor (_31356_, _31355_, _02210_);
  nand (_31357_, _31356_, _31354_);
  and (_31358_, _02210_, _01805_);
  nor (_31359_, _31358_, _02331_);
  and (_31360_, _31359_, _31357_);
  and (_31361_, _02331_, \oc8051_golden_model_1.PC [1]);
  or (_31363_, _31361_, _31360_);
  nand (_31364_, _31363_, _30883_);
  and (_31365_, _02893_, _01722_);
  nor (_31366_, _31365_, _10629_);
  nand (_31367_, _31366_, _31364_);
  nor (_31368_, _07587_, \oc8051_golden_model_1.PC [1]);
  and (_31369_, _31145_, _07587_);
  or (_31370_, _31369_, _31368_);
  and (_31371_, _31370_, _10629_);
  nor (_31372_, _31371_, _10634_);
  and (_31374_, _31372_, _31367_);
  or (_31375_, _31374_, _31128_);
  nand (_31376_, _31375_, _10135_);
  nor (_31377_, _10135_, _01412_);
  nor (_31378_, _31377_, _02206_);
  nand (_31379_, _31378_, _31376_);
  and (_31380_, _02206_, _01805_);
  nor (_31381_, _31380_, _02342_);
  and (_31382_, _31381_, _31379_);
  and (_31383_, _02342_, \oc8051_golden_model_1.PC [1]);
  or (_31385_, _31383_, _31382_);
  nand (_31386_, _31385_, _30879_);
  and (_31387_, _02893_, _01728_);
  nor (_31388_, _31387_, _10649_);
  nand (_31389_, _31388_, _31386_);
  nor (_31390_, _31145_, \oc8051_golden_model_1.PSW [7]);
  and (_31391_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  nor (_31392_, _31391_, _10650_);
  not (_31393_, _31392_);
  nor (_31394_, _31393_, _31390_);
  nor (_31396_, _31394_, _10654_);
  and (_31397_, _31396_, _31389_);
  or (_31398_, _31397_, _31127_);
  nand (_31399_, _31398_, _07339_);
  nor (_31400_, _07339_, _01412_);
  nor (_31401_, _31400_, _02202_);
  and (_31402_, _31401_, _31399_);
  and (_31403_, _02202_, _01805_);
  or (_31404_, _31403_, _02334_);
  nor (_31405_, _31404_, _31402_);
  and (_31407_, _02334_, \oc8051_golden_model_1.PC [1]);
  or (_31408_, _31407_, _31405_);
  nand (_31409_, _31408_, _30876_);
  and (_31410_, _02893_, _01736_);
  nor (_31411_, _31410_, _10122_);
  and (_31412_, _31411_, _31409_);
  nor (_31413_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_31414_, _31145_, \oc8051_golden_model_1.PSW [7]);
  or (_31415_, _31414_, _31413_);
  and (_31416_, _31415_, _10122_);
  or (_31418_, _31416_, _31412_);
  nand (_31419_, _31418_, _10120_);
  nor (_31420_, _10120_, _01805_);
  nor (_31421_, _31420_, _07386_);
  nand (_31422_, _31421_, _31419_);
  nor (_31423_, _07385_, _01412_);
  nor (_31424_, _31423_, _07415_);
  nand (_31425_, _31424_, _31422_);
  and (_31426_, _07415_, _10226_);
  nor (_31427_, _31426_, _02350_);
  and (_31429_, _31427_, _31425_);
  nor (_31430_, _05075_, _09472_);
  or (_31431_, _31430_, _31429_);
  nand (_31432_, _31431_, _04964_);
  and (_31433_, _02893_, _01726_);
  nor (_31434_, _31433_, _02200_);
  and (_31435_, _31434_, _31432_);
  nor (_31436_, _08690_, _10226_);
  and (_31437_, _31135_, _08690_);
  nor (_31438_, _31437_, _31436_);
  nor (_31440_, _31438_, _10689_);
  or (_31441_, _31440_, _31435_);
  nand (_31442_, _31441_, _10118_);
  nor (_31443_, _10118_, _01805_);
  nor (_31444_, _31443_, _07489_);
  nand (_31445_, _31444_, _31442_);
  nor (_31446_, _07488_, _01412_);
  nor (_31447_, _31446_, _07533_);
  nand (_31448_, _31447_, _31445_);
  and (_31449_, _07533_, _10226_);
  nor (_31450_, _31449_, _02083_);
  and (_31451_, _31450_, _31448_);
  nor (_31452_, _05075_, _02084_);
  or (_31453_, _31452_, _31451_);
  nand (_31454_, _31453_, _10712_);
  and (_31455_, _02893_, _01738_);
  nor (_31456_, _31455_, _02243_);
  nand (_31457_, _31456_, _31454_);
  nor (_31458_, _31135_, _08690_);
  and (_31459_, _08690_, _10226_);
  nor (_31461_, _31459_, _31458_);
  and (_31462_, _31461_, _02243_);
  nor (_31463_, _23255_, _04970_);
  not (_31464_, _31463_);
  nor (_31465_, _31464_, _31462_);
  and (_31466_, _31465_, _31457_);
  nor (_31467_, _31463_, _10226_);
  or (_31468_, _31467_, _31466_);
  nand (_31469_, _31468_, _31126_);
  nor (_31470_, _31126_, _10226_);
  nor (_31472_, _31470_, _02366_);
  and (_31473_, _31472_, _31469_);
  or (_31474_, _31473_, _31125_);
  nand (_31475_, _31474_, _07581_);
  nor (_31476_, _07581_, _01805_);
  nor (_31477_, _31476_, _03537_);
  nand (_31478_, _31477_, _31475_);
  and (_31479_, _03537_, _02893_);
  nor (_31480_, _31479_, _01697_);
  nand (_31481_, _31480_, _31478_);
  and (_31483_, _31461_, _01697_);
  nor (_31484_, _31483_, _05338_);
  and (_31485_, _31484_, _31481_);
  nor (_31486_, _05337_, _10226_);
  or (_31487_, _31486_, _31485_);
  nand (_31488_, _31487_, _03326_);
  and (_31489_, _02222_, _01731_);
  nor (_31490_, _31489_, _01805_);
  or (_31491_, _31490_, _23298_);
  nand (_31492_, _31491_, _31488_);
  nand (_31494_, _02786_, _10226_);
  nand (_31495_, _31494_, _31492_);
  nand (_31496_, _31495_, _02082_);
  not (_31497_, _10751_);
  and (_31498_, _02081_, _01412_);
  nor (_31499_, _31498_, _31497_);
  and (_31500_, _31499_, _31496_);
  nor (_31501_, _10751_, _10226_);
  or (_31502_, _31501_, _31500_);
  nand (_31503_, _31502_, _23330_);
  and (_31505_, _30863_, _02893_);
  nor (_31506_, _31505_, _10762_);
  nand (_31507_, _31506_, _31503_);
  and (_31508_, _10762_, _10226_);
  not (_31509_, _31508_);
  nand (_31510_, _31509_, _31507_);
  or (_31511_, _31510_, _39633_);
  or (_31512_, _39632_, \oc8051_golden_model_1.PC [1]);
  and (_31513_, _31512_, _39026_);
  and (_41794_, _31513_, _31511_);
  and (_31515_, _02081_, _01701_);
  nor (_31516_, _10118_, _01782_);
  nor (_31517_, _10120_, _01782_);
  nor (_31518_, _10133_, _01782_);
  nor (_31519_, _10139_, _01782_);
  nor (_31520_, _10147_, _01782_);
  not (_31521_, _02124_);
  nor (_31522_, _10542_, _01782_);
  nor (_31523_, _10153_, _01782_);
  nor (_31524_, _31255_, _01701_);
  and (_31526_, _08881_, _01783_);
  and (_31527_, _10235_, _10232_);
  nor (_31528_, _31527_, _10236_);
  and (_31529_, _31528_, _10482_);
  and (_31530_, _10223_, _08842_);
  nor (_31531_, _31530_, _31529_);
  nor (_31532_, _31531_, _08836_);
  not (_31533_, _31528_);
  and (_31534_, _31533_, _10295_);
  and (_31535_, _10293_, _10224_);
  nor (_31537_, _31535_, _31534_);
  or (_31538_, _31537_, _03006_);
  and (_31539_, _10435_, _01701_);
  and (_31540_, _10387_, _10384_);
  nor (_31541_, _31540_, _10388_);
  and (_31542_, _31541_, _10437_);
  nor (_31543_, _31542_, _31539_);
  nand (_31544_, _31543_, _04535_);
  nor (_31545_, _10312_, _01782_);
  not (_31546_, _31545_);
  and (_31548_, _02062_, _01702_);
  nor (_31549_, _02062_, \oc8051_golden_model_1.PC [2]);
  and (_31550_, _31549_, _10302_);
  nor (_31551_, _31550_, _31548_);
  nor (_31552_, _31551_, _06855_);
  nor (_31553_, _31552_, _02060_);
  and (_31554_, _31553_, _31546_);
  not (_31555_, _06859_);
  nor (_31556_, _02494_, _01747_);
  or (_31557_, _31556_, _31555_);
  nor (_31559_, _31557_, _31554_);
  nor (_31560_, _06859_, _01782_);
  nor (_31561_, _31560_, _02160_);
  not (_31562_, _31561_);
  nor (_31563_, _31562_, _31559_);
  and (_31564_, _02160_, _01701_);
  or (_31565_, _31564_, _31563_);
  and (_31566_, _31565_, _10299_);
  and (_31567_, _06845_, _01782_);
  or (_31568_, _31567_, _31566_);
  and (_31570_, _31568_, _01752_);
  nor (_31571_, _02494_, _01752_);
  nor (_31572_, _31571_, _04535_);
  not (_31573_, _31572_);
  nor (_31574_, _31573_, _31570_);
  nor (_31575_, _31574_, _02079_);
  and (_31576_, _31575_, _31544_);
  and (_31577_, _02079_, _01782_);
  or (_31578_, _31577_, _02158_);
  or (_31579_, _31578_, _31576_);
  nand (_31581_, _31579_, _31538_);
  nand (_31582_, _31581_, _10287_);
  nor (_31583_, _10287_, _01782_);
  nor (_31584_, _31583_, _02057_);
  nand (_31585_, _31584_, _31582_);
  and (_31586_, _02057_, _01701_);
  nor (_31587_, _31586_, _03446_);
  nand (_31588_, _31587_, _31585_);
  and (_31589_, _02494_, _03446_);
  nor (_31590_, _31589_, _02155_);
  nand (_31592_, _31590_, _31588_);
  and (_31593_, _02155_, _01701_);
  nor (_31594_, _31593_, _22169_);
  nand (_31595_, _31594_, _31592_);
  nor (_31596_, _10452_, _01782_);
  nor (_31597_, _31596_, _02153_);
  nand (_31598_, _31597_, _31595_);
  and (_31599_, _02153_, _01701_);
  nor (_31600_, _31599_, _10462_);
  nand (_31601_, _31600_, _31598_);
  nor (_31603_, _10460_, _01782_);
  nor (_31604_, _31603_, _02053_);
  nand (_31605_, _31604_, _31601_);
  and (_31606_, _02053_, _01701_);
  nor (_31607_, _31606_, _10464_);
  nand (_31608_, _31607_, _31605_);
  and (_31609_, _02494_, _10464_);
  nor (_31610_, _31609_, _02052_);
  nand (_31611_, _31610_, _31608_);
  and (_31612_, _02052_, _01701_);
  nor (_31613_, _31612_, _10475_);
  nand (_31614_, _31613_, _31611_);
  and (_31615_, _10223_, _08770_);
  nor (_31616_, _31533_, _08770_);
  or (_31617_, _31616_, _31615_);
  nor (_31618_, _31617_, _10471_);
  nor (_31619_, _31618_, _08790_);
  nand (_31620_, _31619_, _31614_);
  nand (_31621_, _31620_, _02547_);
  or (_31622_, _31621_, _31532_);
  nor (_31624_, _31533_, _08877_);
  not (_31625_, _31624_);
  and (_31626_, _10223_, _08877_);
  nor (_31627_, _31626_, _02547_);
  and (_31628_, _31627_, _31625_);
  nor (_31629_, _31628_, _02246_);
  nand (_31630_, _31629_, _31622_);
  nor (_31631_, _31528_, _08922_);
  and (_31632_, _10224_, _08922_);
  or (_31633_, _31632_, _08917_);
  nor (_31635_, _31633_, _31631_);
  nor (_31636_, _31635_, _08881_);
  and (_31637_, _31636_, _31630_);
  or (_31638_, _31637_, _31526_);
  nand (_31639_, _31638_, _02047_);
  and (_31640_, _02046_, _01702_);
  nor (_31641_, _31640_, _03310_);
  nand (_31642_, _31641_, _31639_);
  nor (_31643_, _02494_, _01750_);
  nor (_31644_, _31643_, _31256_);
  and (_31646_, _31644_, _31642_);
  or (_31647_, _31646_, _31524_);
  nand (_31648_, _31647_, _10158_);
  nor (_31649_, _10158_, _01782_);
  nor (_31650_, _31649_, _02182_);
  nand (_31651_, _31650_, _31648_);
  and (_31652_, _02182_, _01701_);
  nor (_31653_, _31652_, _10513_);
  nand (_31654_, _31653_, _31651_);
  and (_31655_, _02494_, _10513_);
  nor (_31657_, _31655_, _02181_);
  nand (_31658_, _31657_, _31654_);
  and (_31659_, _02181_, _01701_);
  nor (_31660_, _31659_, _10517_);
  and (_31661_, _31660_, _31658_);
  or (_31662_, _31661_, _31523_);
  nand (_31663_, _31662_, _07016_);
  nor (_31664_, _07016_, _01701_);
  nor (_31665_, _31664_, _01876_);
  nand (_31666_, _31665_, _31663_);
  nor (_31668_, _01783_, _01778_);
  nor (_31669_, _31668_, _02042_);
  and (_31670_, _31669_, _31666_);
  and (_31671_, _02042_, _01702_);
  or (_31672_, _31671_, _31670_);
  nand (_31673_, _31672_, _04460_);
  and (_31674_, _02494_, _01767_);
  nor (_31675_, _31674_, _02218_);
  nand (_31676_, _31675_, _31673_);
  nor (_31677_, _05443_, _02031_);
  and (_31679_, _02644_, _01701_);
  and (_31680_, _10223_, _02218_);
  nor (_31681_, _31680_, _31679_);
  and (_31682_, _31681_, _31677_);
  nand (_31683_, _31682_, _31676_);
  nor (_31684_, _10534_, _01701_);
  nor (_31685_, _31684_, _01765_);
  nand (_31686_, _31685_, _31683_);
  and (_31687_, _10223_, _01765_);
  nor (_31688_, _31687_, _10546_);
  and (_31690_, _31688_, _31686_);
  or (_31691_, _31690_, _31522_);
  nand (_31692_, _31691_, _31521_);
  and (_31693_, _02124_, _01702_);
  nor (_31694_, _31693_, _01711_);
  nand (_31695_, _31694_, _31692_);
  nor (_31696_, _02494_, _01712_);
  nor (_31697_, _31696_, _10550_);
  nand (_31698_, _31697_, _31695_);
  nor (_31699_, _31541_, _10551_);
  nor (_31701_, _31699_, _03344_);
  nand (_31702_, _31701_, _31698_);
  and (_31703_, _03344_, _01701_);
  and (_31704_, _02130_, _01717_);
  nor (_31705_, _31704_, _04915_);
  not (_31706_, _31705_);
  nor (_31707_, _31706_, _31703_);
  nand (_31708_, _31707_, _31702_);
  and (_31709_, _02133_, _01717_);
  nor (_31710_, _31705_, _01701_);
  nor (_31712_, _31710_, _31709_);
  nand (_31713_, _31712_, _31708_);
  and (_31714_, _31709_, _01701_);
  nor (_31715_, _31714_, _22538_);
  nand (_31716_, _31715_, _31713_);
  and (_31717_, _22538_, _01702_);
  nor (_31718_, _31717_, _01994_);
  nand (_31719_, _31718_, _31716_);
  and (_31720_, _10223_, _01994_);
  nor (_31721_, _31720_, _07239_);
  and (_31723_, _31721_, _31719_);
  and (_31724_, _07239_, _01702_);
  or (_31725_, _31724_, _31723_);
  nand (_31726_, _31725_, _10150_);
  nor (_31727_, _10150_, _01798_);
  nor (_31728_, _31727_, _02123_);
  nand (_31729_, _31728_, _31726_);
  and (_31730_, _02123_, _01701_);
  nor (_31731_, _31730_, _01718_);
  nand (_31732_, _31731_, _31729_);
  and (_31734_, _02494_, _01718_);
  nor (_31735_, _31734_, _10604_);
  nand (_31736_, _31735_, _31732_);
  nor (_31737_, _31541_, _07587_);
  and (_31738_, _07587_, _01702_);
  nor (_31739_, _31738_, _10605_);
  not (_31740_, _31739_);
  nor (_31741_, _31740_, _31737_);
  nor (_31742_, _31741_, _10609_);
  and (_31743_, _31742_, _31736_);
  or (_31745_, _31743_, _31520_);
  nand (_31746_, _31745_, _10618_);
  nor (_31747_, _10618_, _01701_);
  nor (_31748_, _31747_, _02210_);
  nand (_31749_, _31748_, _31746_);
  and (_31750_, _10223_, _02210_);
  nor (_31751_, _31750_, _02331_);
  and (_31752_, _31751_, _31749_);
  and (_31753_, _02331_, _01702_);
  or (_31754_, _31753_, _31752_);
  nand (_31756_, _31754_, _30883_);
  and (_31757_, _02494_, _01722_);
  nor (_31758_, _31757_, _10629_);
  nand (_31759_, _31758_, _31756_);
  nor (_31760_, _07587_, _01702_);
  and (_31761_, _31541_, _07587_);
  or (_31762_, _31761_, _31760_);
  and (_31763_, _31762_, _10629_);
  nor (_31764_, _31763_, _10634_);
  and (_31765_, _31764_, _31759_);
  or (_31767_, _31765_, _31519_);
  nand (_31768_, _31767_, _10135_);
  nor (_31769_, _10135_, _01701_);
  nor (_31770_, _31769_, _02206_);
  nand (_31771_, _31770_, _31768_);
  and (_31772_, _10223_, _02206_);
  nor (_31773_, _31772_, _02342_);
  and (_31774_, _31773_, _31771_);
  and (_31775_, _02342_, _01702_);
  or (_31776_, _31775_, _31774_);
  nand (_31777_, _31776_, _30879_);
  and (_31778_, _02494_, _01728_);
  nor (_31779_, _31778_, _10649_);
  nand (_31780_, _31779_, _31777_);
  or (_31781_, _31541_, \oc8051_golden_model_1.PSW [7]);
  or (_31782_, _01701_, _06707_);
  and (_31783_, _31782_, _10649_);
  and (_31784_, _31783_, _31781_);
  nor (_31785_, _31784_, _10654_);
  and (_31786_, _31785_, _31780_);
  or (_31788_, _31786_, _31518_);
  nand (_31789_, _31788_, _07339_);
  nor (_31790_, _07339_, _01701_);
  nor (_31791_, _31790_, _02202_);
  nand (_31792_, _31791_, _31789_);
  and (_31793_, _10223_, _02202_);
  nor (_31794_, _31793_, _02334_);
  and (_31795_, _31794_, _31792_);
  and (_31796_, _02334_, _01702_);
  or (_31797_, _31796_, _31795_);
  nand (_31799_, _31797_, _30876_);
  and (_31800_, _02494_, _01736_);
  nor (_31801_, _31800_, _10122_);
  nand (_31802_, _31801_, _31799_);
  nor (_31803_, _31541_, _06707_);
  nor (_31804_, _01701_, \oc8051_golden_model_1.PSW [7]);
  nor (_31805_, _31804_, _10123_);
  not (_31806_, _31805_);
  nor (_31807_, _31806_, _31803_);
  nor (_31808_, _31807_, _10671_);
  and (_31810_, _31808_, _31802_);
  or (_31811_, _31810_, _31517_);
  nand (_31812_, _31811_, _07385_);
  nor (_31813_, _07385_, _01701_);
  nor (_31814_, _31813_, _07415_);
  nand (_31815_, _31814_, _31812_);
  and (_31816_, _07415_, _01782_);
  nor (_31817_, _31816_, _02350_);
  and (_31818_, _31817_, _31815_);
  nor (_31819_, _05211_, _09472_);
  or (_31821_, _31819_, _31818_);
  nand (_31822_, _31821_, _04964_);
  and (_31823_, _02494_, _01726_);
  nor (_31824_, _31823_, _02200_);
  nand (_31825_, _31824_, _31822_);
  and (_31826_, _31533_, _08690_);
  nor (_31827_, _10223_, _08690_);
  or (_31828_, _31827_, _10689_);
  nor (_31829_, _31828_, _31826_);
  nor (_31830_, _31829_, _10693_);
  and (_31832_, _31830_, _31825_);
  or (_31833_, _31832_, _31516_);
  nand (_31834_, _31833_, _07488_);
  nor (_31835_, _07488_, _01701_);
  nor (_31836_, _31835_, _07533_);
  nand (_31837_, _31836_, _31834_);
  and (_31838_, _07533_, _01782_);
  nor (_31839_, _31838_, _02083_);
  and (_31840_, _31839_, _31837_);
  nor (_31841_, _05211_, _02084_);
  or (_31843_, _31841_, _31840_);
  nand (_31844_, _31843_, _10712_);
  and (_31845_, _02494_, _01738_);
  nor (_31846_, _31845_, _02243_);
  nand (_31847_, _31846_, _31844_);
  nor (_31848_, _31528_, _08690_);
  and (_31849_, _10224_, _08690_);
  nor (_31850_, _31849_, _31848_);
  and (_31851_, _31850_, _02243_);
  nor (_31852_, _31851_, _10723_);
  nand (_31854_, _31852_, _31847_);
  nor (_31855_, _10722_, _01782_);
  nor (_31856_, _31855_, _02366_);
  nand (_31857_, _31856_, _31854_);
  not (_31858_, _07581_);
  and (_31859_, _02366_, _01701_);
  nor (_31860_, _31859_, _31858_);
  and (_31861_, _31860_, _31857_);
  nor (_31862_, _07581_, _01782_);
  or (_31863_, _31862_, _31861_);
  nand (_31865_, _31863_, _01990_);
  and (_31866_, _03537_, _02494_);
  nor (_31867_, _31866_, _01697_);
  nand (_31868_, _31867_, _31865_);
  and (_31869_, _31850_, _01697_);
  nor (_31870_, _31869_, _10744_);
  nand (_31871_, _31870_, _31868_);
  and (_31872_, _10744_, _01783_);
  nor (_31873_, _31872_, _02081_);
  and (_31874_, _31873_, _31871_);
  or (_31876_, _31874_, _31515_);
  nand (_31877_, _31876_, _10751_);
  nor (_31878_, _10751_, _01783_);
  nor (_31879_, _31878_, _30863_);
  nand (_31880_, _31879_, _31877_);
  and (_31881_, _30863_, _02494_);
  nor (_31882_, _31881_, _10762_);
  nand (_31883_, _31882_, _31880_);
  and (_31884_, _10762_, _01782_);
  not (_31885_, _31884_);
  and (_31887_, _31885_, _31883_);
  nand (_31888_, _31887_, _39632_);
  or (_31889_, _39632_, \oc8051_golden_model_1.PC [2]);
  and (_31890_, _31889_, _39026_);
  and (_41795_, _31890_, _31888_);
  and (_31891_, _02081_, _01825_);
  and (_31892_, _02366_, _01825_);
  nor (_31893_, _10118_, _02266_);
  nor (_31894_, _10120_, _02266_);
  nor (_31895_, _10133_, _02266_);
  nor (_31897_, _10139_, _02266_);
  nor (_31898_, _10147_, _02266_);
  nor (_31899_, _04919_, _01825_);
  and (_31900_, _10218_, _02218_);
  nor (_31901_, _31255_, _01825_);
  or (_31902_, _10295_, _10218_);
  or (_31903_, _10221_, _10220_);
  and (_31904_, _31903_, _10237_);
  nor (_31905_, _31903_, _10237_);
  nor (_31906_, _31905_, _31904_);
  or (_31908_, _31906_, _10293_);
  and (_31909_, _31908_, _31902_);
  or (_31910_, _31909_, _03006_);
  and (_31911_, _10435_, _01825_);
  or (_31912_, _10377_, _10376_);
  and (_31913_, _31912_, _10389_);
  nor (_31914_, _31912_, _10389_);
  nor (_31915_, _31914_, _31913_);
  and (_31916_, _31915_, _10437_);
  nor (_31917_, _31916_, _31911_);
  nand (_31919_, _31917_, _04535_);
  nor (_31920_, _10301_, \oc8051_golden_model_1.PC [3]);
  nor (_31921_, _31920_, _02062_);
  and (_31922_, _02062_, _01825_);
  nor (_31923_, _31922_, _06855_);
  not (_31924_, _31923_);
  nor (_31925_, _31924_, _31921_);
  not (_31926_, _31925_);
  nor (_31927_, _10312_, _02266_);
  nor (_31928_, _31927_, _02060_);
  and (_31930_, _31928_, _31926_);
  nor (_31931_, _02324_, _01747_);
  or (_31932_, _31931_, _31555_);
  nor (_31933_, _31932_, _31930_);
  nor (_31934_, _06859_, _02266_);
  nor (_31935_, _31934_, _02160_);
  not (_31936_, _31935_);
  nor (_31937_, _31936_, _31933_);
  and (_31938_, _02160_, _01825_);
  or (_31939_, _31938_, _31937_);
  and (_31940_, _31939_, _10299_);
  and (_31941_, _06845_, _02266_);
  or (_31942_, _31941_, _31940_);
  and (_31943_, _31942_, _01752_);
  nor (_31944_, _02324_, _01752_);
  or (_31945_, _31944_, _04535_);
  nor (_31946_, _31945_, _31943_);
  nor (_31947_, _31946_, _02079_);
  and (_31948_, _31947_, _31919_);
  and (_31949_, _02079_, _02266_);
  or (_31951_, _31949_, _02158_);
  or (_31952_, _31951_, _31948_);
  nand (_31953_, _31952_, _31910_);
  nand (_31954_, _31953_, _10287_);
  nor (_31955_, _10287_, _02266_);
  nor (_31956_, _31955_, _02057_);
  nand (_31957_, _31956_, _31954_);
  and (_31958_, _02057_, _01825_);
  nor (_31959_, _31958_, _03446_);
  nand (_31960_, _31959_, _31957_);
  and (_31962_, _02324_, _03446_);
  nor (_31963_, _31962_, _02155_);
  nand (_31964_, _31963_, _31960_);
  and (_31965_, _02155_, _01825_);
  nor (_31966_, _31965_, _22169_);
  nand (_31967_, _31966_, _31964_);
  nor (_31968_, _10452_, _02266_);
  nor (_31969_, _31968_, _02153_);
  nand (_31970_, _31969_, _31967_);
  and (_31971_, _02153_, _01825_);
  nor (_31973_, _31971_, _10462_);
  nand (_31974_, _31973_, _31970_);
  nor (_31975_, _10460_, _02266_);
  nor (_31976_, _31975_, _02053_);
  nand (_31977_, _31976_, _31974_);
  and (_31978_, _02053_, _01825_);
  nor (_31979_, _31978_, _10464_);
  nand (_31980_, _31979_, _31977_);
  and (_31981_, _02324_, _10464_);
  nor (_31982_, _31981_, _02052_);
  nand (_31984_, _31982_, _31980_);
  and (_31985_, _02052_, _01825_);
  nor (_31986_, _31985_, _10475_);
  nand (_31987_, _31986_, _31984_);
  and (_31988_, _10218_, _08770_);
  not (_31989_, _31906_);
  nor (_31990_, _31989_, _08770_);
  or (_31991_, _31990_, _31988_);
  nor (_31992_, _31991_, _10471_);
  nor (_31993_, _31992_, _08790_);
  nand (_31995_, _31993_, _31987_);
  or (_31996_, _31989_, _08842_);
  or (_31997_, _10219_, _10482_);
  nand (_31998_, _31997_, _31996_);
  nand (_31999_, _31998_, _08790_);
  and (_32000_, _31999_, _02547_);
  nand (_32001_, _32000_, _31995_);
  nor (_32002_, _31989_, _08877_);
  not (_32003_, _32002_);
  and (_32004_, _10218_, _08877_);
  nor (_32006_, _32004_, _02547_);
  and (_32007_, _32006_, _32003_);
  nor (_32008_, _32007_, _02246_);
  nand (_32009_, _32008_, _32001_);
  nand (_32010_, _10218_, _08922_);
  not (_32011_, _08922_);
  nand (_32012_, _31906_, _32011_);
  and (_32013_, _32012_, _32010_);
  or (_32014_, _32013_, _08917_);
  and (_32015_, _32014_, _32009_);
  or (_32017_, _32015_, _08881_);
  nand (_32018_, _08881_, _02266_);
  and (_32019_, _32018_, _32017_);
  nand (_32020_, _32019_, _02047_);
  and (_32021_, _02046_, _02264_);
  nor (_32022_, _32021_, _03310_);
  nand (_32023_, _32022_, _32020_);
  nor (_32024_, _02324_, _01750_);
  nor (_32025_, _32024_, _31256_);
  and (_32026_, _32025_, _32023_);
  or (_32028_, _32026_, _31901_);
  nand (_32029_, _32028_, _10158_);
  nor (_32030_, _10158_, _02266_);
  nor (_32031_, _32030_, _02182_);
  nand (_32032_, _32031_, _32029_);
  and (_32033_, _02182_, _01825_);
  nor (_32034_, _32033_, _10513_);
  nand (_32035_, _32034_, _32032_);
  and (_32036_, _02324_, _10513_);
  nor (_32037_, _32036_, _02181_);
  nand (_32039_, _32037_, _32035_);
  and (_32040_, _02181_, _01825_);
  nor (_32041_, _32040_, _10517_);
  and (_32042_, _32041_, _32039_);
  nor (_32043_, _10153_, _02266_);
  or (_32044_, _32043_, _32042_);
  nand (_32045_, _32044_, _07016_);
  nor (_32046_, _07016_, _01825_);
  nor (_32047_, _32046_, _01876_);
  and (_32048_, _32047_, _32045_);
  nor (_32050_, _01778_, _01830_);
  or (_32051_, _32050_, _02042_);
  nor (_32052_, _32051_, _32048_);
  and (_32053_, _02042_, _02264_);
  or (_32054_, _32053_, _32052_);
  nand (_32055_, _32054_, _04460_);
  and (_32056_, _02324_, _01767_);
  nor (_32057_, _32056_, _02218_);
  nand (_32058_, _32057_, _32055_);
  nand (_32059_, _32058_, _10534_);
  or (_32061_, _32059_, _31900_);
  nor (_32062_, _10534_, _01825_);
  nor (_32063_, _32062_, _01765_);
  nand (_32064_, _32063_, _32061_);
  and (_32065_, _10218_, _01765_);
  nor (_32066_, _32065_, _10546_);
  nand (_32067_, _32066_, _32064_);
  nor (_32068_, _10542_, _02266_);
  nor (_32069_, _32068_, _02124_);
  nand (_32070_, _32069_, _32067_);
  and (_32072_, _02124_, _01825_);
  nor (_32073_, _32072_, _01711_);
  nand (_32074_, _32073_, _32070_);
  and (_32075_, _02324_, _01711_);
  nor (_32076_, _32075_, _10550_);
  nand (_32077_, _32076_, _32074_);
  and (_32078_, _31915_, _10550_);
  nor (_32079_, _32078_, _04920_);
  and (_32080_, _32079_, _32077_);
  or (_32081_, _32080_, _31899_);
  nand (_32083_, _32081_, _01995_);
  and (_32084_, _10219_, _01994_);
  nor (_32085_, _32084_, _07239_);
  nand (_32086_, _32085_, _32083_);
  and (_32087_, _07239_, _01825_);
  nor (_32088_, _32087_, _10149_);
  nand (_32089_, _32088_, _32086_);
  nor (_32090_, _10150_, _01845_);
  nor (_32091_, _32090_, _02123_);
  and (_32092_, _32091_, _32089_);
  and (_32094_, _02123_, _01825_);
  or (_32095_, _32094_, _01718_);
  or (_32096_, _32095_, _32092_);
  and (_32097_, _02324_, _01718_);
  nor (_32098_, _32097_, _10604_);
  nand (_32099_, _32098_, _32096_);
  and (_32100_, _07587_, _01825_);
  and (_32101_, _31915_, _10611_);
  or (_32102_, _32101_, _32100_);
  and (_32103_, _32102_, _10604_);
  nor (_32104_, _32103_, _10609_);
  and (_32105_, _32104_, _32099_);
  or (_32106_, _32105_, _31898_);
  nand (_32107_, _32106_, _10618_);
  nor (_32108_, _10618_, _01825_);
  nor (_32109_, _32108_, _02210_);
  and (_32110_, _32109_, _32107_);
  and (_32111_, _10218_, _02210_);
  or (_32112_, _32111_, _02331_);
  nor (_32113_, _32112_, _32110_);
  and (_32115_, _02331_, _02264_);
  or (_32116_, _32115_, _32113_);
  nand (_32117_, _32116_, _30883_);
  and (_32118_, _02324_, _01722_);
  nor (_32119_, _32118_, _10629_);
  nand (_32120_, _32119_, _32117_);
  nor (_32121_, _07587_, _02264_);
  and (_32122_, _31915_, _07587_);
  or (_32123_, _32122_, _32121_);
  and (_32124_, _32123_, _10629_);
  nor (_32126_, _32124_, _10634_);
  and (_32127_, _32126_, _32120_);
  or (_32128_, _32127_, _31897_);
  nand (_32129_, _32128_, _10135_);
  nor (_32130_, _10135_, _01825_);
  nor (_32131_, _32130_, _02206_);
  and (_32132_, _32131_, _32129_);
  and (_32133_, _10218_, _02206_);
  or (_32134_, _32133_, _02342_);
  nor (_32135_, _32134_, _32132_);
  and (_32137_, _02342_, _02264_);
  or (_32138_, _32137_, _32135_);
  nand (_32139_, _32138_, _30879_);
  and (_32140_, _02324_, _01728_);
  nor (_32141_, _32140_, _10649_);
  nand (_32142_, _32141_, _32139_);
  or (_32143_, _31915_, \oc8051_golden_model_1.PSW [7]);
  or (_32144_, _01825_, _06707_);
  and (_32145_, _32144_, _10649_);
  and (_32146_, _32145_, _32143_);
  nor (_32148_, _32146_, _10654_);
  and (_32149_, _32148_, _32142_);
  or (_32150_, _32149_, _31895_);
  nand (_32151_, _32150_, _07339_);
  nor (_32152_, _07339_, _01825_);
  nor (_32153_, _32152_, _02202_);
  and (_32154_, _32153_, _32151_);
  and (_32155_, _10218_, _02202_);
  or (_32156_, _32155_, _02334_);
  nor (_32157_, _32156_, _32154_);
  and (_32159_, _02334_, _02264_);
  or (_32160_, _32159_, _32157_);
  nand (_32161_, _32160_, _30876_);
  and (_32162_, _02324_, _01736_);
  nor (_32163_, _32162_, _10122_);
  nand (_32164_, _32163_, _32161_);
  nor (_32165_, _31915_, _06707_);
  nor (_32166_, _01825_, \oc8051_golden_model_1.PSW [7]);
  nor (_32167_, _32166_, _10123_);
  not (_32168_, _32167_);
  nor (_32170_, _32168_, _32165_);
  nor (_32171_, _32170_, _10671_);
  and (_32172_, _32171_, _32164_);
  or (_32173_, _32172_, _31894_);
  nand (_32174_, _32173_, _07385_);
  nor (_32175_, _07385_, _01825_);
  nor (_32176_, _32175_, _07415_);
  nand (_32177_, _32176_, _32174_);
  and (_32178_, _07415_, _02266_);
  nor (_32179_, _32178_, _02350_);
  and (_32181_, _32179_, _32177_);
  nor (_32182_, _05166_, _09472_);
  or (_32183_, _32182_, _32181_);
  nand (_32184_, _32183_, _04964_);
  and (_32185_, _02324_, _01726_);
  nor (_32186_, _32185_, _02200_);
  nand (_32187_, _32186_, _32184_);
  and (_32188_, _31989_, _08690_);
  nor (_32189_, _10218_, _08690_);
  or (_32190_, _32189_, _10689_);
  nor (_32192_, _32190_, _32188_);
  nor (_32193_, _32192_, _10693_);
  and (_32194_, _32193_, _32187_);
  or (_32195_, _32194_, _31893_);
  nand (_32196_, _32195_, _07488_);
  nor (_32197_, _07488_, _01825_);
  nor (_32198_, _32197_, _07533_);
  nand (_32199_, _32198_, _32196_);
  and (_32200_, _07533_, _02266_);
  nor (_32201_, _32200_, _02083_);
  and (_32203_, _32201_, _32199_);
  nor (_32204_, _05166_, _02084_);
  or (_32205_, _32204_, _32203_);
  nand (_32206_, _32205_, _10712_);
  and (_32207_, _02324_, _01738_);
  nor (_32208_, _32207_, _02243_);
  nand (_32209_, _32208_, _32206_);
  nor (_32210_, _31906_, _08690_);
  and (_32211_, _10219_, _08690_);
  nor (_32212_, _32211_, _32210_);
  and (_32214_, _32212_, _02243_);
  nor (_32215_, _32214_, _10723_);
  nand (_32216_, _32215_, _32209_);
  nor (_32217_, _10722_, _02266_);
  nor (_32218_, _32217_, _02366_);
  and (_32219_, _32218_, _32216_);
  or (_32220_, _32219_, _31892_);
  nand (_32221_, _32220_, _07581_);
  nor (_32222_, _07581_, _01830_);
  nor (_32223_, _32222_, _03537_);
  nand (_32225_, _32223_, _32221_);
  and (_32226_, _03537_, _02324_);
  nor (_32227_, _32226_, _01697_);
  nand (_32228_, _32227_, _32225_);
  and (_32229_, _32212_, _01697_);
  nor (_32230_, _32229_, _10744_);
  nand (_32231_, _32230_, _32228_);
  and (_32232_, _10744_, _01830_);
  nor (_32233_, _32232_, _02081_);
  and (_32234_, _32233_, _32231_);
  or (_32236_, _32234_, _31891_);
  nand (_32237_, _32236_, _10751_);
  nor (_32238_, _10751_, _01830_);
  nor (_32239_, _32238_, _30863_);
  nand (_32240_, _32239_, _32237_);
  and (_32241_, _30863_, _02324_);
  nor (_32242_, _32241_, _10762_);
  and (_32243_, _32242_, _32240_);
  and (_32244_, _10762_, _02266_);
  or (_32245_, _32244_, _32243_);
  or (_32247_, _32245_, _39633_);
  or (_32248_, _39632_, \oc8051_golden_model_1.PC [3]);
  and (_32249_, _32248_, _39026_);
  and (_41796_, _32249_, _32247_);
  not (_32250_, \oc8051_golden_model_1.PC [4]);
  nor (_32251_, _01426_, _32250_);
  and (_32252_, _01426_, _32250_);
  nor (_32253_, _32252_, _32251_);
  not (_32254_, _32253_);
  and (_32255_, _32254_, _10744_);
  nor (_32257_, _10374_, _07587_);
  and (_32258_, _10394_, _10391_);
  nor (_32259_, _32258_, _10395_);
  and (_32260_, _32259_, _07587_);
  or (_32261_, _32260_, _32257_);
  and (_32262_, _32261_, _10629_);
  nor (_32263_, _10373_, _04919_);
  and (_32264_, _10214_, _02218_);
  nor (_32265_, _31255_, _10373_);
  and (_32266_, _10374_, _02053_);
  nor (_32267_, _32253_, _10452_);
  and (_32268_, _10242_, _10239_);
  nor (_32269_, _32268_, _10243_);
  or (_32270_, _32269_, _10293_);
  or (_32271_, _10295_, _10214_);
  and (_32272_, _32271_, _02158_);
  and (_32273_, _32272_, _32270_);
  and (_32274_, _10435_, _10373_);
  and (_32275_, _32259_, _10437_);
  nor (_32276_, _32275_, _32274_);
  nand (_32278_, _32276_, _04535_);
  not (_32279_, _10442_);
  and (_32280_, _04784_, _02060_);
  and (_32281_, _10374_, _02062_);
  or (_32282_, _32281_, _06855_);
  or (_32283_, _10301_, _32250_);
  and (_32284_, _32283_, _02063_);
  or (_32285_, _32284_, _32282_);
  or (_32286_, _32254_, _10312_);
  and (_32287_, _32286_, _01747_);
  and (_32289_, _32287_, _32285_);
  or (_32290_, _32289_, _31555_);
  or (_32291_, _32290_, _32280_);
  or (_32292_, _32254_, _06859_);
  and (_32293_, _32292_, _06847_);
  and (_32294_, _32293_, _32291_);
  and (_32295_, _10374_, _02160_);
  or (_32296_, _32295_, _32294_);
  nor (_32297_, _32296_, _06845_);
  and (_32298_, _32253_, _06845_);
  or (_32300_, _32298_, _32297_);
  and (_32301_, _32300_, _01752_);
  nor (_32302_, _04784_, _01752_);
  nor (_32303_, _32302_, _04535_);
  not (_32304_, _32303_);
  nor (_32305_, _32304_, _32301_);
  nor (_32306_, _32305_, _32279_);
  and (_32307_, _32306_, _32278_);
  or (_32308_, _32307_, _32273_);
  and (_32309_, _32308_, _10287_);
  nor (_32311_, _32254_, _10448_);
  or (_32312_, _32311_, _02057_);
  or (_32313_, _32312_, _32309_);
  and (_32314_, _10374_, _02057_);
  nor (_32315_, _32314_, _03446_);
  and (_32316_, _32315_, _32313_);
  nor (_32317_, _04784_, _01745_);
  or (_32318_, _32317_, _02155_);
  nor (_32319_, _32318_, _32316_);
  and (_32320_, _10374_, _02155_);
  or (_32322_, _32320_, _32319_);
  and (_32323_, _32322_, _10452_);
  or (_32324_, _32323_, _32267_);
  nand (_32325_, _32324_, _02549_);
  and (_32326_, _10374_, _02153_);
  nor (_32327_, _32326_, _10462_);
  nand (_32328_, _32327_, _32325_);
  nor (_32329_, _32254_, _10460_);
  nor (_32330_, _32329_, _02053_);
  and (_32331_, _32330_, _32328_);
  or (_32333_, _32331_, _32266_);
  nand (_32334_, _32333_, _01757_);
  and (_32335_, _04784_, _10464_);
  nor (_32336_, _32335_, _02052_);
  nand (_32337_, _32336_, _32334_);
  and (_32338_, _10373_, _02052_);
  nor (_32339_, _32338_, _10475_);
  nand (_32340_, _32339_, _32337_);
  and (_32341_, _10214_, _08770_);
  not (_32342_, _32269_);
  nor (_32344_, _32342_, _08770_);
  or (_32345_, _32344_, _10471_);
  nor (_32346_, _32345_, _32341_);
  or (_32347_, _08790_, _02171_);
  nor (_32348_, _32347_, _32346_);
  nand (_32349_, _32348_, _32340_);
  and (_32350_, _10214_, _08877_);
  nor (_32351_, _32342_, _08877_);
  nor (_32352_, _32351_, _32350_);
  nor (_32353_, _32352_, _02547_);
  and (_32355_, _10215_, _08842_);
  and (_32356_, _32342_, _10482_);
  nor (_32357_, _32356_, _32355_);
  and (_32358_, _32357_, _08790_);
  nor (_32359_, _32358_, _32353_);
  nand (_32360_, _32359_, _32349_);
  nand (_32361_, _32360_, _08917_);
  and (_32362_, _10215_, _08922_);
  nor (_32363_, _32269_, _08922_);
  or (_32364_, _32363_, _08917_);
  or (_32366_, _32364_, _32362_);
  and (_32367_, _32366_, _08882_);
  and (_32368_, _32367_, _32361_);
  and (_32369_, _32254_, _08881_);
  or (_32370_, _32369_, _32368_);
  nand (_32371_, _32370_, _02047_);
  and (_32372_, _10374_, _02046_);
  nor (_32373_, _32372_, _03310_);
  nand (_32374_, _32373_, _32371_);
  nor (_32375_, _04784_, _01750_);
  nor (_32377_, _32375_, _31256_);
  and (_32378_, _32377_, _32374_);
  or (_32379_, _32378_, _32265_);
  nand (_32380_, _32379_, _10158_);
  nor (_32381_, _32253_, _10158_);
  nor (_32382_, _32381_, _02182_);
  nand (_32383_, _32382_, _32380_);
  and (_32384_, _10373_, _02182_);
  nor (_32385_, _32384_, _10513_);
  nand (_32386_, _32385_, _32383_);
  and (_32388_, _04784_, _10513_);
  nor (_32389_, _32388_, _02181_);
  and (_32390_, _32389_, _32386_);
  and (_32391_, _10373_, _02181_);
  or (_32392_, _32391_, _32390_);
  nand (_32393_, _32392_, _10153_);
  nor (_32394_, _32254_, _10153_);
  nor (_32395_, _32394_, _07017_);
  nand (_32396_, _32395_, _32393_);
  nor (_32397_, _10373_, _07016_);
  nor (_32399_, _32397_, _01876_);
  nand (_32400_, _32399_, _32396_);
  nor (_32401_, _32254_, _01778_);
  nor (_32402_, _32401_, _02042_);
  and (_32403_, _32402_, _32400_);
  and (_32404_, _10374_, _02042_);
  or (_32405_, _32404_, _32403_);
  nand (_32406_, _32405_, _04460_);
  and (_32407_, _04784_, _01767_);
  nor (_32408_, _32407_, _02218_);
  nand (_32410_, _32408_, _32406_);
  nand (_32411_, _32410_, _10534_);
  or (_32412_, _32411_, _32264_);
  nor (_32413_, _10373_, _10534_);
  nor (_32414_, _32413_, _01765_);
  nand (_32415_, _32414_, _32412_);
  and (_32416_, _10214_, _01765_);
  nor (_32417_, _32416_, _10546_);
  nand (_32418_, _32417_, _32415_);
  nor (_32419_, _32253_, _10542_);
  nor (_32421_, _32419_, _02124_);
  nand (_32422_, _32421_, _32418_);
  and (_32423_, _10373_, _02124_);
  nor (_32424_, _32423_, _01711_);
  nand (_32425_, _32424_, _32422_);
  and (_32426_, _04784_, _01711_);
  nor (_32427_, _32426_, _10550_);
  nand (_32428_, _32427_, _32425_);
  and (_32429_, _32259_, _10550_);
  nor (_32430_, _32429_, _04920_);
  and (_32431_, _32430_, _32428_);
  or (_32432_, _32431_, _32263_);
  nand (_32433_, _32432_, _01995_);
  and (_32434_, _10215_, _01994_);
  nor (_32435_, _32434_, _07239_);
  and (_32436_, _32435_, _32433_);
  and (_32437_, _10373_, _07239_);
  or (_32438_, _32437_, _32436_);
  nand (_32439_, _32438_, _10150_);
  and (_32440_, _10580_, _10577_);
  nor (_32442_, _32440_, _10581_);
  and (_32443_, _32442_, _10149_);
  nor (_32444_, _32443_, _02123_);
  and (_32445_, _32444_, _32439_);
  and (_32446_, _10374_, _02123_);
  or (_32447_, _32446_, _32445_);
  nand (_32448_, _32447_, _03308_);
  and (_32449_, _04784_, _01718_);
  nor (_32450_, _32449_, _10604_);
  and (_32451_, _32450_, _32448_);
  and (_32453_, _10373_, _07587_);
  and (_32454_, _32259_, _10611_);
  or (_32455_, _32454_, _32453_);
  and (_32456_, _32455_, _10604_);
  or (_32457_, _32456_, _32451_);
  nand (_32458_, _32457_, _10147_);
  nor (_32459_, _32254_, _10147_);
  nor (_32460_, _32459_, _10619_);
  nand (_32461_, _32460_, _32458_);
  nor (_32462_, _10618_, _10373_);
  nor (_32464_, _32462_, _02210_);
  nand (_32465_, _32464_, _32461_);
  and (_32466_, _10214_, _02210_);
  nor (_32467_, _32466_, _02331_);
  and (_32468_, _32467_, _32465_);
  and (_32469_, _10374_, _02331_);
  or (_32470_, _32469_, _32468_);
  nand (_32471_, _32470_, _30883_);
  and (_32472_, _04784_, _01722_);
  nor (_32473_, _32472_, _10629_);
  and (_32475_, _32473_, _32471_);
  or (_32476_, _32475_, _32262_);
  nand (_32477_, _32476_, _10139_);
  nor (_32478_, _32254_, _10139_);
  nor (_32479_, _32478_, _10136_);
  nand (_32480_, _32479_, _32477_);
  nor (_32481_, _10373_, _10135_);
  nor (_32482_, _32481_, _02206_);
  nand (_32483_, _32482_, _32480_);
  and (_32484_, _10214_, _02206_);
  nor (_32486_, _32484_, _02342_);
  and (_32487_, _32486_, _32483_);
  and (_32488_, _10374_, _02342_);
  or (_32489_, _32488_, _32487_);
  nand (_32490_, _32489_, _30879_);
  and (_32491_, _04784_, _01728_);
  nor (_32492_, _32491_, _10649_);
  nand (_32493_, _32492_, _32490_);
  nand (_32494_, _10373_, \oc8051_golden_model_1.PSW [7]);
  nand (_32495_, _32259_, _06707_);
  and (_32497_, _32495_, _32494_);
  or (_32498_, _32497_, _10650_);
  nand (_32499_, _32498_, _32493_);
  nand (_32500_, _32499_, _10133_);
  nor (_32501_, _32254_, _10133_);
  nor (_32502_, _32501_, _07340_);
  nand (_32503_, _32502_, _32500_);
  nor (_32504_, _10373_, _07339_);
  nor (_32505_, _32504_, _02202_);
  nand (_32506_, _32505_, _32503_);
  and (_32508_, _10214_, _02202_);
  nor (_32509_, _32508_, _02334_);
  and (_32510_, _32509_, _32506_);
  and (_32511_, _10374_, _02334_);
  or (_32512_, _32511_, _32510_);
  nand (_32513_, _32512_, _30876_);
  and (_32514_, _04784_, _01736_);
  nor (_32515_, _32514_, _10122_);
  nand (_32516_, _32515_, _32513_);
  nand (_32517_, _10373_, _06707_);
  nand (_32519_, _32259_, \oc8051_golden_model_1.PSW [7]);
  and (_32520_, _32519_, _32517_);
  or (_32521_, _32520_, _10123_);
  nand (_32522_, _32521_, _32516_);
  nand (_32523_, _32522_, _10120_);
  nor (_32524_, _32254_, _10120_);
  nor (_32525_, _32524_, _07386_);
  nand (_32526_, _32525_, _32523_);
  nor (_32527_, _10373_, _07385_);
  nor (_32528_, _32527_, _07415_);
  nand (_32530_, _32528_, _32526_);
  and (_32531_, _32253_, _07415_);
  nor (_32532_, _32531_, _02350_);
  and (_32533_, _32532_, _32530_);
  nor (_32534_, _05303_, _09472_);
  or (_32535_, _32534_, _32533_);
  nand (_32536_, _32535_, _04964_);
  and (_32537_, _04784_, _01726_);
  nor (_32538_, _32537_, _02200_);
  and (_32539_, _32538_, _32536_);
  nor (_32541_, _10215_, _08690_);
  and (_32542_, _32269_, _08690_);
  nor (_32543_, _32542_, _32541_);
  nor (_32544_, _32543_, _10689_);
  or (_32545_, _32544_, _32539_);
  nand (_32546_, _32545_, _10118_);
  nor (_32547_, _32254_, _10118_);
  nor (_32548_, _32547_, _07489_);
  nand (_32549_, _32548_, _32546_);
  nor (_32550_, _10373_, _07488_);
  nor (_32552_, _32550_, _07533_);
  nand (_32553_, _32552_, _32549_);
  and (_32554_, _32253_, _07533_);
  nor (_32555_, _32554_, _02083_);
  nand (_32556_, _32555_, _32553_);
  nor (_32557_, _05303_, _02084_);
  nor (_32558_, _32557_, _01738_);
  nand (_32559_, _32558_, _32556_);
  nor (_32560_, _04784_, _10712_);
  nor (_32561_, _32560_, _02243_);
  nand (_32562_, _32561_, _32559_);
  and (_32563_, _10215_, _08690_);
  nor (_32564_, _32269_, _08690_);
  nor (_32565_, _32564_, _32563_);
  nor (_32566_, _32565_, _02367_);
  nor (_32567_, _32566_, _10723_);
  nand (_32568_, _32567_, _32562_);
  nor (_32569_, _32254_, _10722_);
  nor (_32570_, _32569_, _02366_);
  nand (_32571_, _32570_, _32568_);
  and (_32573_, _10374_, _02366_);
  nor (_32574_, _32573_, _31858_);
  nand (_32575_, _32574_, _32571_);
  nor (_32576_, _32254_, _07581_);
  nor (_32577_, _32576_, _03537_);
  nand (_32578_, _32577_, _32575_);
  and (_32579_, _04784_, _03537_);
  nor (_32580_, _32579_, _01697_);
  nand (_32581_, _32580_, _32578_);
  and (_32582_, _32565_, _01697_);
  nor (_32584_, _32582_, _10744_);
  and (_32585_, _32584_, _32581_);
  or (_32586_, _32585_, _32255_);
  nand (_32587_, _32586_, _02082_);
  and (_32588_, _10374_, _02081_);
  nor (_32589_, _32588_, _31497_);
  nand (_32590_, _32589_, _32587_);
  nor (_32591_, _32254_, _10751_);
  nor (_32592_, _32591_, _30863_);
  nand (_32593_, _32592_, _32590_);
  and (_32595_, _30863_, _04784_);
  nor (_32596_, _32595_, _10762_);
  nand (_32597_, _32596_, _32593_);
  and (_32598_, _32253_, _10762_);
  not (_32599_, _32598_);
  and (_32600_, _32599_, _32597_);
  nand (_32601_, _32600_, _39632_);
  or (_32602_, _39632_, \oc8051_golden_model_1.PC [4]);
  and (_32603_, _32602_, _39026_);
  and (_41797_, _32603_, _32601_);
  and (_32605_, _10368_, _02081_);
  and (_32606_, _10368_, _02366_);
  nor (_32607_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_32608_, _10368_, _01439_);
  nor (_32609_, _32608_, _32607_);
  nor (_32610_, _32609_, _10118_);
  nor (_32611_, _32609_, _10120_);
  nor (_32612_, _32609_, _10133_);
  nor (_32613_, _32609_, _10139_);
  nor (_32614_, _32609_, _10147_);
  nor (_32616_, _10368_, _04919_);
  nor (_32617_, _31255_, _10368_);
  or (_32618_, _10295_, _10209_);
  or (_32619_, _10212_, _10211_);
  not (_32620_, _32619_);
  nor (_32621_, _32620_, _10244_);
  and (_32622_, _32620_, _10244_);
  nor (_32623_, _32622_, _32621_);
  not (_32624_, _32623_);
  or (_32625_, _32624_, _10293_);
  and (_32627_, _32625_, _32618_);
  or (_32628_, _32627_, _03006_);
  or (_32629_, _10371_, _10370_);
  not (_32630_, _32629_);
  nor (_32631_, _32630_, _10396_);
  and (_32632_, _32630_, _10396_);
  nor (_32633_, _32632_, _32631_);
  nor (_32634_, _32633_, _10435_);
  and (_32635_, _10435_, _10368_);
  nor (_32636_, _32635_, _32634_);
  nand (_32638_, _32636_, _04535_);
  nor (_32639_, _10301_, \oc8051_golden_model_1.PC [5]);
  nor (_32640_, _32639_, _02062_);
  and (_32641_, _10368_, _02062_);
  nor (_32642_, _32641_, _06855_);
  not (_32643_, _32642_);
  nor (_32644_, _32643_, _32640_);
  not (_32645_, _32644_);
  nor (_32646_, _32609_, _10312_);
  nor (_32647_, _32646_, _02060_);
  and (_32649_, _32647_, _32645_);
  nor (_32650_, _04815_, _01747_);
  or (_32651_, _32650_, _31555_);
  nor (_32652_, _32651_, _32649_);
  nor (_32653_, _32609_, _06859_);
  nor (_32654_, _32653_, _02160_);
  not (_32655_, _32654_);
  nor (_32656_, _32655_, _32652_);
  and (_32657_, _10368_, _02160_);
  or (_32658_, _32657_, _32656_);
  and (_32660_, _32658_, _10299_);
  and (_32661_, _32609_, _06845_);
  or (_32662_, _32661_, _32660_);
  and (_32663_, _32662_, _01752_);
  nor (_32664_, _04815_, _01752_);
  or (_32665_, _32664_, _04535_);
  nor (_32666_, _32665_, _32663_);
  nor (_32667_, _32666_, _02079_);
  and (_32668_, _32667_, _32638_);
  and (_32669_, _32609_, _02079_);
  or (_32671_, _32669_, _02158_);
  or (_32672_, _32671_, _32668_);
  nand (_32673_, _32672_, _32628_);
  nand (_32674_, _32673_, _10287_);
  nor (_32675_, _32609_, _10287_);
  nor (_32676_, _32675_, _02057_);
  nand (_32677_, _32676_, _32674_);
  and (_32678_, _10368_, _02057_);
  nor (_32679_, _32678_, _03446_);
  nand (_32680_, _32679_, _32677_);
  and (_32682_, _04815_, _03446_);
  nor (_32683_, _32682_, _02155_);
  nand (_32684_, _32683_, _32680_);
  and (_32685_, _10368_, _02155_);
  nor (_32686_, _32685_, _22169_);
  nand (_32687_, _32686_, _32684_);
  nor (_32688_, _32609_, _10452_);
  nor (_32689_, _32688_, _02153_);
  nand (_32690_, _32689_, _32687_);
  and (_32691_, _10368_, _02153_);
  nor (_32693_, _32691_, _10462_);
  nand (_32694_, _32693_, _32690_);
  nor (_32695_, _32609_, _10460_);
  nor (_32696_, _32695_, _02053_);
  nand (_32697_, _32696_, _32694_);
  and (_32698_, _10368_, _02053_);
  nor (_32699_, _32698_, _10464_);
  nand (_32700_, _32699_, _32697_);
  and (_32701_, _04815_, _10464_);
  nor (_32702_, _32701_, _02052_);
  nand (_32703_, _32702_, _32700_);
  and (_32704_, _10368_, _02052_);
  nor (_32705_, _32704_, _10475_);
  nand (_32706_, _32705_, _32703_);
  and (_32707_, _10209_, _08770_);
  nor (_32708_, _32623_, _08770_);
  or (_32709_, _32708_, _32707_);
  nor (_32710_, _32709_, _10471_);
  nor (_32711_, _32710_, _08790_);
  nand (_32712_, _32711_, _32706_);
  or (_32713_, _32623_, _08842_);
  or (_32714_, _10210_, _10482_);
  nand (_32715_, _32714_, _32713_);
  nand (_32716_, _32715_, _08790_);
  and (_32717_, _32716_, _02547_);
  nand (_32718_, _32717_, _32712_);
  nor (_32719_, _32623_, _08877_);
  not (_32720_, _32719_);
  and (_32721_, _10209_, _08877_);
  nor (_32722_, _32721_, _02547_);
  and (_32723_, _32722_, _32720_);
  nor (_32724_, _32723_, _02246_);
  nand (_32725_, _32724_, _32718_);
  nand (_32726_, _10209_, _08922_);
  or (_32727_, _32623_, _08922_);
  and (_32728_, _32727_, _32726_);
  or (_32729_, _32728_, _08917_);
  and (_32730_, _32729_, _32725_);
  or (_32731_, _32730_, _08881_);
  nand (_32732_, _32609_, _08881_);
  and (_32734_, _32732_, _32731_);
  nand (_32735_, _32734_, _02047_);
  and (_32736_, _10369_, _02046_);
  nor (_32737_, _32736_, _03310_);
  nand (_32738_, _32737_, _32735_);
  nor (_32739_, _04815_, _01750_);
  nor (_32740_, _32739_, _31256_);
  and (_32741_, _32740_, _32738_);
  or (_32742_, _32741_, _32617_);
  nand (_32743_, _32742_, _10158_);
  nor (_32745_, _32609_, _10158_);
  nor (_32746_, _32745_, _02182_);
  nand (_32747_, _32746_, _32743_);
  and (_32748_, _10368_, _02182_);
  nor (_32749_, _32748_, _10513_);
  nand (_32750_, _32749_, _32747_);
  and (_32751_, _04815_, _10513_);
  nor (_32752_, _32751_, _02181_);
  nand (_32753_, _32752_, _32750_);
  and (_32754_, _10368_, _02181_);
  nor (_32755_, _32754_, _10517_);
  and (_32756_, _32755_, _32753_);
  nor (_32757_, _32609_, _10153_);
  or (_32758_, _32757_, _32756_);
  nand (_32759_, _32758_, _07016_);
  nor (_32760_, _10368_, _07016_);
  nor (_32761_, _32760_, _01876_);
  and (_32762_, _32761_, _32759_);
  not (_32763_, _32609_);
  nor (_32764_, _32763_, _01778_);
  or (_32766_, _32764_, _02042_);
  nor (_32767_, _32766_, _32762_);
  and (_32768_, _10369_, _02042_);
  or (_32769_, _32768_, _32767_);
  nand (_32770_, _32769_, _04460_);
  and (_32771_, _04815_, _01767_);
  nor (_32772_, _32771_, _02218_);
  nand (_32773_, _32772_, _32770_);
  and (_32774_, _10209_, _02218_);
  not (_32775_, _32774_);
  and (_32777_, _32775_, _10534_);
  nand (_32778_, _32777_, _32773_);
  nor (_32779_, _10368_, _10534_);
  nor (_32780_, _32779_, _01765_);
  nand (_32781_, _32780_, _32778_);
  and (_32782_, _10209_, _01765_);
  nor (_32783_, _32782_, _10546_);
  nand (_32784_, _32783_, _32781_);
  nor (_32785_, _32609_, _10542_);
  nor (_32786_, _32785_, _02124_);
  nand (_32788_, _32786_, _32784_);
  and (_32789_, _10368_, _02124_);
  nor (_32790_, _32789_, _01711_);
  nand (_32791_, _32790_, _32788_);
  and (_32792_, _04815_, _01711_);
  nor (_32793_, _32792_, _10550_);
  nand (_32794_, _32793_, _32791_);
  nor (_32795_, _32633_, _10551_);
  nor (_32796_, _32795_, _04920_);
  and (_32797_, _32796_, _32794_);
  or (_32799_, _32797_, _32616_);
  nand (_32800_, _32799_, _01995_);
  and (_32801_, _10210_, _01994_);
  nor (_32802_, _32801_, _07239_);
  nand (_32803_, _32802_, _32800_);
  and (_32804_, _10368_, _07239_);
  nor (_32805_, _32804_, _10149_);
  nand (_32806_, _32805_, _32803_);
  and (_32807_, _10582_, _10575_);
  nor (_32808_, _32807_, _10583_);
  nor (_32810_, _32808_, _10150_);
  nor (_32811_, _32810_, _02123_);
  nand (_32812_, _32811_, _32806_);
  and (_32813_, _10368_, _02123_);
  nor (_32814_, _32813_, _01718_);
  nand (_32815_, _32814_, _32812_);
  and (_32816_, _04815_, _01718_);
  nor (_32817_, _32816_, _10604_);
  nand (_32818_, _32817_, _32815_);
  and (_32819_, _32633_, _10611_);
  and (_32821_, _10369_, _07587_);
  nor (_32822_, _32821_, _10605_);
  not (_32823_, _32822_);
  nor (_32824_, _32823_, _32819_);
  nor (_32825_, _32824_, _10609_);
  and (_32826_, _32825_, _32818_);
  or (_32827_, _32826_, _32614_);
  nand (_32828_, _32827_, _10618_);
  nor (_32829_, _10618_, _10368_);
  nor (_32830_, _32829_, _02210_);
  nand (_32832_, _32830_, _32828_);
  and (_32833_, _10209_, _02210_);
  nor (_32834_, _32833_, _02331_);
  and (_32835_, _32834_, _32832_);
  and (_32836_, _10369_, _02331_);
  or (_32837_, _32836_, _32835_);
  nand (_32838_, _32837_, _30883_);
  and (_32839_, _04815_, _01722_);
  nor (_32840_, _32839_, _10629_);
  nand (_32841_, _32840_, _32838_);
  and (_32843_, _10368_, _10611_);
  nor (_32844_, _32633_, _10611_);
  or (_32845_, _32844_, _32843_);
  and (_32846_, _32845_, _10629_);
  nor (_32847_, _32846_, _10634_);
  and (_32848_, _32847_, _32841_);
  or (_32849_, _32848_, _32613_);
  nand (_32850_, _32849_, _10135_);
  nor (_32851_, _10368_, _10135_);
  nor (_32852_, _32851_, _02206_);
  nand (_32854_, _32852_, _32850_);
  and (_32855_, _10209_, _02206_);
  nor (_32856_, _32855_, _02342_);
  and (_32857_, _32856_, _32854_);
  and (_32858_, _10369_, _02342_);
  or (_32859_, _32858_, _32857_);
  nand (_32860_, _32859_, _30879_);
  and (_32861_, _04815_, _01728_);
  nor (_32862_, _32861_, _10649_);
  nand (_32863_, _32862_, _32860_);
  nand (_32865_, _32633_, _06707_);
  or (_32866_, _10368_, _06707_);
  and (_32867_, _32866_, _10649_);
  and (_32868_, _32867_, _32865_);
  nor (_32869_, _32868_, _10654_);
  and (_32870_, _32869_, _32863_);
  or (_32871_, _32870_, _32612_);
  nand (_32872_, _32871_, _07339_);
  nor (_32873_, _10368_, _07339_);
  nor (_32874_, _32873_, _02202_);
  nand (_32876_, _32874_, _32872_);
  and (_32877_, _10209_, _02202_);
  nor (_32878_, _32877_, _02334_);
  and (_32879_, _32878_, _32876_);
  and (_32880_, _10369_, _02334_);
  or (_32881_, _32880_, _32879_);
  nand (_32882_, _32881_, _30876_);
  and (_32883_, _04815_, _01736_);
  nor (_32884_, _32883_, _10122_);
  nand (_32885_, _32884_, _32882_);
  and (_32887_, _10368_, _06707_);
  nor (_32888_, _32633_, _06707_);
  or (_32889_, _32888_, _32887_);
  and (_32890_, _32889_, _10122_);
  nor (_32891_, _32890_, _10671_);
  and (_32892_, _32891_, _32885_);
  or (_32893_, _32892_, _32611_);
  nand (_32894_, _32893_, _07385_);
  nor (_32895_, _10368_, _07385_);
  nor (_32896_, _32895_, _07415_);
  nand (_32898_, _32896_, _32894_);
  and (_32899_, _32609_, _07415_);
  nor (_32900_, _32899_, _02350_);
  and (_32901_, _32900_, _32898_);
  nor (_32902_, _05258_, _09472_);
  or (_32903_, _32902_, _32901_);
  nand (_32904_, _32903_, _04964_);
  and (_32905_, _04815_, _01726_);
  nor (_32906_, _32905_, _02200_);
  nand (_32907_, _32906_, _32904_);
  and (_32909_, _32623_, _08690_);
  nor (_32910_, _10209_, _08690_);
  or (_32911_, _32910_, _10689_);
  nor (_32912_, _32911_, _32909_);
  nor (_32913_, _32912_, _10693_);
  and (_32914_, _32913_, _32907_);
  or (_32915_, _32914_, _32610_);
  nand (_32916_, _32915_, _07488_);
  nor (_32917_, _10368_, _07488_);
  nor (_32918_, _32917_, _07533_);
  nand (_32920_, _32918_, _32916_);
  and (_32921_, _32609_, _07533_);
  nor (_32922_, _32921_, _02083_);
  and (_32923_, _32922_, _32920_);
  nor (_32924_, _05258_, _02084_);
  or (_32925_, _32924_, _32923_);
  nand (_32926_, _32925_, _10712_);
  and (_32927_, _04815_, _01738_);
  nor (_32928_, _32927_, _02243_);
  nand (_32929_, _32928_, _32926_);
  and (_32931_, _10210_, _08690_);
  nor (_32932_, _32624_, _08690_);
  nor (_32933_, _32932_, _32931_);
  and (_32934_, _32933_, _02243_);
  nor (_32935_, _32934_, _10723_);
  nand (_32936_, _32935_, _32929_);
  nor (_32937_, _32609_, _10722_);
  nor (_32938_, _32937_, _02366_);
  and (_32939_, _32938_, _32936_);
  or (_32940_, _32939_, _32606_);
  nand (_32942_, _32940_, _07581_);
  nor (_32943_, _32763_, _07581_);
  nor (_32944_, _32943_, _03537_);
  nand (_32945_, _32944_, _32942_);
  and (_32946_, _04815_, _03537_);
  nor (_32947_, _32946_, _01697_);
  nand (_32948_, _32947_, _32945_);
  and (_32949_, _32933_, _01697_);
  nor (_32950_, _32949_, _10744_);
  nand (_32951_, _32950_, _32948_);
  and (_32953_, _32763_, _10744_);
  nor (_32954_, _32953_, _02081_);
  and (_32955_, _32954_, _32951_);
  or (_32956_, _32955_, _32605_);
  nand (_32957_, _32956_, _10751_);
  nor (_32958_, _32763_, _10751_);
  nor (_32959_, _32958_, _30863_);
  nand (_32960_, _32959_, _32957_);
  and (_32961_, _30863_, _04815_);
  nor (_32962_, _32961_, _10762_);
  nand (_32964_, _32962_, _32960_);
  and (_32965_, _32609_, _10762_);
  not (_32966_, _32965_);
  and (_32967_, _32966_, _32964_);
  nand (_32968_, _32967_, _39632_);
  or (_32969_, _39632_, \oc8051_golden_model_1.PC [5]);
  and (_32970_, _32969_, _39026_);
  and (_41798_, _32970_, _32968_);
  and (_32971_, _04752_, _03537_);
  and (_32972_, _04538_, _10107_);
  and (_32974_, _32972_, \oc8051_golden_model_1.PC [6]);
  nor (_32975_, _32972_, \oc8051_golden_model_1.PC [6]);
  nor (_32976_, _32975_, _32974_);
  not (_32977_, _32976_);
  and (_32978_, _32977_, _07533_);
  and (_32979_, _10202_, _02218_);
  nor (_32980_, _31255_, _10360_);
  and (_32981_, _32977_, _08881_);
  and (_32982_, _10201_, _08877_);
  and (_32983_, _10246_, _10206_);
  nor (_32985_, _32983_, _10247_);
  not (_32986_, _32985_);
  nor (_32987_, _32986_, _08877_);
  nor (_32988_, _32987_, _32982_);
  or (_32989_, _32988_, _02547_);
  and (_32990_, _10361_, _02053_);
  nor (_32991_, _32976_, _10452_);
  or (_32992_, _32985_, _10293_);
  or (_32993_, _10295_, _10201_);
  and (_32994_, _32993_, _02158_);
  and (_32996_, _32994_, _32992_);
  and (_32997_, _10435_, _10360_);
  and (_32998_, _10398_, _10365_);
  nor (_32999_, _32998_, _10399_);
  and (_33000_, _32999_, _10437_);
  nor (_33001_, _33000_, _32997_);
  nand (_33002_, _33001_, _04535_);
  and (_33003_, _04752_, _02060_);
  and (_33004_, _10361_, _02062_);
  or (_33005_, _33004_, _06855_);
  nand (_33007_, _10302_, \oc8051_golden_model_1.PC [6]);
  and (_33008_, _33007_, _02063_);
  or (_33009_, _33008_, _33005_);
  or (_33010_, _32977_, _10312_);
  and (_33011_, _33010_, _01747_);
  and (_33012_, _33011_, _33009_);
  or (_33013_, _33012_, _31555_);
  or (_33014_, _33013_, _33003_);
  or (_33015_, _32977_, _06859_);
  and (_33016_, _33015_, _06847_);
  and (_33018_, _33016_, _33014_);
  and (_33019_, _10361_, _02160_);
  or (_33020_, _33019_, _33018_);
  nor (_33021_, _33020_, _06845_);
  and (_33022_, _32976_, _06845_);
  or (_33023_, _33022_, _33021_);
  and (_33024_, _33023_, _01752_);
  nor (_33025_, _04752_, _01752_);
  nor (_33026_, _33025_, _04535_);
  not (_33027_, _33026_);
  nor (_33029_, _33027_, _33024_);
  nor (_33030_, _33029_, _32279_);
  and (_33031_, _33030_, _33002_);
  or (_33032_, _33031_, _32996_);
  and (_33033_, _33032_, _10287_);
  nor (_33034_, _32977_, _10448_);
  or (_33035_, _33034_, _02057_);
  or (_33036_, _33035_, _33033_);
  and (_33037_, _10361_, _02057_);
  nor (_33038_, _33037_, _03446_);
  and (_33040_, _33038_, _33036_);
  nor (_33041_, _04752_, _01745_);
  or (_33042_, _33041_, _02155_);
  nor (_33043_, _33042_, _33040_);
  and (_33044_, _10361_, _02155_);
  or (_33045_, _33044_, _33043_);
  and (_33046_, _33045_, _10452_);
  or (_33047_, _33046_, _32991_);
  nand (_33048_, _33047_, _02549_);
  and (_33049_, _10361_, _02153_);
  nor (_33051_, _33049_, _10462_);
  nand (_33052_, _33051_, _33048_);
  nor (_33053_, _32977_, _10460_);
  nor (_33054_, _33053_, _02053_);
  and (_33055_, _33054_, _33052_);
  or (_33056_, _33055_, _32990_);
  nand (_33057_, _33056_, _01757_);
  and (_33058_, _04752_, _10464_);
  nor (_33059_, _33058_, _02052_);
  nand (_33060_, _33059_, _33057_);
  and (_33062_, _10360_, _02052_);
  nor (_33063_, _33062_, _10475_);
  and (_33064_, _33063_, _33060_);
  and (_33065_, _10201_, _08770_);
  nor (_33066_, _32986_, _08770_);
  or (_33067_, _33066_, _33065_);
  nor (_33068_, _33067_, _10471_);
  or (_33069_, _33068_, _33064_);
  and (_33070_, _33069_, _08836_);
  and (_33071_, _10201_, _08842_);
  and (_33073_, _32985_, _10482_);
  or (_33074_, _33073_, _08836_);
  nor (_33075_, _33074_, _33071_);
  or (_33076_, _33075_, _33070_);
  or (_33077_, _33076_, _02171_);
  and (_33078_, _33077_, _32989_);
  or (_33079_, _33078_, _02246_);
  and (_33080_, _10201_, _08922_);
  and (_33081_, _32985_, _32011_);
  nor (_33082_, _33081_, _33080_);
  nor (_33084_, _33082_, _08917_);
  nor (_33085_, _33084_, _08881_);
  and (_33086_, _33085_, _33079_);
  or (_33087_, _33086_, _32981_);
  nand (_33088_, _33087_, _02047_);
  and (_33089_, _10361_, _02046_);
  nor (_33090_, _33089_, _03310_);
  nand (_33091_, _33090_, _33088_);
  nor (_33092_, _04752_, _01750_);
  nor (_33093_, _33092_, _31256_);
  and (_33095_, _33093_, _33091_);
  or (_33096_, _33095_, _32980_);
  nand (_33097_, _33096_, _10158_);
  nor (_33098_, _32976_, _10158_);
  nor (_33099_, _33098_, _02182_);
  nand (_33100_, _33099_, _33097_);
  and (_33101_, _10360_, _02182_);
  not (_33102_, _33101_);
  and (_33103_, _33102_, _10514_);
  and (_33104_, _33103_, _33100_);
  and (_33106_, _04752_, _10513_);
  and (_33107_, _10361_, _02181_);
  or (_33108_, _33107_, _33106_);
  or (_33109_, _33108_, _33104_);
  nand (_33110_, _33109_, _10153_);
  nor (_33111_, _32976_, _10153_);
  nor (_33112_, _33111_, _07017_);
  and (_33113_, _33112_, _33110_);
  nor (_33114_, _10361_, _07016_);
  or (_33115_, _33114_, _01876_);
  nor (_33116_, _33115_, _33113_);
  nor (_33117_, _32976_, _01778_);
  or (_33118_, _33117_, _33116_);
  nand (_33119_, _33118_, _02043_);
  and (_33120_, _10361_, _02042_);
  nor (_33121_, _33120_, _01767_);
  nand (_33122_, _33121_, _33119_);
  nor (_33123_, _04752_, _04460_);
  nor (_33124_, _33123_, _02218_);
  nand (_33125_, _33124_, _33122_);
  nand (_33127_, _33125_, _10534_);
  or (_33128_, _33127_, _32979_);
  nor (_33129_, _10361_, _10534_);
  nor (_33130_, _33129_, _01765_);
  nand (_33131_, _33130_, _33128_);
  and (_33132_, _10202_, _01765_);
  nor (_33133_, _33132_, _10546_);
  nand (_33134_, _33133_, _33131_);
  nor (_33135_, _32977_, _10542_);
  nor (_33136_, _33135_, _02124_);
  and (_33138_, _33136_, _33134_);
  and (_33139_, _10361_, _02124_);
  or (_33140_, _33139_, _33138_);
  nand (_33141_, _33140_, _01712_);
  and (_33142_, _04752_, _01711_);
  nor (_33143_, _33142_, _10550_);
  nand (_33144_, _33143_, _33141_);
  and (_33145_, _32999_, _10550_);
  nor (_33146_, _33145_, _04920_);
  and (_33147_, _33146_, _33144_);
  nor (_33149_, _10360_, _04919_);
  or (_33150_, _33149_, _33147_);
  nand (_33151_, _33150_, _01995_);
  and (_33152_, _10202_, _01994_);
  nor (_33153_, _33152_, _07239_);
  nand (_33154_, _33153_, _33151_);
  and (_33155_, _10360_, _07239_);
  nor (_33156_, _33155_, _10149_);
  nand (_33157_, _33156_, _33154_);
  and (_33158_, _10584_, _10571_);
  nor (_33160_, _33158_, _10585_);
  nor (_33161_, _33160_, _10150_);
  nor (_33162_, _33161_, _02123_);
  nand (_33163_, _33162_, _33157_);
  and (_33164_, _10360_, _02123_);
  nor (_33165_, _33164_, _01718_);
  nand (_33166_, _33165_, _33163_);
  and (_33167_, _04752_, _01718_);
  nor (_33168_, _33167_, _10604_);
  nand (_33169_, _33168_, _33166_);
  nor (_33171_, _32999_, _07587_);
  and (_33172_, _10361_, _07587_);
  nor (_33173_, _33172_, _10605_);
  not (_33174_, _33173_);
  nor (_33175_, _33174_, _33171_);
  nor (_33176_, _33175_, _10609_);
  nand (_33177_, _33176_, _33169_);
  nor (_33178_, _32976_, _10147_);
  nor (_33179_, _33178_, _10619_);
  nand (_33180_, _33179_, _33177_);
  nor (_33182_, _10618_, _10361_);
  nor (_33183_, _33182_, _02210_);
  and (_33184_, _33183_, _33180_);
  and (_33185_, _10202_, _02210_);
  or (_33186_, _33185_, _33184_);
  nand (_33187_, _33186_, _03061_);
  and (_33188_, _10361_, _02331_);
  nor (_33189_, _33188_, _01722_);
  and (_33190_, _33189_, _33187_);
  nor (_33191_, _04752_, _30883_);
  or (_33193_, _33191_, _33190_);
  nand (_33194_, _33193_, _10630_);
  and (_33195_, _10360_, _10611_);
  and (_33196_, _32999_, _07587_);
  or (_33197_, _33196_, _33195_);
  and (_33198_, _33197_, _10629_);
  nor (_33199_, _33198_, _10634_);
  nand (_33200_, _33199_, _33194_);
  nor (_33201_, _32976_, _10139_);
  nor (_33202_, _33201_, _10136_);
  nand (_33204_, _33202_, _33200_);
  nor (_33205_, _10361_, _10135_);
  nor (_33206_, _33205_, _02206_);
  and (_33207_, _33206_, _33204_);
  and (_33208_, _10202_, _02206_);
  or (_33209_, _33208_, _33207_);
  nand (_33210_, _33209_, _03065_);
  and (_33211_, _10361_, _02342_);
  nor (_33212_, _33211_, _01728_);
  and (_33213_, _33212_, _33210_);
  nor (_33215_, _04752_, _30879_);
  or (_33216_, _33215_, _33213_);
  nand (_33217_, _33216_, _10650_);
  or (_33218_, _32999_, \oc8051_golden_model_1.PSW [7]);
  or (_33219_, _10360_, _06707_);
  and (_33220_, _33219_, _10649_);
  and (_33221_, _33220_, _33218_);
  nor (_33222_, _33221_, _10654_);
  nand (_33223_, _33222_, _33217_);
  nor (_33224_, _32976_, _10133_);
  nor (_33226_, _33224_, _07340_);
  nand (_33227_, _33226_, _33223_);
  nor (_33228_, _10361_, _07339_);
  nor (_33229_, _33228_, _02202_);
  and (_33230_, _33229_, _33227_);
  and (_33231_, _10202_, _02202_);
  or (_33232_, _33231_, _33230_);
  nand (_33233_, _33232_, _04958_);
  and (_33234_, _10361_, _02334_);
  nor (_33235_, _33234_, _01736_);
  and (_33237_, _33235_, _33233_);
  nor (_33238_, _04752_, _30876_);
  or (_33239_, _33238_, _33237_);
  nand (_33240_, _33239_, _10123_);
  and (_33241_, _10360_, _06707_);
  and (_33242_, _32999_, \oc8051_golden_model_1.PSW [7]);
  or (_33243_, _33242_, _33241_);
  and (_33244_, _33243_, _10122_);
  nor (_33245_, _33244_, _10671_);
  nand (_33246_, _33245_, _33240_);
  nor (_33248_, _32976_, _10120_);
  nor (_33249_, _33248_, _07386_);
  nand (_33250_, _33249_, _33246_);
  nor (_33251_, _10361_, _07385_);
  nor (_33252_, _33251_, _07415_);
  nand (_33253_, _33252_, _33250_);
  and (_33254_, _32977_, _07415_);
  nor (_33255_, _33254_, _02350_);
  nand (_33256_, _33255_, _33253_);
  and (_33257_, _05029_, _02350_);
  nor (_33259_, _33257_, _01726_);
  nand (_33260_, _33259_, _33256_);
  and (_33261_, _04752_, _01726_);
  nor (_33262_, _33261_, _02200_);
  nand (_33263_, _33262_, _33260_);
  and (_33264_, _32986_, _08690_);
  nor (_33265_, _10201_, _08690_);
  or (_33266_, _33265_, _10689_);
  nor (_33267_, _33266_, _33264_);
  nor (_33268_, _33267_, _10693_);
  nand (_33270_, _33268_, _33263_);
  nor (_33271_, _32976_, _10118_);
  nor (_33272_, _33271_, _07489_);
  nand (_33273_, _33272_, _33270_);
  nor (_33274_, _10361_, _07488_);
  nor (_33275_, _33274_, _07533_);
  and (_33276_, _33275_, _33273_);
  or (_33277_, _33276_, _32978_);
  nand (_33278_, _33277_, _02084_);
  nor (_33279_, _05029_, _02084_);
  nor (_33281_, _33279_, _01738_);
  nand (_33282_, _33281_, _33278_);
  nor (_33283_, _04752_, _10712_);
  nor (_33284_, _33283_, _02243_);
  and (_33285_, _33284_, _33282_);
  and (_33286_, _10202_, _08690_);
  nor (_33287_, _32985_, _08690_);
  nor (_33288_, _33287_, _33286_);
  nor (_33289_, _33288_, _02367_);
  or (_33290_, _33289_, _33285_);
  and (_33292_, _33290_, _10722_);
  nor (_33293_, _32976_, _10722_);
  or (_33294_, _33293_, _33292_);
  nand (_33295_, _33294_, _02778_);
  and (_33296_, _10361_, _02366_);
  nor (_33297_, _33296_, _31858_);
  nand (_33298_, _33297_, _33295_);
  nor (_33299_, _32977_, _07581_);
  nor (_33300_, _33299_, _03537_);
  and (_33301_, _33300_, _33298_);
  or (_33303_, _33301_, _32971_);
  nand (_33304_, _33303_, _01698_);
  nor (_33305_, _33288_, _01698_);
  nor (_33306_, _33305_, _10744_);
  nand (_33307_, _33306_, _33304_);
  and (_33308_, _32976_, _10744_);
  nor (_33309_, _33308_, _02081_);
  nand (_33310_, _33309_, _33307_);
  and (_33311_, _10361_, _02081_);
  nor (_33312_, _33311_, _31497_);
  nand (_33314_, _33312_, _33310_);
  nor (_33315_, _32977_, _10751_);
  nor (_33316_, _33315_, _30863_);
  nand (_33317_, _33316_, _33314_);
  and (_33318_, _30863_, _04752_);
  nor (_33319_, _33318_, _10762_);
  nand (_33320_, _33319_, _33317_);
  and (_33321_, _32976_, _10762_);
  not (_33322_, _33321_);
  and (_33323_, _33322_, _33320_);
  nand (_33325_, _33323_, _39632_);
  or (_33326_, _39632_, \oc8051_golden_model_1.PC [6]);
  and (_33327_, _33326_, _39026_);
  and (_41799_, _33327_, _33325_);
  and (_33328_, _04543_, _02081_);
  nor (_33329_, _10108_, \oc8051_golden_model_1.PC [7]);
  nor (_33330_, _33329_, _10109_);
  nor (_33331_, _33330_, _10118_);
  nor (_33332_, _33330_, _10120_);
  nor (_33333_, _33330_, _10133_);
  nor (_33335_, _33330_, _10139_);
  nor (_33336_, _33330_, _10147_);
  nor (_33337_, _04919_, _04543_);
  and (_33338_, _05322_, _02218_);
  nor (_33339_, _31255_, _04543_);
  or (_33340_, _10295_, _05322_);
  or (_33341_, _10197_, _10198_);
  and (_33342_, _33341_, _10248_);
  nor (_33343_, _33341_, _10248_);
  nor (_33344_, _33343_, _33342_);
  or (_33346_, _33344_, _10293_);
  and (_33347_, _33346_, _33340_);
  or (_33348_, _33347_, _03006_);
  and (_33349_, _10435_, _04543_);
  or (_33350_, _10356_, _10357_);
  and (_33351_, _33350_, _10400_);
  nor (_33352_, _33350_, _10400_);
  nor (_33353_, _33352_, _33351_);
  and (_33354_, _33353_, _10437_);
  nor (_33355_, _33354_, _33349_);
  nand (_33357_, _33355_, _04535_);
  nor (_33358_, _10301_, \oc8051_golden_model_1.PC [7]);
  nor (_33359_, _33358_, _02062_);
  and (_33360_, _04543_, _02062_);
  nor (_33361_, _33360_, _06855_);
  not (_33362_, _33361_);
  nor (_33363_, _33362_, _33359_);
  not (_33364_, _33363_);
  nor (_33365_, _33330_, _10312_);
  nor (_33366_, _33365_, _02060_);
  and (_33368_, _33366_, _33364_);
  nor (_33369_, _04458_, _01747_);
  or (_33370_, _33369_, _31555_);
  nor (_33371_, _33370_, _33368_);
  nor (_33372_, _33330_, _06859_);
  nor (_33373_, _33372_, _02160_);
  not (_33374_, _33373_);
  nor (_33375_, _33374_, _33371_);
  and (_33376_, _04543_, _02160_);
  or (_33377_, _33376_, _33375_);
  and (_33379_, _33377_, _10299_);
  and (_33380_, _33330_, _06845_);
  or (_33381_, _33380_, _33379_);
  and (_33382_, _33381_, _01752_);
  nor (_33383_, _04458_, _01752_);
  nor (_33384_, _33383_, _04535_);
  not (_33385_, _33384_);
  nor (_33386_, _33385_, _33382_);
  nor (_33387_, _33386_, _02079_);
  and (_33388_, _33387_, _33357_);
  and (_33390_, _33330_, _02079_);
  or (_33391_, _33390_, _02158_);
  or (_33392_, _33391_, _33388_);
  nand (_33393_, _33392_, _33348_);
  nand (_33394_, _33393_, _10287_);
  nor (_33395_, _33330_, _10287_);
  nor (_33396_, _33395_, _02057_);
  nand (_33397_, _33396_, _33394_);
  and (_33398_, _04543_, _02057_);
  nor (_33399_, _33398_, _03446_);
  nand (_33401_, _33399_, _33397_);
  and (_33402_, _04458_, _03446_);
  nor (_33403_, _33402_, _02155_);
  nand (_33404_, _33403_, _33401_);
  and (_33405_, _04543_, _02155_);
  nor (_33406_, _33405_, _22169_);
  nand (_33407_, _33406_, _33404_);
  nor (_33408_, _33330_, _10452_);
  nor (_33409_, _33408_, _02153_);
  nand (_33410_, _33409_, _33407_);
  and (_33412_, _04543_, _02153_);
  nor (_33413_, _33412_, _10462_);
  nand (_33414_, _33413_, _33410_);
  nor (_33415_, _33330_, _10460_);
  nor (_33416_, _33415_, _02053_);
  nand (_33417_, _33416_, _33414_);
  and (_33418_, _04543_, _02053_);
  nor (_33419_, _33418_, _10464_);
  nand (_33420_, _33419_, _33417_);
  and (_33421_, _04458_, _10464_);
  nor (_33423_, _33421_, _02052_);
  nand (_33424_, _33423_, _33420_);
  and (_33425_, _04543_, _02052_);
  nor (_33426_, _33425_, _10475_);
  nand (_33427_, _33426_, _33424_);
  and (_33428_, _08770_, _05322_);
  not (_33429_, _33344_);
  nor (_33430_, _33429_, _08770_);
  or (_33431_, _33430_, _10471_);
  nor (_33432_, _33431_, _33428_);
  nor (_33434_, _33432_, _32347_);
  nand (_33435_, _33434_, _33427_);
  and (_33436_, _08877_, _05322_);
  nor (_33437_, _33429_, _08877_);
  nor (_33438_, _33437_, _33436_);
  nor (_33439_, _33438_, _02547_);
  or (_33440_, _10482_, _05323_);
  or (_33441_, _33429_, _08842_);
  nand (_33442_, _33441_, _33440_);
  and (_33443_, _33442_, _08790_);
  nor (_33445_, _33443_, _33439_);
  nand (_33446_, _33445_, _33435_);
  nand (_33447_, _33446_, _08917_);
  nand (_33448_, _08922_, _05322_);
  nand (_33449_, _33344_, _32011_);
  and (_33450_, _33449_, _33448_);
  or (_33451_, _33450_, _08917_);
  and (_33452_, _33451_, _33447_);
  or (_33453_, _33452_, _08881_);
  nand (_33454_, _33330_, _08881_);
  and (_33456_, _33454_, _33453_);
  nand (_33457_, _33456_, _02047_);
  and (_33458_, _04544_, _02046_);
  nor (_33459_, _33458_, _03310_);
  nand (_33460_, _33459_, _33457_);
  nor (_33461_, _04458_, _01750_);
  nor (_33462_, _33461_, _31256_);
  and (_33463_, _33462_, _33460_);
  or (_33464_, _33463_, _33339_);
  nand (_33465_, _33464_, _10158_);
  nor (_33467_, _33330_, _10158_);
  nor (_33468_, _33467_, _02182_);
  nand (_33469_, _33468_, _33465_);
  and (_33470_, _04543_, _02182_);
  nor (_33471_, _33470_, _10513_);
  nand (_33472_, _33471_, _33469_);
  and (_33473_, _04458_, _10513_);
  nor (_33474_, _33473_, _02181_);
  nand (_33475_, _33474_, _33472_);
  and (_33476_, _04543_, _02181_);
  nor (_33478_, _33476_, _10517_);
  and (_33479_, _33478_, _33475_);
  nor (_33480_, _33330_, _10153_);
  or (_33481_, _33480_, _33479_);
  nand (_33482_, _33481_, _07016_);
  nor (_33483_, _07016_, _04543_);
  nor (_33484_, _33483_, _01876_);
  and (_33485_, _33484_, _33482_);
  not (_33486_, _33330_);
  nor (_33487_, _33486_, _01778_);
  or (_33489_, _33487_, _02042_);
  nor (_33490_, _33489_, _33485_);
  and (_33491_, _04544_, _02042_);
  or (_33492_, _33491_, _33490_);
  nand (_33493_, _33492_, _04460_);
  and (_33494_, _04458_, _01767_);
  nor (_33495_, _33494_, _02218_);
  nand (_33496_, _33495_, _33493_);
  nand (_33497_, _33496_, _10534_);
  or (_33498_, _33497_, _33338_);
  nor (_33500_, _10534_, _04543_);
  nor (_33501_, _33500_, _01765_);
  nand (_33502_, _33501_, _33498_);
  and (_33503_, _05322_, _01765_);
  nor (_33504_, _33503_, _10546_);
  nand (_33505_, _33504_, _33502_);
  nor (_33506_, _33330_, _10542_);
  nor (_33507_, _33506_, _02124_);
  nand (_33508_, _33507_, _33505_);
  and (_33509_, _04543_, _02124_);
  nor (_33510_, _33509_, _01711_);
  nand (_33511_, _33510_, _33508_);
  and (_33512_, _04458_, _01711_);
  nor (_33513_, _33512_, _10550_);
  nand (_33514_, _33513_, _33511_);
  and (_33515_, _33353_, _10550_);
  nor (_33516_, _33515_, _04920_);
  and (_33517_, _33516_, _33514_);
  or (_33518_, _33517_, _33337_);
  nand (_33519_, _33518_, _01995_);
  and (_33521_, _05323_, _01994_);
  nor (_33522_, _33521_, _07239_);
  nand (_33523_, _33522_, _33519_);
  and (_33524_, _07239_, _04543_);
  nor (_33525_, _33524_, _10149_);
  nand (_33526_, _33525_, _33523_);
  or (_33527_, _10566_, _10567_);
  not (_33528_, _33527_);
  and (_33529_, _33528_, _10586_);
  nor (_33530_, _33528_, _10586_);
  nor (_33532_, _33530_, _33529_);
  and (_33533_, _33532_, _10149_);
  nor (_33534_, _33533_, _02123_);
  and (_33535_, _33534_, _33526_);
  and (_33536_, _04543_, _02123_);
  or (_33537_, _33536_, _01718_);
  or (_33538_, _33537_, _33535_);
  and (_33539_, _04458_, _01718_);
  nor (_33540_, _33539_, _10604_);
  nand (_33541_, _33540_, _33538_);
  nor (_33543_, _33353_, _07587_);
  and (_33544_, _07587_, _04544_);
  nor (_33545_, _33544_, _10605_);
  not (_33546_, _33545_);
  nor (_33547_, _33546_, _33543_);
  nor (_33548_, _33547_, _10609_);
  and (_33549_, _33548_, _33541_);
  or (_33550_, _33549_, _33336_);
  nand (_33551_, _33550_, _10618_);
  nor (_33552_, _10618_, _04543_);
  nor (_33554_, _33552_, _02210_);
  nand (_33555_, _33554_, _33551_);
  and (_33556_, _05322_, _02210_);
  nor (_33557_, _33556_, _02331_);
  and (_33558_, _33557_, _33555_);
  and (_33559_, _04544_, _02331_);
  or (_33560_, _33559_, _33558_);
  nand (_33561_, _33560_, _30883_);
  and (_33562_, _04458_, _01722_);
  nor (_33563_, _33562_, _10629_);
  nand (_33565_, _33563_, _33561_);
  and (_33566_, _10611_, _04543_);
  and (_33567_, _33353_, _07587_);
  or (_33568_, _33567_, _33566_);
  and (_33569_, _33568_, _10629_);
  nor (_33570_, _33569_, _10634_);
  and (_33571_, _33570_, _33565_);
  or (_33572_, _33571_, _33335_);
  nand (_33573_, _33572_, _10135_);
  nor (_33574_, _10135_, _04543_);
  nor (_33576_, _33574_, _02206_);
  nand (_33577_, _33576_, _33573_);
  and (_33578_, _05322_, _02206_);
  nor (_33579_, _33578_, _02342_);
  and (_33580_, _33579_, _33577_);
  and (_33581_, _04544_, _02342_);
  or (_33582_, _33581_, _33580_);
  nand (_33583_, _33582_, _30879_);
  and (_33584_, _04458_, _01728_);
  nor (_33585_, _33584_, _10649_);
  nand (_33587_, _33585_, _33583_);
  or (_33588_, _33353_, \oc8051_golden_model_1.PSW [7]);
  or (_33589_, _04543_, _06707_);
  and (_33590_, _33589_, _10649_);
  and (_33591_, _33590_, _33588_);
  nor (_33592_, _33591_, _10654_);
  and (_33593_, _33592_, _33587_);
  or (_33594_, _33593_, _33333_);
  nand (_33595_, _33594_, _07339_);
  nor (_33596_, _07339_, _04543_);
  nor (_33598_, _33596_, _02202_);
  and (_33599_, _33598_, _33595_);
  and (_33600_, _05322_, _02202_);
  or (_33601_, _33600_, _02334_);
  nor (_33602_, _33601_, _33599_);
  and (_33603_, _04544_, _02334_);
  or (_33604_, _33603_, _33602_);
  nand (_33605_, _33604_, _30876_);
  and (_33606_, _04458_, _01736_);
  nor (_33607_, _33606_, _10122_);
  nand (_33609_, _33607_, _33605_);
  and (_33610_, _04543_, _06707_);
  and (_33611_, _33353_, \oc8051_golden_model_1.PSW [7]);
  or (_33612_, _33611_, _33610_);
  and (_33613_, _33612_, _10122_);
  nor (_33614_, _33613_, _10671_);
  and (_33615_, _33614_, _33609_);
  or (_33616_, _33615_, _33332_);
  nand (_33617_, _33616_, _07385_);
  nor (_33618_, _07385_, _04543_);
  nor (_33620_, _33618_, _07415_);
  nand (_33621_, _33620_, _33617_);
  and (_33622_, _33330_, _07415_);
  nor (_33623_, _33622_, _02350_);
  and (_33624_, _33623_, _33621_);
  and (_33625_, _04698_, _02350_);
  or (_33626_, _33625_, _33624_);
  nand (_33627_, _33626_, _04964_);
  and (_33628_, _04458_, _01726_);
  nor (_33629_, _33628_, _02200_);
  nand (_33631_, _33629_, _33627_);
  and (_33632_, _33429_, _08690_);
  nor (_33633_, _08690_, _05322_);
  or (_33634_, _33633_, _10689_);
  nor (_33635_, _33634_, _33632_);
  nor (_33636_, _33635_, _10693_);
  and (_33637_, _33636_, _33631_);
  or (_33638_, _33637_, _33331_);
  nand (_33639_, _33638_, _07488_);
  nor (_33640_, _07488_, _04543_);
  nor (_33642_, _33640_, _07533_);
  nand (_33643_, _33642_, _33639_);
  and (_33644_, _33330_, _07533_);
  nor (_33645_, _33644_, _02083_);
  and (_33646_, _33645_, _33643_);
  and (_33647_, _04698_, _02083_);
  or (_33648_, _33647_, _33646_);
  nand (_33649_, _33648_, _10712_);
  and (_33650_, _04458_, _01738_);
  nor (_33651_, _33650_, _02243_);
  nand (_33653_, _33651_, _33649_);
  nor (_33654_, _33344_, _08690_);
  and (_33655_, _08690_, _05323_);
  nor (_33656_, _33655_, _33654_);
  and (_33657_, _33656_, _02243_);
  nor (_33658_, _33657_, _10723_);
  nand (_33659_, _33658_, _33653_);
  nor (_33660_, _33330_, _10722_);
  nor (_33661_, _33660_, _02366_);
  nand (_33662_, _33661_, _33659_);
  and (_33664_, _04543_, _02366_);
  nor (_33665_, _33664_, _31858_);
  and (_33666_, _33665_, _33662_);
  nor (_33667_, _33330_, _07581_);
  or (_33668_, _33667_, _33666_);
  nand (_33669_, _33668_, _01990_);
  and (_33670_, _04458_, _03537_);
  nor (_33671_, _33670_, _01697_);
  nand (_33672_, _33671_, _33669_);
  and (_33673_, _33656_, _01697_);
  nor (_33675_, _33673_, _10744_);
  nand (_33676_, _33675_, _33672_);
  and (_33677_, _33486_, _10744_);
  nor (_33678_, _33677_, _02081_);
  and (_33679_, _33678_, _33676_);
  or (_33680_, _33679_, _33328_);
  nand (_33681_, _33680_, _10751_);
  nor (_33682_, _33486_, _10751_);
  nor (_33683_, _33682_, _30863_);
  nand (_33684_, _33683_, _33681_);
  and (_33686_, _30863_, _04458_);
  nor (_33687_, _33686_, _10762_);
  nand (_33688_, _33687_, _33684_);
  and (_33689_, _33330_, _10762_);
  not (_33690_, _33689_);
  and (_33691_, _33690_, _33688_);
  nand (_33692_, _33691_, _39632_);
  or (_33693_, _39632_, \oc8051_golden_model_1.PC [7]);
  and (_33694_, _33693_, _39026_);
  and (_41800_, _33694_, _33692_);
  nor (_33696_, _10762_, _01732_);
  nor (_33697_, _10755_, _02027_);
  nor (_33698_, _05395_, _02027_);
  nor (_33699_, _10122_, _01736_);
  nor (_33700_, _10404_, _04919_);
  and (_33701_, _10404_, _02124_);
  and (_33702_, _10252_, _08877_);
  nor (_33703_, _10256_, _10250_);
  nor (_33704_, _33703_, _10257_);
  not (_33705_, _33704_);
  nor (_33707_, _33705_, _08877_);
  nor (_33708_, _33707_, _33702_);
  nor (_33709_, _33708_, _02547_);
  and (_33710_, _10252_, _08842_);
  and (_33711_, _33704_, _10482_);
  nor (_33712_, _33711_, _33710_);
  nor (_33713_, _33712_, _08836_);
  and (_33714_, _10404_, _02053_);
  and (_33715_, _10404_, _02057_);
  or (_33716_, _10295_, _10252_);
  or (_33718_, _33704_, _10293_);
  and (_33719_, _33718_, _33716_);
  or (_33720_, _33719_, _03006_);
  and (_33721_, _10435_, _10404_);
  nor (_33722_, _10407_, _10402_);
  nor (_33723_, _33722_, _10408_);
  and (_33724_, _33723_, _10437_);
  nor (_33725_, _33724_, _33721_);
  nand (_33726_, _33725_, _04535_);
  nor (_33727_, _10109_, \oc8051_golden_model_1.PC [8]);
  and (_33729_, _10109_, \oc8051_golden_model_1.PC [8]);
  nor (_33730_, _33729_, _33727_);
  nor (_33731_, _33730_, _06859_);
  nor (_33732_, _33730_, _10312_);
  nor (_33733_, _10301_, \oc8051_golden_model_1.PC [8]);
  nor (_33734_, _06855_, _02062_);
  and (_33735_, _33734_, _33733_);
  nor (_33736_, _33735_, _33732_);
  not (_33737_, _33736_);
  and (_33738_, _33737_, _10311_);
  nor (_33740_, _33738_, _33731_);
  nor (_33741_, _33740_, _02160_);
  nor (_33742_, _02160_, _02062_);
  nor (_33743_, _33742_, _10404_);
  nor (_33744_, _33743_, _06845_);
  not (_33745_, _33744_);
  nor (_33746_, _33745_, _33741_);
  not (_33747_, _33730_);
  and (_33748_, _33747_, _22054_);
  nor (_33749_, _33748_, _22055_);
  nor (_33751_, _33749_, _33746_);
  nor (_33752_, _33751_, _02079_);
  and (_33753_, _33752_, _33726_);
  and (_33754_, _33730_, _02079_);
  or (_33755_, _33754_, _02158_);
  or (_33756_, _33755_, _33753_);
  nand (_33757_, _33756_, _33720_);
  nand (_33758_, _33757_, _10287_);
  nor (_33759_, _33730_, _10287_);
  nor (_33760_, _33759_, _02057_);
  and (_33762_, _33760_, _33758_);
  or (_33763_, _33762_, _33715_);
  nand (_33764_, _33763_, _10446_);
  and (_33765_, _10404_, _02155_);
  nor (_33766_, _33765_, _22169_);
  nand (_33767_, _33766_, _33764_);
  nor (_33768_, _33730_, _10452_);
  nor (_33769_, _33768_, _02153_);
  nand (_33770_, _33769_, _33767_);
  and (_33771_, _10404_, _02153_);
  nor (_33773_, _33771_, _10462_);
  nand (_33774_, _33773_, _33770_);
  nor (_33775_, _33730_, _10460_);
  nor (_33776_, _33775_, _02053_);
  and (_33777_, _33776_, _33774_);
  or (_33778_, _33777_, _33714_);
  nand (_33779_, _33778_, _10465_);
  and (_33780_, _10404_, _02052_);
  nor (_33781_, _33780_, _10475_);
  nand (_33782_, _33781_, _33779_);
  and (_33783_, _10252_, _08770_);
  nor (_33784_, _33705_, _08770_);
  or (_33785_, _33784_, _10471_);
  nor (_33786_, _33785_, _33783_);
  nor (_33787_, _33786_, _32347_);
  and (_33788_, _33787_, _33782_);
  or (_33789_, _33788_, _33713_);
  or (_33790_, _33789_, _33709_);
  nand (_33791_, _33790_, _08917_);
  and (_33792_, _10253_, _08922_);
  nor (_33794_, _33704_, _08922_);
  or (_33795_, _33794_, _08917_);
  or (_33796_, _33795_, _33792_);
  and (_33797_, _33796_, _08882_);
  nand (_33798_, _33797_, _33791_);
  and (_33799_, _33747_, _08881_);
  nor (_33800_, _33799_, _02046_);
  nand (_33801_, _33800_, _33798_);
  and (_33802_, _10404_, _02046_);
  nor (_33803_, _33802_, _03310_);
  nand (_33805_, _33803_, _33801_);
  nand (_33806_, _33805_, _31255_);
  not (_33807_, _10404_);
  nor (_33808_, _31255_, _33807_);
  nor (_33809_, _33808_, _10159_);
  nand (_33810_, _33809_, _33806_);
  nor (_33811_, _33730_, _10158_);
  nor (_33812_, _33811_, _02182_);
  nand (_33813_, _33812_, _33810_);
  and (_33814_, _10404_, _02182_);
  nor (_33816_, _33814_, _10513_);
  nand (_33817_, _33816_, _33813_);
  nand (_33818_, _33817_, _09032_);
  and (_33819_, _10404_, _02181_);
  nor (_33820_, _33819_, _10517_);
  nand (_33821_, _33820_, _33818_);
  nor (_33822_, _33730_, _10153_);
  nor (_33823_, _33822_, _07017_);
  and (_33824_, _33823_, _33821_);
  nor (_33825_, _33807_, _07016_);
  or (_33827_, _33825_, _01876_);
  nor (_33828_, _33827_, _33824_);
  nor (_33829_, _33730_, _01778_);
  or (_33830_, _33829_, _33828_);
  nand (_33831_, _33830_, _02043_);
  and (_33832_, _33807_, _02042_);
  nor (_33833_, _33832_, _22431_);
  nand (_33834_, _33833_, _33831_);
  and (_33835_, _10252_, _02218_);
  not (_33836_, _33835_);
  and (_33838_, _33836_, _10534_);
  nand (_33839_, _33838_, _33834_);
  nor (_33840_, _10404_, _10534_);
  nor (_33841_, _33840_, _01765_);
  nand (_33842_, _33841_, _33839_);
  and (_33843_, _10252_, _01765_);
  nor (_33844_, _33843_, _10546_);
  nand (_33845_, _33844_, _33842_);
  nor (_33846_, _33730_, _10542_);
  nor (_33847_, _33846_, _02124_);
  and (_33849_, _33847_, _33845_);
  or (_33850_, _33849_, _33701_);
  nand (_33851_, _33850_, _22530_);
  and (_33852_, _33723_, _10550_);
  nor (_33853_, _33852_, _04920_);
  and (_33854_, _33853_, _33851_);
  or (_33855_, _33854_, _33700_);
  nand (_33856_, _33855_, _01995_);
  and (_33857_, _10253_, _01994_);
  nor (_33858_, _33857_, _07239_);
  nand (_33860_, _33858_, _33856_);
  and (_33861_, _10404_, _07239_);
  nor (_33862_, _33861_, _10149_);
  nand (_33863_, _33862_, _33860_);
  nor (_33864_, _10588_, \oc8051_golden_model_1.DPH [0]);
  nor (_33865_, _33864_, _10589_);
  nor (_33866_, _33865_, _10150_);
  nor (_33867_, _33866_, _02123_);
  nand (_33868_, _33867_, _33863_);
  and (_33869_, _10404_, _02123_);
  nor (_33871_, _33869_, _01718_);
  nand (_33872_, _33871_, _33868_);
  nand (_33873_, _33872_, _10605_);
  and (_33874_, _10404_, _07587_);
  and (_33875_, _33723_, _10611_);
  or (_33876_, _33875_, _33874_);
  and (_33877_, _33876_, _10604_);
  nor (_33878_, _33877_, _10609_);
  nand (_33879_, _33878_, _33873_);
  nor (_33880_, _33730_, _10147_);
  nor (_33882_, _33880_, _10619_);
  nand (_33883_, _33882_, _33879_);
  nor (_33884_, _10618_, _33807_);
  nor (_33885_, _33884_, _02210_);
  nand (_33886_, _33885_, _33883_);
  and (_33887_, _10253_, _02210_);
  nor (_33888_, _33887_, _02331_);
  nand (_33889_, _33888_, _33886_);
  and (_33890_, _10404_, _02331_);
  nor (_33891_, _33890_, _01722_);
  nand (_33893_, _33891_, _33889_);
  nand (_33894_, _33893_, _10630_);
  and (_33895_, _10404_, _10611_);
  and (_33896_, _33723_, _07587_);
  or (_33897_, _33896_, _33895_);
  and (_33898_, _33897_, _10629_);
  nor (_33899_, _33898_, _10634_);
  nand (_33900_, _33899_, _33894_);
  nor (_33901_, _33730_, _10139_);
  nor (_33902_, _33901_, _10136_);
  nand (_33904_, _33902_, _33900_);
  nor (_33905_, _33807_, _10135_);
  nor (_33906_, _33905_, _02206_);
  and (_33907_, _33906_, _33904_);
  and (_33908_, _10253_, _02206_);
  or (_33909_, _33908_, _33907_);
  nand (_33910_, _33909_, _03065_);
  nor (_33911_, _10649_, _01728_);
  not (_33912_, _33911_);
  and (_33913_, _33807_, _02342_);
  nor (_33915_, _33913_, _33912_);
  nand (_33916_, _33915_, _33910_);
  or (_33917_, _33723_, \oc8051_golden_model_1.PSW [7]);
  or (_33918_, _10404_, _06707_);
  and (_33919_, _33918_, _10649_);
  and (_33920_, _33919_, _33917_);
  nor (_33921_, _33920_, _10654_);
  nand (_33922_, _33921_, _33916_);
  nor (_33923_, _33730_, _10133_);
  nor (_33924_, _33923_, _07340_);
  and (_33926_, _33924_, _33922_);
  nor (_33927_, _33807_, _07339_);
  or (_33928_, _33927_, _02202_);
  or (_33929_, _33928_, _33926_);
  and (_33930_, _10253_, _02202_);
  nor (_33931_, _33930_, _02334_);
  and (_33932_, _33931_, _33929_);
  and (_33933_, _10404_, _02334_);
  or (_33934_, _33933_, _33932_);
  nand (_33935_, _33934_, _33699_);
  and (_33937_, _10404_, _06707_);
  and (_33938_, _33723_, \oc8051_golden_model_1.PSW [7]);
  or (_33939_, _33938_, _33937_);
  and (_33940_, _33939_, _10122_);
  nor (_33941_, _33940_, _10671_);
  nand (_33942_, _33941_, _33935_);
  nor (_33943_, _33730_, _10120_);
  nor (_33944_, _33943_, _07386_);
  nand (_33945_, _33944_, _33942_);
  nor (_33946_, _33807_, _07385_);
  nor (_33947_, _33946_, _07415_);
  nand (_33948_, _33947_, _33945_);
  and (_33949_, _33747_, _07415_);
  nor (_33950_, _33949_, _02350_);
  nand (_33951_, _33950_, _33948_);
  and (_33952_, _03002_, _02350_);
  nor (_33953_, _33952_, _01726_);
  nand (_33954_, _33953_, _33951_);
  nand (_33955_, _33954_, _10689_);
  and (_33956_, _33705_, _08690_);
  nor (_33958_, _10252_, _08690_);
  or (_33959_, _33958_, _10689_);
  nor (_33960_, _33959_, _33956_);
  nor (_33961_, _33960_, _10693_);
  nand (_33962_, _33961_, _33955_);
  nor (_33963_, _33730_, _10118_);
  nor (_33964_, _33963_, _07489_);
  nand (_33965_, _33964_, _33962_);
  nor (_33966_, _33807_, _07488_);
  nor (_33967_, _33966_, _07533_);
  nand (_33969_, _33967_, _33965_);
  and (_33970_, _33747_, _07533_);
  nor (_33971_, _33970_, _02083_);
  nand (_33972_, _33971_, _33969_);
  and (_33973_, _03002_, _02083_);
  nor (_33974_, _33973_, _01738_);
  nand (_33975_, _33974_, _33972_);
  nand (_33976_, _33975_, _02367_);
  and (_33977_, _10253_, _08690_);
  nor (_33978_, _33704_, _08690_);
  nor (_33980_, _33978_, _33977_);
  and (_33981_, _33980_, _02243_);
  nor (_33982_, _33981_, _10723_);
  nand (_33983_, _33982_, _33976_);
  nor (_33984_, _33730_, _10722_);
  nor (_33985_, _33984_, _02366_);
  nand (_33986_, _33985_, _33983_);
  and (_33987_, _10404_, _02366_);
  nor (_33988_, _33987_, _31858_);
  nand (_33989_, _33988_, _33986_);
  nor (_33991_, _33730_, _07581_);
  nor (_33992_, _33991_, _01989_);
  and (_33993_, _33992_, _33989_);
  or (_33994_, _33993_, _33698_);
  nor (_33995_, _01733_, _01697_);
  nand (_33996_, _33995_, _33994_);
  and (_33997_, _33980_, _01697_);
  nor (_33998_, _33997_, _10744_);
  nand (_33999_, _33998_, _33996_);
  and (_34000_, _33747_, _10744_);
  nor (_34002_, _34000_, _02081_);
  nand (_34003_, _34002_, _33999_);
  and (_34004_, _10404_, _02081_);
  nor (_34005_, _34004_, _31497_);
  nand (_34006_, _34005_, _34003_);
  nor (_34007_, _33730_, _10751_);
  nor (_34008_, _34007_, _02198_);
  and (_34009_, _34008_, _34006_);
  or (_34010_, _34009_, _33697_);
  nand (_34011_, _34010_, _33696_);
  and (_34013_, _33730_, _10762_);
  not (_34014_, _34013_);
  and (_34015_, _34014_, _34011_);
  nand (_34016_, _34015_, _39632_);
  or (_34017_, _39632_, \oc8051_golden_model_1.PC [8]);
  and (_34018_, _34017_, _39026_);
  and (_41802_, _34018_, _34016_);
  nor (_34019_, _02859_, _10755_);
  nor (_34020_, _02859_, _05395_);
  not (_34021_, \oc8051_golden_model_1.PC [9]);
  and (_34023_, _05320_, _10107_);
  and (_34024_, _34023_, \oc8051_golden_model_1.PC [8]);
  nor (_34025_, _34024_, _34021_);
  and (_34026_, _34024_, _34021_);
  or (_34027_, _34026_, _34025_);
  nor (_34028_, _34027_, _10118_);
  nor (_34029_, _34027_, _10120_);
  and (_34030_, _10192_, _02202_);
  nor (_34031_, _34027_, _10133_);
  and (_34032_, _10192_, _02206_);
  nor (_34034_, _34027_, _10139_);
  and (_34035_, _10192_, _02210_);
  nor (_34036_, _34027_, _10147_);
  nor (_34037_, _10352_, _04919_);
  and (_34038_, _10352_, _02124_);
  and (_34039_, _10352_, _02181_);
  nor (_34040_, _34027_, _10158_);
  not (_34041_, _34027_);
  and (_34042_, _34041_, _08881_);
  and (_34043_, _10352_, _02155_);
  and (_34045_, _10312_, _06859_);
  nor (_34046_, _34045_, _34027_);
  nor (_34047_, _10301_, \oc8051_golden_model_1.PC [9]);
  and (_34048_, _34047_, _33734_);
  and (_34049_, _34048_, _10311_);
  nor (_34050_, _34049_, _34046_);
  nor (_34051_, _34050_, _02160_);
  nor (_34052_, _33742_, _10352_);
  nor (_34053_, _34052_, _06845_);
  not (_34054_, _34053_);
  nor (_34056_, _34054_, _34051_);
  and (_34057_, _34027_, _06845_);
  not (_34058_, _34057_);
  and (_34059_, _34058_, _22054_);
  not (_34060_, _34059_);
  nor (_34061_, _34060_, _34056_);
  nor (_34062_, _10408_, _10405_);
  and (_34063_, _34062_, _10355_);
  nor (_34064_, _34062_, _10355_);
  nor (_34065_, _34064_, _34063_);
  nor (_34067_, _34065_, _10435_);
  and (_34068_, _10435_, _10352_);
  or (_34069_, _34068_, _34067_);
  nor (_34070_, _34069_, _04534_);
  nor (_34071_, _34070_, _34061_);
  nor (_34072_, _34071_, _02079_);
  and (_34073_, _34041_, _02079_);
  nor (_34074_, _34073_, _34072_);
  and (_34075_, _34074_, _03006_);
  nor (_34076_, _10257_, _10254_);
  and (_34077_, _34076_, _10196_);
  nor (_34078_, _34076_, _10196_);
  nor (_34079_, _34078_, _34077_);
  and (_34080_, _34079_, _10295_);
  nor (_34081_, _30930_, _10192_);
  or (_34082_, _34081_, _03006_);
  nor (_34083_, _34082_, _34080_);
  or (_34084_, _34083_, _10288_);
  nor (_34085_, _34084_, _34075_);
  nor (_34086_, _34027_, _10287_);
  nor (_34088_, _34086_, _02057_);
  not (_34089_, _34088_);
  nor (_34090_, _34089_, _34085_);
  and (_34091_, _10352_, _02057_);
  or (_34092_, _34091_, _03446_);
  nor (_34093_, _34092_, _34090_);
  nor (_34094_, _34093_, _02155_);
  or (_34095_, _34094_, _22169_);
  or (_34096_, _34095_, _34043_);
  nor (_34097_, _34027_, _10452_);
  nor (_34099_, _34097_, _02153_);
  nand (_34100_, _34099_, _34096_);
  and (_34101_, _10352_, _02153_);
  nor (_34102_, _34101_, _10462_);
  nand (_34103_, _34102_, _34100_);
  nor (_34104_, _34027_, _10460_);
  nor (_34105_, _34104_, _02053_);
  nand (_34106_, _34105_, _34103_);
  and (_34107_, _10352_, _02053_);
  nor (_34108_, _34107_, _10464_);
  nand (_34110_, _34108_, _34106_);
  nand (_34111_, _34110_, _03114_);
  and (_34112_, _10352_, _02052_);
  nor (_34113_, _34112_, _10475_);
  nand (_34114_, _34113_, _34111_);
  and (_34115_, _10192_, _08770_);
  nor (_34116_, _34079_, _08770_);
  or (_34117_, _34116_, _10471_);
  nor (_34118_, _34117_, _34115_);
  nor (_34119_, _34118_, _32347_);
  nand (_34121_, _34119_, _34114_);
  nor (_34122_, _34079_, _08877_);
  and (_34123_, _10192_, _08877_);
  nor (_34124_, _34123_, _34122_);
  nor (_34125_, _34124_, _02547_);
  not (_34126_, _34079_);
  and (_34127_, _34126_, _10482_);
  and (_34128_, _10192_, _08842_);
  nor (_34129_, _34128_, _34127_);
  nor (_34130_, _34129_, _08836_);
  nor (_34132_, _34130_, _34125_);
  nand (_34133_, _34132_, _34121_);
  nand (_34134_, _34133_, _08917_);
  and (_34135_, _10192_, _08922_);
  nor (_34136_, _34079_, _08922_);
  or (_34137_, _34136_, _34135_);
  and (_34138_, _34137_, _02246_);
  nor (_34139_, _34138_, _08881_);
  and (_34140_, _34139_, _34134_);
  or (_34141_, _34140_, _34042_);
  nand (_34143_, _34141_, _02047_);
  not (_34144_, _10352_);
  and (_34145_, _34144_, _02046_);
  nand (_34146_, _31252_, _22230_);
  nor (_34147_, _34146_, _34145_);
  nand (_34148_, _34147_, _34143_);
  nor (_34149_, _31255_, _34144_);
  nor (_34150_, _34149_, _10159_);
  and (_34151_, _34150_, _34148_);
  or (_34152_, _34151_, _34040_);
  nand (_34154_, _34152_, _08505_);
  and (_34155_, _34144_, _02182_);
  not (_34156_, _34155_);
  and (_34157_, _34156_, _10514_);
  and (_34158_, _34157_, _34154_);
  or (_34159_, _34158_, _34039_);
  nand (_34160_, _34159_, _10153_);
  nor (_34161_, _34041_, _10153_);
  nor (_34162_, _34161_, _07017_);
  nand (_34163_, _34162_, _34160_);
  nor (_34165_, _10352_, _07016_);
  nor (_34166_, _34165_, _01876_);
  nand (_34167_, _34166_, _34163_);
  nor (_34168_, _34041_, _01778_);
  nor (_34169_, _34168_, _02042_);
  nand (_34170_, _34169_, _34167_);
  and (_34171_, _34144_, _02042_);
  nor (_34172_, _34171_, _22431_);
  nand (_34173_, _34172_, _34170_);
  and (_34174_, _10192_, _02218_);
  not (_34176_, _34174_);
  and (_34177_, _34176_, _10534_);
  nand (_34178_, _34177_, _34173_);
  nor (_34179_, _10352_, _10534_);
  nor (_34180_, _34179_, _01765_);
  nand (_34181_, _34180_, _34178_);
  and (_34182_, _10192_, _01765_);
  nor (_34183_, _34182_, _10546_);
  nand (_34184_, _34183_, _34181_);
  nor (_34185_, _34027_, _10542_);
  nor (_34187_, _34185_, _02124_);
  and (_34188_, _34187_, _34184_);
  or (_34189_, _34188_, _34038_);
  nand (_34190_, _34189_, _22530_);
  nor (_34191_, _34065_, _10551_);
  nor (_34192_, _34191_, _04920_);
  and (_34193_, _34192_, _34190_);
  or (_34194_, _34193_, _34037_);
  nand (_34195_, _34194_, _01995_);
  and (_34196_, _10193_, _01994_);
  nor (_34197_, _34196_, _07239_);
  nand (_34198_, _34197_, _34195_);
  and (_34199_, _10352_, _07239_);
  nor (_34200_, _34199_, _10149_);
  nand (_34201_, _34200_, _34198_);
  nor (_34202_, _10589_, \oc8051_golden_model_1.DPH [1]);
  nor (_34203_, _34202_, _10590_);
  nor (_34204_, _34203_, _10150_);
  nor (_34205_, _34204_, _02123_);
  nand (_34206_, _34205_, _34201_);
  and (_34208_, _10352_, _02123_);
  nor (_34209_, _34208_, _01718_);
  nand (_34210_, _34209_, _34206_);
  nand (_34211_, _34210_, _10605_);
  and (_34212_, _34065_, _10611_);
  nor (_34213_, _10352_, _10611_);
  nor (_34214_, _34213_, _10605_);
  not (_34215_, _34214_);
  nor (_34216_, _34215_, _34212_);
  nor (_34217_, _34216_, _10609_);
  and (_34219_, _34217_, _34211_);
  or (_34220_, _34219_, _34036_);
  nand (_34221_, _34220_, _10618_);
  nor (_34222_, _10618_, _10352_);
  nor (_34223_, _34222_, _02210_);
  and (_34224_, _34223_, _34221_);
  or (_34225_, _34224_, _34035_);
  nand (_34226_, _34225_, _03061_);
  and (_34227_, _10352_, _02331_);
  nor (_34228_, _34227_, _01722_);
  nand (_34230_, _34228_, _34226_);
  nand (_34231_, _34230_, _10630_);
  and (_34232_, _34065_, _07587_);
  nor (_34233_, _10352_, _07587_);
  nor (_34234_, _34233_, _10630_);
  not (_34235_, _34234_);
  nor (_34236_, _34235_, _34232_);
  nor (_34237_, _34236_, _10634_);
  and (_34238_, _34237_, _34231_);
  or (_34239_, _34238_, _34034_);
  nand (_34241_, _34239_, _10135_);
  nor (_34242_, _10352_, _10135_);
  nor (_34243_, _34242_, _02206_);
  and (_34244_, _34243_, _34241_);
  or (_34245_, _34244_, _34032_);
  nand (_34246_, _34245_, _03065_);
  and (_34247_, _10352_, _02342_);
  nor (_34248_, _34247_, _01728_);
  nand (_34249_, _34248_, _34246_);
  nand (_34250_, _34249_, _10650_);
  nand (_34252_, _34065_, _06707_);
  or (_34253_, _10352_, _06707_);
  and (_34254_, _34253_, _10649_);
  and (_34255_, _34254_, _34252_);
  nor (_34256_, _34255_, _10654_);
  and (_34257_, _34256_, _34250_);
  or (_34258_, _34257_, _34031_);
  nand (_34259_, _34258_, _07339_);
  nor (_34260_, _10352_, _07339_);
  nor (_34261_, _34260_, _02202_);
  and (_34263_, _34261_, _34259_);
  or (_34264_, _34263_, _34030_);
  nand (_34265_, _34264_, _04958_);
  and (_34266_, _10352_, _02334_);
  nor (_34267_, _34266_, _01736_);
  nand (_34268_, _34267_, _34265_);
  nand (_34269_, _34268_, _10123_);
  and (_34270_, _10352_, _06707_);
  nor (_34271_, _34065_, _06707_);
  or (_34272_, _34271_, _34270_);
  and (_34274_, _34272_, _10122_);
  nor (_34275_, _34274_, _10671_);
  and (_34276_, _34275_, _34269_);
  or (_34277_, _34276_, _34029_);
  nand (_34278_, _34277_, _07385_);
  nor (_34279_, _10352_, _07385_);
  nor (_34280_, _34279_, _07415_);
  nand (_34281_, _34280_, _34278_);
  and (_34282_, _34027_, _07415_);
  nor (_34283_, _34282_, _02350_);
  nand (_34285_, _34283_, _34281_);
  nor (_34286_, _02200_, _01726_);
  not (_34287_, _34286_);
  and (_34288_, _03161_, _02350_);
  nor (_34289_, _34288_, _34287_);
  nand (_34290_, _34289_, _34285_);
  nor (_34291_, _10192_, _08690_);
  and (_34292_, _34079_, _08690_);
  or (_34293_, _34292_, _10689_);
  or (_34294_, _34293_, _34291_);
  and (_34295_, _34294_, _10118_);
  and (_34296_, _34295_, _34290_);
  or (_34297_, _34296_, _34028_);
  nand (_34298_, _34297_, _07488_);
  nor (_34299_, _10352_, _07488_);
  nor (_34300_, _34299_, _07533_);
  nand (_34301_, _34300_, _34298_);
  and (_34302_, _34027_, _07533_);
  nor (_34303_, _34302_, _02083_);
  nand (_34304_, _34303_, _34301_);
  and (_34306_, _03161_, _02083_);
  or (_34307_, _02243_, _01738_);
  nor (_34308_, _34307_, _34306_);
  nand (_34309_, _34308_, _34304_);
  and (_34310_, _10193_, _08690_);
  nor (_34311_, _34126_, _08690_);
  nor (_34312_, _34311_, _34310_);
  and (_34313_, _34312_, _02243_);
  nor (_34314_, _34313_, _10723_);
  nand (_34315_, _34314_, _34309_);
  nor (_34317_, _34027_, _10722_);
  nor (_34318_, _34317_, _02366_);
  nand (_34319_, _34318_, _34315_);
  and (_34320_, _10352_, _02366_);
  nor (_34321_, _34320_, _31858_);
  nand (_34322_, _34321_, _34319_);
  nor (_34323_, _34027_, _07581_);
  nor (_34324_, _34323_, _01989_);
  and (_34325_, _34324_, _34322_);
  or (_34326_, _34325_, _34020_);
  nand (_34328_, _34326_, _33995_);
  and (_34329_, _34312_, _01697_);
  nor (_34330_, _34329_, _10744_);
  nand (_34331_, _34330_, _34328_);
  and (_34332_, _34041_, _10744_);
  nor (_34333_, _34332_, _02081_);
  nand (_34334_, _34333_, _34331_);
  and (_34335_, _10352_, _02081_);
  nor (_34336_, _34335_, _31497_);
  nand (_34337_, _34336_, _34334_);
  nor (_34339_, _34027_, _10751_);
  nor (_34340_, _34339_, _02198_);
  and (_34341_, _34340_, _34337_);
  or (_34342_, _34341_, _34019_);
  nand (_34343_, _34342_, _33696_);
  and (_34344_, _34027_, _10762_);
  not (_34345_, _34344_);
  and (_34346_, _34345_, _34343_);
  nand (_34347_, _34346_, _39632_);
  or (_34348_, _39632_, \oc8051_golden_model_1.PC [9]);
  and (_34350_, _34348_, _39026_);
  and (_41803_, _34350_, _34347_);
  and (_34351_, _32974_, \oc8051_golden_model_1.PC [7]);
  and (_34352_, _34351_, \oc8051_golden_model_1.PC [8]);
  and (_34353_, _34352_, \oc8051_golden_model_1.PC [9]);
  and (_34354_, _34353_, \oc8051_golden_model_1.PC [10]);
  nor (_34355_, _34353_, \oc8051_golden_model_1.PC [10]);
  nor (_34356_, _34355_, _34354_);
  and (_34357_, _34356_, _10762_);
  not (_34358_, _34357_);
  and (_34360_, _02452_, _02198_);
  not (_34361_, _34356_);
  and (_34362_, _34361_, _10744_);
  and (_34363_, _02452_, _01989_);
  nor (_34364_, _34356_, _10722_);
  and (_34365_, _34361_, _07533_);
  and (_34366_, _34361_, _07415_);
  and (_34367_, _10186_, _02202_);
  and (_34368_, _10186_, _02206_);
  and (_34369_, _10186_, _02210_);
  nor (_34371_, _10604_, _01718_);
  nor (_34372_, _34361_, _10460_);
  not (_34373_, _10189_);
  nor (_34374_, _10261_, _10258_);
  nor (_34375_, _34374_, _34373_);
  and (_34376_, _34374_, _34373_);
  nor (_34377_, _34376_, _34375_);
  or (_34378_, _34377_, _10293_);
  or (_34379_, _10295_, _10185_);
  and (_34380_, _34379_, _34378_);
  nor (_34382_, _34380_, _03006_);
  not (_34383_, _10349_);
  nor (_34384_, _10412_, _10409_);
  nor (_34385_, _34384_, _34383_);
  and (_34386_, _34384_, _34383_);
  nor (_34387_, _34386_, _34385_);
  and (_34388_, _34387_, _10437_);
  and (_34389_, _10435_, _10346_);
  nor (_34390_, _34389_, _34388_);
  nand (_34391_, _34390_, _04535_);
  nor (_34392_, _34356_, _34045_);
  not (_34393_, _10346_);
  and (_34394_, _34393_, _02062_);
  nor (_34395_, _02062_, \oc8051_golden_model_1.PC [10]);
  and (_34396_, _34395_, _10302_);
  nor (_34397_, _34396_, _34394_);
  nor (_34398_, _34397_, _06855_);
  and (_34399_, _34398_, _10311_);
  nor (_34400_, _34399_, _34392_);
  and (_34401_, _34400_, _06847_);
  and (_34403_, _10346_, _02160_);
  or (_34404_, _34403_, _34401_);
  and (_34405_, _34404_, _10299_);
  and (_34406_, _34356_, _06845_);
  not (_34407_, _34406_);
  and (_34408_, _34407_, _22054_);
  not (_34409_, _34408_);
  nor (_34410_, _34409_, _34405_);
  nor (_34411_, _34410_, _02079_);
  nand (_34412_, _34411_, _34391_);
  and (_34414_, _34356_, _02079_);
  nor (_34415_, _34414_, _02158_);
  and (_34416_, _34415_, _34412_);
  or (_34417_, _34416_, _34382_);
  nand (_34418_, _34417_, _10287_);
  nor (_34419_, _34356_, _10287_);
  nor (_34420_, _34419_, _02057_);
  nand (_34421_, _34420_, _34418_);
  and (_34422_, _10346_, _02057_);
  not (_34423_, _34422_);
  and (_34425_, _34423_, _10446_);
  and (_34426_, _34425_, _34421_);
  and (_34427_, _34393_, _02155_);
  or (_34428_, _34427_, _34426_);
  and (_34429_, _34428_, _10452_);
  nor (_34430_, _34356_, _10452_);
  or (_34431_, _34430_, _34429_);
  nand (_34432_, _34431_, _02549_);
  and (_34433_, _34393_, _02153_);
  nor (_34434_, _34433_, _10462_);
  and (_34436_, _34434_, _34432_);
  or (_34437_, _34436_, _34372_);
  nand (_34438_, _34437_, _02054_);
  and (_34439_, _10346_, _02053_);
  nor (_34440_, _34439_, _10464_);
  nand (_34441_, _34440_, _34438_);
  nand (_34442_, _34441_, _03114_);
  and (_34443_, _10346_, _02052_);
  nor (_34444_, _34443_, _10475_);
  nand (_34445_, _34444_, _34442_);
  and (_34447_, _10185_, _08770_);
  not (_34448_, _34377_);
  nor (_34449_, _34448_, _08770_);
  or (_34450_, _34449_, _10471_);
  nor (_34451_, _34450_, _34447_);
  nor (_34452_, _34451_, _32347_);
  nand (_34453_, _34452_, _34445_);
  nor (_34454_, _34448_, _08877_);
  and (_34455_, _10185_, _08877_);
  nor (_34456_, _34455_, _34454_);
  nor (_34458_, _34456_, _02547_);
  or (_34459_, _34448_, _08842_);
  or (_34460_, _10186_, _10482_);
  nand (_34461_, _34460_, _34459_);
  and (_34462_, _34461_, _08790_);
  nor (_34463_, _34462_, _34458_);
  nand (_34464_, _34463_, _34453_);
  nand (_34465_, _34464_, _08917_);
  and (_34466_, _10185_, _08922_);
  and (_34467_, _34377_, _32011_);
  or (_34469_, _34467_, _34466_);
  and (_34470_, _34469_, _02246_);
  nor (_34471_, _34470_, _08881_);
  nand (_34472_, _34471_, _34465_);
  and (_34473_, _34361_, _08881_);
  not (_34474_, _34473_);
  and (_34475_, _31254_, _02148_);
  and (_34476_, _34475_, _34474_);
  and (_34477_, _34476_, _34472_);
  nor (_34478_, _34475_, _34393_);
  nor (_34480_, _34478_, _10159_);
  nand (_34481_, _34480_, _01750_);
  or (_34482_, _34481_, _34477_);
  nor (_34483_, _34356_, _10158_);
  nor (_34484_, _34483_, _02182_);
  nand (_34485_, _34484_, _34482_);
  nand (_34486_, _34485_, _01755_);
  nand (_34487_, _34486_, _09032_);
  nor (_34488_, _34393_, _02183_);
  nor (_34489_, _34488_, _10517_);
  nand (_34491_, _34489_, _34487_);
  nor (_34492_, _34356_, _10153_);
  nor (_34493_, _34492_, _07017_);
  nand (_34494_, _34493_, _34491_);
  nor (_34495_, _34393_, _07016_);
  nor (_34496_, _34495_, _01876_);
  nand (_34497_, _34496_, _34494_);
  nor (_34498_, _34356_, _01778_);
  nor (_34499_, _34498_, _02042_);
  and (_34500_, _34499_, _34497_);
  and (_34502_, _10346_, _02042_);
  nor (_34503_, _34502_, _34500_);
  and (_34504_, _34503_, _22430_);
  and (_34505_, _10186_, _02218_);
  or (_34506_, _34505_, _34504_);
  and (_34507_, _34506_, _10534_);
  nor (_34508_, _10346_, _10534_);
  or (_34509_, _34508_, _34507_);
  nand (_34510_, _34509_, _02037_);
  and (_34511_, _10186_, _01765_);
  nor (_34513_, _34511_, _10546_);
  and (_34514_, _34513_, _34510_);
  nor (_34515_, _34361_, _10542_);
  or (_34516_, _34515_, _34514_);
  nand (_34517_, _34516_, _31521_);
  and (_34518_, _10346_, _02124_);
  not (_34519_, _34518_);
  and (_34520_, _34519_, _22530_);
  nand (_34521_, _34520_, _34517_);
  nor (_34522_, _34387_, _10551_);
  nor (_34524_, _34522_, _04920_);
  and (_34525_, _34524_, _34521_);
  nor (_34526_, _34393_, _04919_);
  or (_34527_, _34526_, _01994_);
  or (_34528_, _34527_, _34525_);
  and (_34529_, _10186_, _01994_);
  nor (_34530_, _34529_, _07239_);
  nand (_34531_, _34530_, _34528_);
  and (_34532_, _10346_, _07239_);
  nor (_34533_, _34532_, _10149_);
  nand (_34535_, _34533_, _34531_);
  nor (_34536_, _10590_, \oc8051_golden_model_1.DPH [2]);
  nor (_34537_, _34536_, _10591_);
  nor (_34538_, _34537_, _10150_);
  nor (_34539_, _34538_, _02123_);
  and (_34540_, _34539_, _34535_);
  and (_34541_, _10346_, _02123_);
  or (_34542_, _34541_, _34540_);
  nand (_34543_, _34542_, _34371_);
  and (_34544_, _10346_, _07587_);
  and (_34546_, _34387_, _10611_);
  or (_34547_, _34546_, _34544_);
  and (_34548_, _34547_, _10604_);
  nor (_34549_, _34548_, _10609_);
  nand (_34550_, _34549_, _34543_);
  nor (_34551_, _34356_, _10147_);
  nor (_34552_, _34551_, _10619_);
  nand (_34553_, _34552_, _34550_);
  nor (_34554_, _10618_, _34393_);
  nor (_34555_, _34554_, _02210_);
  and (_34557_, _34555_, _34553_);
  or (_34558_, _34557_, _34369_);
  nand (_34559_, _34558_, _03061_);
  and (_34560_, _34393_, _02331_);
  nor (_34561_, _34560_, _22715_);
  nand (_34562_, _34561_, _34559_);
  and (_34563_, _10346_, _10611_);
  and (_34564_, _34387_, _07587_);
  or (_34565_, _34564_, _34563_);
  and (_34566_, _34565_, _10629_);
  nor (_34568_, _34566_, _10634_);
  nand (_34569_, _34568_, _34562_);
  nor (_34570_, _34356_, _10139_);
  nor (_34571_, _34570_, _10136_);
  nand (_34572_, _34571_, _34569_);
  nor (_34573_, _34393_, _10135_);
  nor (_34574_, _34573_, _02206_);
  and (_34575_, _34574_, _34572_);
  or (_34576_, _34575_, _34368_);
  nand (_34577_, _34576_, _03065_);
  and (_34579_, _34393_, _02342_);
  nor (_34580_, _34579_, _33912_);
  nand (_34581_, _34580_, _34577_);
  or (_34582_, _34387_, \oc8051_golden_model_1.PSW [7]);
  or (_34583_, _10346_, _06707_);
  and (_34584_, _34583_, _10649_);
  and (_34585_, _34584_, _34582_);
  nor (_34586_, _34585_, _10654_);
  nand (_34587_, _34586_, _34581_);
  nor (_34588_, _34356_, _10133_);
  nor (_34590_, _34588_, _07340_);
  nand (_34591_, _34590_, _34587_);
  nor (_34592_, _34393_, _07339_);
  nor (_34593_, _34592_, _02202_);
  and (_34594_, _34593_, _34591_);
  or (_34595_, _34594_, _34367_);
  nand (_34596_, _34595_, _04958_);
  and (_34597_, _34393_, _02334_);
  not (_34598_, _34597_);
  and (_34599_, _34598_, _33699_);
  nand (_34601_, _34599_, _34596_);
  and (_34602_, _10346_, _06707_);
  and (_34603_, _34387_, \oc8051_golden_model_1.PSW [7]);
  or (_34604_, _34603_, _34602_);
  and (_34605_, _34604_, _10122_);
  nor (_34606_, _34605_, _10671_);
  nand (_34607_, _34606_, _34601_);
  nor (_34608_, _34356_, _10120_);
  nor (_34609_, _34608_, _07386_);
  nand (_34610_, _34609_, _34607_);
  nor (_34612_, _34393_, _07385_);
  nor (_34613_, _34612_, _07415_);
  and (_34614_, _34613_, _34610_);
  or (_34615_, _34614_, _34366_);
  nand (_34616_, _34615_, _09472_);
  and (_34617_, _03624_, _02350_);
  nor (_34618_, _34617_, _34287_);
  nand (_34619_, _34618_, _34616_);
  nor (_34620_, _10185_, _08690_);
  and (_34621_, _34448_, _08690_);
  or (_34622_, _34621_, _10689_);
  nor (_34623_, _34622_, _34620_);
  nor (_34624_, _34623_, _10693_);
  nand (_34625_, _34624_, _34619_);
  nor (_34626_, _34356_, _10118_);
  nor (_34627_, _34626_, _07489_);
  nand (_34628_, _34627_, _34625_);
  nor (_34629_, _34393_, _07488_);
  nor (_34630_, _34629_, _07533_);
  and (_34631_, _34630_, _34628_);
  or (_34633_, _34631_, _34365_);
  nand (_34634_, _34633_, _02084_);
  and (_34635_, _03624_, _02083_);
  nor (_34636_, _34635_, _34307_);
  nand (_34637_, _34636_, _34634_);
  nor (_34638_, _34377_, _08690_);
  and (_34639_, _10186_, _08690_);
  nor (_34640_, _34639_, _34638_);
  and (_34641_, _34640_, _02243_);
  nor (_34642_, _34641_, _10723_);
  and (_34644_, _34642_, _34637_);
  or (_34645_, _34644_, _34364_);
  nand (_34646_, _34645_, _02778_);
  and (_34647_, _34393_, _02366_);
  nor (_34648_, _34647_, _31858_);
  nand (_34649_, _34648_, _34646_);
  nor (_34650_, _34361_, _07581_);
  nor (_34651_, _34650_, _01989_);
  nand (_34652_, _34651_, _34649_);
  nand (_34653_, _34652_, _33995_);
  or (_34655_, _34653_, _34363_);
  and (_34656_, _34640_, _01697_);
  nor (_34657_, _34656_, _10744_);
  and (_34658_, _34657_, _34655_);
  or (_34659_, _34658_, _34362_);
  nand (_34660_, _34659_, _02082_);
  and (_34661_, _34393_, _02081_);
  nor (_34662_, _34661_, _31497_);
  nand (_34663_, _34662_, _34660_);
  nor (_34664_, _34361_, _10751_);
  nor (_34666_, _34664_, _02198_);
  nand (_34667_, _34666_, _34663_);
  nand (_34668_, _34667_, _33696_);
  or (_34669_, _34668_, _34360_);
  and (_34670_, _34669_, _34358_);
  nand (_34671_, _34670_, _39632_);
  or (_34672_, _39632_, \oc8051_golden_model_1.PC [10]);
  and (_34673_, _34672_, _39026_);
  and (_41804_, _34673_, _34671_);
  nand (_34674_, _03434_, _02083_);
  nor (_34676_, _10110_, _10176_);
  and (_34677_, _10110_, _10176_);
  or (_34678_, _34677_, _34676_);
  or (_34679_, _34678_, _10118_);
  or (_34680_, _34678_, _10120_);
  or (_34681_, _34678_, _10133_);
  or (_34682_, _34678_, _10139_);
  or (_34683_, _34678_, _10147_);
  or (_34684_, _10341_, _04919_);
  and (_34685_, _10179_, _01765_);
  or (_34686_, _34678_, _10153_);
  not (_34687_, _34678_);
  nor (_34688_, _34687_, _10158_);
  nand (_34689_, _10180_, _08877_);
  nor (_34690_, _34375_, _10187_);
  and (_34691_, _34690_, _10183_);
  nor (_34692_, _34690_, _10183_);
  or (_34693_, _34692_, _34691_);
  or (_34694_, _34693_, _08877_);
  and (_34695_, _34694_, _02171_);
  and (_34697_, _34695_, _34689_);
  nand (_34698_, _10180_, _08770_);
  or (_34699_, _34693_, _08770_);
  and (_34700_, _34699_, _10475_);
  and (_34701_, _34700_, _34698_);
  and (_34702_, _10341_, _02153_);
  or (_34703_, _10447_, _10341_);
  or (_34704_, _10295_, _10179_);
  or (_34705_, _34693_, _10293_);
  and (_34706_, _34705_, _02158_);
  and (_34708_, _34706_, _34704_);
  and (_34709_, _10435_, _10341_);
  nor (_34710_, _34385_, _10347_);
  nor (_34711_, _34710_, _10344_);
  and (_34712_, _34710_, _10344_);
  or (_34713_, _34712_, _34711_);
  and (_34714_, _34713_, _10437_);
  or (_34715_, _34714_, _04534_);
  or (_34716_, _34715_, _34709_);
  nand (_34717_, _34687_, _06845_);
  or (_34719_, _34678_, _34045_);
  nand (_34720_, _01747_, _10176_);
  nor (_34721_, _34720_, _02062_);
  and (_34722_, _34721_, _10312_);
  nand (_34723_, _34722_, _30897_);
  and (_34724_, _34723_, _34719_);
  or (_34725_, _34724_, _02160_);
  and (_34726_, _34725_, _34717_);
  or (_34727_, _34726_, _10323_);
  nor (_34728_, _10317_, _10323_);
  or (_34730_, _34728_, _10341_);
  and (_34731_, _34730_, _34727_);
  or (_34732_, _34731_, _04535_);
  and (_34733_, _34732_, _10442_);
  and (_34734_, _34733_, _34716_);
  or (_34735_, _34734_, _34708_);
  and (_34736_, _34735_, _10287_);
  not (_34737_, _10447_);
  nor (_34738_, _34687_, _10448_);
  or (_34739_, _34738_, _34737_);
  or (_34741_, _34739_, _34736_);
  and (_34742_, _34741_, _34703_);
  or (_34743_, _34742_, _22169_);
  or (_34744_, _34678_, _10452_);
  and (_34745_, _34744_, _02549_);
  and (_34746_, _34745_, _34743_);
  or (_34747_, _34746_, _34702_);
  and (_34748_, _34747_, _10460_);
  or (_34749_, _34687_, _10460_);
  nand (_34750_, _34749_, _10466_);
  or (_34751_, _34750_, _34748_);
  or (_34752_, _10466_, _10341_);
  and (_34753_, _34752_, _10471_);
  and (_34754_, _34753_, _34751_);
  or (_34755_, _34754_, _34701_);
  or (_34756_, _34755_, _08790_);
  and (_34757_, _10179_, _08842_);
  and (_34758_, _34693_, _10482_);
  or (_34759_, _34758_, _08836_);
  or (_34760_, _34759_, _34757_);
  and (_34761_, _34760_, _02547_);
  and (_34762_, _34761_, _34756_);
  or (_34763_, _34762_, _34697_);
  and (_34764_, _34763_, _08917_);
  or (_34765_, _34693_, _08922_);
  nand (_34766_, _10180_, _08922_);
  and (_34767_, _34766_, _02246_);
  and (_34768_, _34767_, _34765_);
  or (_34769_, _34768_, _34764_);
  and (_34770_, _34769_, _08882_);
  nand (_34772_, _34678_, _08881_);
  nand (_34773_, _34772_, _10506_);
  or (_34774_, _34773_, _34770_);
  or (_34775_, _10506_, _10341_);
  and (_34776_, _34775_, _10158_);
  and (_34777_, _34776_, _34774_);
  or (_34778_, _34777_, _34688_);
  and (_34779_, _34778_, _10515_);
  not (_34780_, _10515_);
  and (_34781_, _34780_, _10341_);
  or (_34783_, _34781_, _10517_);
  or (_34784_, _34783_, _34779_);
  and (_34785_, _34784_, _34686_);
  or (_34786_, _34785_, _07017_);
  or (_34787_, _10341_, _07016_);
  and (_34788_, _34787_, _01778_);
  and (_34789_, _34788_, _34786_);
  or (_34790_, _34687_, _01778_);
  nand (_34791_, _34790_, _10527_);
  or (_34792_, _34791_, _34789_);
  or (_34794_, _10527_, _10341_);
  and (_34795_, _34794_, _07633_);
  and (_34796_, _34795_, _34792_);
  nand (_34797_, _10179_, _02218_);
  nand (_34798_, _34797_, _10534_);
  or (_34799_, _34798_, _34796_);
  or (_34800_, _10341_, _10534_);
  and (_34801_, _34800_, _02037_);
  and (_34802_, _34801_, _34799_);
  or (_34803_, _34802_, _34685_);
  and (_34804_, _34803_, _10542_);
  nor (_34805_, _34687_, _10542_);
  or (_34806_, _34805_, _10545_);
  or (_34807_, _34806_, _34804_);
  or (_34808_, _10544_, _10341_);
  and (_34809_, _34808_, _10551_);
  and (_34810_, _34809_, _34807_);
  and (_34811_, _34713_, _10550_);
  or (_34812_, _34811_, _04920_);
  or (_34813_, _34812_, _34810_);
  and (_34815_, _34813_, _34684_);
  or (_34816_, _34815_, _01994_);
  nand (_34817_, _10180_, _01994_);
  and (_34818_, _34817_, _07240_);
  and (_34819_, _34818_, _34816_);
  and (_34820_, _10341_, _07239_);
  or (_34821_, _34820_, _34819_);
  and (_34822_, _34821_, _10150_);
  or (_34823_, _10591_, \oc8051_golden_model_1.DPH [3]);
  nor (_34824_, _10592_, _10150_);
  and (_34826_, _34824_, _34823_);
  or (_34827_, _34826_, _10601_);
  or (_34828_, _34827_, _34822_);
  or (_34829_, _10600_, _10341_);
  and (_34830_, _34829_, _10605_);
  and (_34831_, _34830_, _34828_);
  or (_34832_, _34713_, _07587_);
  or (_34833_, _10341_, _10611_);
  and (_34834_, _34833_, _10604_);
  and (_34835_, _34834_, _34832_);
  or (_34836_, _34835_, _10609_);
  or (_34837_, _34836_, _34831_);
  and (_34838_, _34837_, _34683_);
  or (_34839_, _34838_, _10619_);
  or (_34840_, _10618_, _10341_);
  and (_34841_, _34840_, _03059_);
  and (_34842_, _34841_, _34839_);
  nand (_34843_, _10179_, _02210_);
  nand (_34844_, _34843_, _10625_);
  or (_34845_, _34844_, _34842_);
  or (_34847_, _10625_, _10341_);
  and (_34848_, _34847_, _10630_);
  and (_34849_, _34848_, _34845_);
  or (_34850_, _34713_, _10611_);
  or (_34851_, _10341_, _07587_);
  and (_34852_, _34851_, _10629_);
  and (_34853_, _34852_, _34850_);
  or (_34854_, _34853_, _10634_);
  or (_34855_, _34854_, _34849_);
  and (_34856_, _34855_, _34682_);
  or (_34857_, _34856_, _10136_);
  or (_34858_, _10341_, _10135_);
  and (_34859_, _34858_, _02208_);
  and (_34860_, _34859_, _34857_);
  nand (_34861_, _10179_, _02206_);
  nand (_34862_, _34861_, _09561_);
  or (_34863_, _34862_, _34860_);
  and (_34864_, _10650_, _10341_);
  or (_34865_, _34864_, _22844_);
  and (_34866_, _34865_, _34863_);
  or (_34868_, _34713_, \oc8051_golden_model_1.PSW [7]);
  or (_34869_, _10341_, _06707_);
  and (_34870_, _34869_, _10649_);
  and (_34871_, _34870_, _34868_);
  or (_34872_, _34871_, _10654_);
  or (_34873_, _34872_, _34866_);
  and (_34874_, _34873_, _34681_);
  or (_34875_, _34874_, _07340_);
  or (_34876_, _10341_, _07339_);
  and (_34877_, _34876_, _04953_);
  and (_34879_, _34877_, _34875_);
  nand (_34880_, _10179_, _02202_);
  nand (_34881_, _34880_, _10124_);
  or (_34882_, _34881_, _34879_);
  and (_34883_, _10341_, _10123_);
  or (_34884_, _34883_, _22985_);
  and (_34885_, _34884_, _34882_);
  or (_34886_, _34713_, _06707_);
  or (_34887_, _10341_, \oc8051_golden_model_1.PSW [7]);
  and (_34888_, _34887_, _10122_);
  and (_34890_, _34888_, _34886_);
  or (_34891_, _34890_, _10671_);
  or (_34892_, _34891_, _34885_);
  and (_34893_, _34892_, _34680_);
  or (_34894_, _34893_, _07386_);
  or (_34895_, _10341_, _07385_);
  and (_34896_, _34895_, _07416_);
  and (_34897_, _34896_, _34894_);
  and (_34898_, _34678_, _07415_);
  or (_34899_, _34898_, _02350_);
  or (_34901_, _34899_, _34897_);
  nand (_34902_, _03434_, _02350_);
  and (_34903_, _34902_, _34901_);
  or (_34904_, _34903_, _01726_);
  or (_34905_, _10341_, _04964_);
  and (_34906_, _34905_, _10689_);
  and (_34907_, _34906_, _34904_);
  or (_34908_, _34693_, _10694_);
  or (_34909_, _10179_, _08690_);
  and (_34910_, _34909_, _02200_);
  and (_34912_, _34910_, _34908_);
  or (_34913_, _34912_, _10693_);
  or (_34914_, _34913_, _34907_);
  and (_34915_, _34914_, _34679_);
  or (_34916_, _34915_, _07489_);
  or (_34917_, _10341_, _07488_);
  and (_34918_, _34917_, _07534_);
  and (_34919_, _34918_, _34916_);
  and (_34920_, _34678_, _07533_);
  or (_34921_, _34920_, _02083_);
  or (_34923_, _34921_, _34919_);
  and (_34924_, _34923_, _34674_);
  or (_34925_, _34924_, _01738_);
  or (_34926_, _10341_, _10712_);
  and (_34927_, _34926_, _02367_);
  and (_34928_, _34927_, _34925_);
  or (_34929_, _34693_, _08690_);
  nand (_34930_, _10180_, _08690_);
  and (_34931_, _34930_, _34929_);
  and (_34932_, _34931_, _02243_);
  or (_34934_, _34932_, _10723_);
  or (_34935_, _34934_, _34928_);
  or (_34936_, _34678_, _10722_);
  and (_34937_, _34936_, _02778_);
  and (_34938_, _34937_, _34935_);
  nand (_34939_, _10341_, _02366_);
  nand (_34940_, _34939_, _07581_);
  or (_34941_, _34940_, _34938_);
  or (_34942_, _34678_, _07581_);
  and (_34943_, _34942_, _05395_);
  and (_34945_, _34943_, _34941_);
  nor (_34946_, _05395_, _01983_);
  or (_34947_, _34946_, _01733_);
  or (_34948_, _34947_, _34945_);
  or (_34949_, _10341_, _10738_);
  and (_34950_, _34949_, _01698_);
  and (_34951_, _34950_, _34948_);
  and (_34952_, _34931_, _01697_);
  or (_34953_, _34952_, _10744_);
  or (_34954_, _34953_, _34951_);
  nand (_34956_, _34687_, _10744_);
  and (_34957_, _34956_, _02082_);
  and (_34958_, _34957_, _34954_);
  nand (_34959_, _10341_, _02081_);
  nand (_34960_, _34959_, _10751_);
  or (_34961_, _34960_, _34958_);
  or (_34962_, _34678_, _10751_);
  and (_34963_, _34962_, _10755_);
  and (_34964_, _34963_, _34961_);
  nor (_34965_, _10755_, _01983_);
  or (_34967_, _34965_, _01732_);
  or (_34968_, _34967_, _34964_);
  or (_34969_, _10341_, _10764_);
  and (_34970_, _34969_, _10763_);
  and (_34971_, _34970_, _34968_);
  and (_34972_, _34678_, _10762_);
  or (_34973_, _34972_, _34971_);
  or (_34974_, _34973_, _39633_);
  or (_34975_, _39632_, \oc8051_golden_model_1.PC [11]);
  and (_34976_, _34975_, _39026_);
  and (_41805_, _34976_, _34974_);
  nor (_34978_, _10111_, \oc8051_golden_model_1.PC [12]);
  nor (_34979_, _34978_, _10112_);
  not (_34980_, _34979_);
  and (_34981_, _34980_, _07533_);
  not (_34982_, _10338_);
  nor (_34983_, _34982_, _10124_);
  nor (_34984_, _34982_, _09561_);
  nor (_34985_, _10625_, _34982_);
  nor (_34986_, _10600_, _34982_);
  and (_34988_, _10174_, _02218_);
  nor (_34989_, _34979_, _10452_);
  and (_34990_, _34979_, _02079_);
  and (_34991_, _10435_, _10338_);
  and (_34992_, _10419_, _10416_);
  nor (_34993_, _34992_, _10420_);
  and (_34994_, _34993_, _10437_);
  nor (_34995_, _34994_, _34991_);
  and (_34996_, _34995_, _04535_);
  and (_34997_, _34045_, _10299_);
  nor (_34999_, _34997_, _34980_);
  and (_35000_, _10338_, _10317_);
  nand (_35001_, _01747_, \oc8051_golden_model_1.PC [12]);
  nor (_35002_, _35001_, _02160_);
  and (_35003_, _33734_, _10302_);
  and (_35004_, _35003_, _35002_);
  and (_35005_, _35004_, _06859_);
  or (_35006_, _35005_, _35000_);
  and (_35007_, _35006_, _10299_);
  nor (_35008_, _35007_, _34999_);
  nor (_35010_, _35008_, _10323_);
  nor (_35011_, _34982_, _01752_);
  nor (_35012_, _35011_, _04535_);
  not (_35013_, _35012_);
  nor (_35014_, _35013_, _35010_);
  or (_35015_, _35014_, _02079_);
  nor (_35016_, _35015_, _34996_);
  or (_35017_, _35016_, _34990_);
  and (_35018_, _35017_, _03006_);
  and (_35019_, _10268_, _10265_);
  nor (_35021_, _35019_, _10269_);
  or (_35022_, _35021_, _10293_);
  or (_35023_, _10295_, _10173_);
  and (_35024_, _35023_, _35022_);
  and (_35025_, _35024_, _02158_);
  nor (_35026_, _35025_, _35018_);
  nand (_35027_, _35026_, _10287_);
  nor (_35028_, _34979_, _10287_);
  nor (_35029_, _35028_, _34737_);
  nand (_35030_, _35029_, _35027_);
  nor (_35032_, _10447_, _34982_);
  nor (_35033_, _35032_, _22169_);
  and (_35034_, _35033_, _35030_);
  or (_35035_, _35034_, _34989_);
  nand (_35036_, _35035_, _02549_);
  and (_35037_, _34982_, _02153_);
  nor (_35038_, _35037_, _10462_);
  and (_35039_, _35038_, _35036_);
  nor (_35040_, _34980_, _10460_);
  or (_35041_, _35040_, _35039_);
  nand (_35042_, _35041_, _10466_);
  nor (_35043_, _10466_, _34982_);
  nor (_35044_, _35043_, _10475_);
  and (_35045_, _35044_, _35042_);
  and (_35046_, _10173_, _08770_);
  not (_35047_, _35021_);
  nor (_35048_, _35047_, _08770_);
  or (_35049_, _35048_, _35046_);
  nor (_35050_, _35049_, _10471_);
  or (_35051_, _35050_, _35045_);
  nand (_35053_, _35051_, _08836_);
  or (_35054_, _35047_, _08842_);
  nand (_35055_, _10173_, _08842_);
  and (_35056_, _35055_, _08790_);
  nand (_35057_, _35056_, _35054_);
  and (_35058_, _35057_, _35053_);
  nand (_35059_, _35058_, _08692_);
  nor (_35060_, _35021_, _08922_);
  and (_35061_, _10174_, _08922_);
  nor (_35062_, _35061_, _08917_);
  not (_35064_, _35062_);
  nor (_35065_, _35064_, _35060_);
  nor (_35066_, _35065_, _08881_);
  nor (_35067_, _35021_, _08877_);
  and (_35068_, _10174_, _08877_);
  or (_35069_, _35068_, _02547_);
  or (_35070_, _35069_, _35067_);
  and (_35071_, _35070_, _35066_);
  and (_35072_, _35071_, _35059_);
  and (_35073_, _34980_, _08881_);
  or (_35075_, _35073_, _35072_);
  and (_35076_, _35075_, _10506_);
  nor (_35077_, _10506_, _10338_);
  or (_35078_, _35077_, _35076_);
  nand (_35079_, _35078_, _10158_);
  nor (_35080_, _34979_, _10158_);
  nor (_35081_, _35080_, _34780_);
  nand (_35082_, _35081_, _35079_);
  nor (_35083_, _10515_, _34982_);
  nor (_35084_, _35083_, _10517_);
  nand (_35086_, _35084_, _35082_);
  nor (_35087_, _34979_, _10153_);
  nor (_35088_, _35087_, _07017_);
  nand (_35089_, _35088_, _35086_);
  nor (_35090_, _34982_, _07016_);
  nor (_35091_, _35090_, _01876_);
  nand (_35092_, _35091_, _35089_);
  nor (_35093_, _34979_, _01778_);
  nor (_35094_, _35093_, _10528_);
  nand (_35095_, _35094_, _35092_);
  nor (_35097_, _10527_, _34982_);
  nor (_35098_, _35097_, _02218_);
  nand (_35099_, _35098_, _35095_);
  nand (_35100_, _35099_, _10534_);
  or (_35101_, _35100_, _34988_);
  nor (_35102_, _34982_, _10534_);
  nor (_35103_, _35102_, _01765_);
  nand (_35104_, _35103_, _35101_);
  and (_35105_, _10174_, _01765_);
  nor (_35106_, _35105_, _10546_);
  nand (_35108_, _35106_, _35104_);
  nor (_35109_, _34980_, _10542_);
  nor (_35110_, _35109_, _10545_);
  nand (_35111_, _35110_, _35108_);
  nor (_35112_, _10544_, _10338_);
  nor (_35113_, _35112_, _10550_);
  and (_35114_, _35113_, _35111_);
  and (_35115_, _34993_, _10550_);
  nor (_35116_, _35115_, _35114_);
  or (_35117_, _35116_, _04920_);
  or (_35119_, _34982_, _04919_);
  and (_35120_, _35119_, _01995_);
  nand (_35121_, _35120_, _35117_);
  and (_35122_, _10174_, _01994_);
  nor (_35123_, _35122_, _07239_);
  nand (_35124_, _35123_, _35121_);
  and (_35125_, _10338_, _07239_);
  nor (_35126_, _35125_, _10149_);
  nand (_35127_, _35126_, _35124_);
  nor (_35128_, _10592_, \oc8051_golden_model_1.DPH [4]);
  nor (_35130_, _35128_, _10593_);
  nor (_35131_, _35130_, _10150_);
  nor (_35132_, _35131_, _10601_);
  and (_35133_, _35132_, _35127_);
  or (_35134_, _35133_, _34986_);
  nand (_35135_, _35134_, _10605_);
  nor (_35136_, _34993_, _07587_);
  nor (_35137_, _10338_, _10611_);
  nor (_35138_, _35137_, _10605_);
  not (_35139_, _35138_);
  nor (_35141_, _35139_, _35136_);
  nor (_35142_, _35141_, _10609_);
  nand (_35143_, _35142_, _35135_);
  nor (_35144_, _34979_, _10147_);
  nor (_35145_, _35144_, _10619_);
  nand (_35146_, _35145_, _35143_);
  nor (_35147_, _10618_, _34982_);
  nor (_35148_, _35147_, _02210_);
  nand (_35149_, _35148_, _35146_);
  and (_35150_, _10174_, _02210_);
  nor (_35151_, _35150_, _10626_);
  and (_35152_, _35151_, _35149_);
  or (_35153_, _35152_, _34985_);
  nand (_35154_, _35153_, _10630_);
  and (_35155_, _10338_, _10611_);
  and (_35156_, _34993_, _07587_);
  or (_35157_, _35156_, _35155_);
  and (_35158_, _35157_, _10629_);
  nor (_35159_, _35158_, _10634_);
  nand (_35160_, _35159_, _35154_);
  nor (_35162_, _34979_, _10139_);
  nor (_35163_, _35162_, _10136_);
  nand (_35164_, _35163_, _35160_);
  nor (_35165_, _34982_, _10135_);
  nor (_35166_, _35165_, _02206_);
  nand (_35167_, _35166_, _35164_);
  and (_35168_, _10174_, _02206_);
  nor (_35169_, _35168_, _09562_);
  and (_35170_, _35169_, _35167_);
  or (_35171_, _35170_, _34984_);
  nand (_35172_, _35171_, _10650_);
  or (_35173_, _34993_, \oc8051_golden_model_1.PSW [7]);
  or (_35174_, _10338_, _06707_);
  and (_35175_, _35174_, _10649_);
  and (_35176_, _35175_, _35173_);
  nor (_35177_, _35176_, _10654_);
  nand (_35178_, _35177_, _35172_);
  nor (_35179_, _34979_, _10133_);
  nor (_35180_, _35179_, _07340_);
  nand (_35181_, _35180_, _35178_);
  nor (_35183_, _34982_, _07339_);
  nor (_35184_, _35183_, _02202_);
  nand (_35185_, _35184_, _35181_);
  and (_35186_, _10174_, _02202_);
  nor (_35187_, _35186_, _10666_);
  and (_35188_, _35187_, _35185_);
  or (_35189_, _35188_, _34983_);
  nand (_35190_, _35189_, _10123_);
  nor (_35191_, _34993_, _06707_);
  nor (_35192_, _10338_, \oc8051_golden_model_1.PSW [7]);
  nor (_35193_, _35192_, _10123_);
  not (_35194_, _35193_);
  nor (_35195_, _35194_, _35191_);
  nor (_35196_, _35195_, _10671_);
  nand (_35197_, _35196_, _35190_);
  nor (_35198_, _34979_, _10120_);
  nor (_35199_, _35198_, _07386_);
  nand (_35200_, _35199_, _35197_);
  nor (_35201_, _34982_, _07385_);
  nor (_35202_, _35201_, _07415_);
  nand (_35204_, _35202_, _35200_);
  and (_35205_, _34980_, _07415_);
  nor (_35206_, _35205_, _02350_);
  and (_35207_, _35206_, _35204_);
  nor (_35208_, _04372_, _09472_);
  or (_35209_, _35208_, _01726_);
  or (_35210_, _35209_, _35207_);
  and (_35211_, _34982_, _01726_);
  nor (_35212_, _35211_, _02200_);
  nand (_35213_, _35212_, _35210_);
  nor (_35215_, _10173_, _08690_);
  and (_35216_, _35047_, _08690_);
  or (_35217_, _35216_, _10689_);
  nor (_35218_, _35217_, _35215_);
  nor (_35219_, _35218_, _10693_);
  nand (_35220_, _35219_, _35213_);
  nor (_35221_, _34979_, _10118_);
  nor (_35222_, _35221_, _07489_);
  nand (_35223_, _35222_, _35220_);
  nor (_35224_, _34982_, _07488_);
  nor (_35226_, _35224_, _07533_);
  and (_35227_, _35226_, _35223_);
  or (_35228_, _35227_, _34981_);
  nand (_35229_, _35228_, _02084_);
  and (_35230_, _04372_, _02083_);
  nor (_35231_, _35230_, _01738_);
  nand (_35232_, _35231_, _35229_);
  and (_35233_, _10338_, _01738_);
  nor (_35234_, _35233_, _02243_);
  nand (_35235_, _35234_, _35232_);
  nor (_35237_, _35021_, _08690_);
  and (_35238_, _10174_, _08690_);
  nor (_35239_, _35238_, _35237_);
  nor (_35240_, _35239_, _02367_);
  nor (_35241_, _35240_, _10723_);
  and (_35242_, _35241_, _35235_);
  nor (_35243_, _34980_, _10722_);
  or (_35244_, _35243_, _02366_);
  or (_35245_, _35244_, _35242_);
  nand (_35246_, _34982_, _02366_);
  and (_35247_, _35246_, _07581_);
  nand (_35248_, _35247_, _35245_);
  nor (_35249_, _34980_, _07581_);
  nor (_35250_, _35249_, _01989_);
  nand (_35251_, _35250_, _35248_);
  and (_35252_, _02825_, _01989_);
  nor (_35253_, _35252_, _01733_);
  nand (_35254_, _35253_, _35251_);
  and (_35255_, _10338_, _01733_);
  nor (_35256_, _35255_, _01697_);
  nand (_35258_, _35256_, _35254_);
  nor (_35259_, _35239_, _01698_);
  nor (_35260_, _35259_, _10744_);
  nand (_35261_, _35260_, _35258_);
  and (_35262_, _34979_, _10744_);
  nor (_35263_, _35262_, _02081_);
  nand (_35264_, _35263_, _35261_);
  and (_35265_, _34982_, _02081_);
  nor (_35266_, _35265_, _31497_);
  nand (_35267_, _35266_, _35264_);
  nor (_35270_, _34980_, _10751_);
  nor (_35271_, _35270_, _02198_);
  nand (_35272_, _35271_, _35267_);
  and (_35273_, _02825_, _02198_);
  nor (_35274_, _35273_, _01732_);
  nand (_35275_, _35274_, _35272_);
  and (_35276_, _10338_, _01732_);
  nor (_35277_, _35276_, _10762_);
  and (_35278_, _35277_, _35275_);
  and (_35279_, _34980_, _10762_);
  or (_35281_, _35279_, _35278_);
  nand (_35282_, _35281_, _39632_);
  or (_35283_, _39632_, \oc8051_golden_model_1.PC [12]);
  and (_35284_, _35283_, _39026_);
  and (_41806_, _35284_, _35282_);
  nor (_35285_, _10112_, \oc8051_golden_model_1.PC [13]);
  nor (_35286_, _35285_, _10113_);
  or (_35287_, _35286_, _10118_);
  or (_35288_, _35286_, _10120_);
  or (_35289_, _35286_, _10133_);
  or (_35291_, _35286_, _10139_);
  or (_35292_, _35286_, _10147_);
  and (_35293_, _10169_, _01765_);
  or (_35294_, _35286_, _10153_);
  not (_35295_, _35286_);
  nor (_35296_, _35295_, _10158_);
  and (_35297_, _10169_, _08842_);
  or (_35298_, _10171_, _10170_);
  not (_35299_, _35298_);
  nor (_35300_, _35299_, _10270_);
  and (_35302_, _35299_, _10270_);
  or (_35303_, _35302_, _35300_);
  and (_35304_, _35303_, _10482_);
  or (_35305_, _35304_, _35297_);
  and (_35306_, _35305_, _08790_);
  not (_35307_, _08770_);
  or (_35308_, _10169_, _35307_);
  or (_35309_, _35303_, _08770_);
  and (_35310_, _35309_, _10475_);
  and (_35311_, _35310_, _35308_);
  and (_35313_, _10334_, _02153_);
  or (_35314_, _10447_, _10334_);
  or (_35315_, _35303_, _10293_);
  or (_35316_, _10295_, _10169_);
  and (_35317_, _35316_, _02158_);
  and (_35318_, _35317_, _35315_);
  or (_35319_, _10336_, _10335_);
  not (_35320_, _35319_);
  nor (_35321_, _35320_, _10421_);
  and (_35322_, _35320_, _10421_);
  or (_35324_, _35322_, _35321_);
  and (_35325_, _35324_, _10437_);
  and (_35326_, _10435_, _10334_);
  or (_35327_, _35326_, _04534_);
  or (_35328_, _35327_, _35325_);
  and (_35329_, _11982_, _10317_);
  nor (_35330_, _02160_, \oc8051_golden_model_1.PC [13]);
  and (_35331_, _35330_, _09495_);
  and (_35332_, _35331_, _10312_);
  and (_35333_, _35332_, _06859_);
  or (_35335_, _35333_, _35329_);
  nand (_35336_, _35335_, _10299_);
  or (_35337_, _35286_, _34997_);
  and (_35338_, _35337_, _01752_);
  and (_35339_, _35338_, _35336_);
  or (_35340_, _11982_, _01752_);
  nand (_35341_, _35340_, _04534_);
  or (_35342_, _35341_, _35339_);
  and (_35343_, _35342_, _10442_);
  and (_35344_, _35343_, _35328_);
  or (_35346_, _35344_, _35318_);
  and (_35347_, _35346_, _10287_);
  nor (_35348_, _35295_, _10448_);
  or (_35349_, _35348_, _34737_);
  or (_35350_, _35349_, _35347_);
  and (_35351_, _35350_, _35314_);
  or (_35352_, _35351_, _22169_);
  or (_35353_, _35286_, _10452_);
  and (_35354_, _35353_, _02549_);
  and (_35355_, _35354_, _35352_);
  or (_35357_, _35355_, _35313_);
  and (_35358_, _35357_, _10460_);
  or (_35359_, _35295_, _10460_);
  nand (_35360_, _35359_, _10466_);
  or (_35361_, _35360_, _35358_);
  or (_35362_, _10466_, _10334_);
  and (_35363_, _35362_, _10471_);
  and (_35364_, _35363_, _35361_);
  or (_35365_, _35364_, _35311_);
  and (_35366_, _35365_, _08836_);
  or (_35368_, _35366_, _35306_);
  and (_35369_, _35368_, _08692_);
  and (_35370_, _10169_, _08877_);
  and (_35371_, _35303_, _10489_);
  or (_35372_, _35371_, _35370_);
  and (_35373_, _35372_, _02171_);
  or (_35374_, _35303_, _08922_);
  or (_35375_, _10169_, _32011_);
  and (_35376_, _35375_, _02246_);
  and (_35377_, _35376_, _35374_);
  or (_35379_, _35377_, _35373_);
  or (_35380_, _35379_, _35369_);
  and (_35381_, _35380_, _08882_);
  nand (_35382_, _35286_, _08881_);
  nand (_35383_, _35382_, _10506_);
  or (_35384_, _35383_, _35381_);
  or (_35385_, _10506_, _10334_);
  and (_35386_, _35385_, _10158_);
  and (_35387_, _35386_, _35384_);
  or (_35388_, _35387_, _35296_);
  and (_35390_, _35388_, _10515_);
  nor (_35391_, _10515_, _11982_);
  or (_35392_, _35391_, _10517_);
  or (_35393_, _35392_, _35390_);
  and (_35394_, _35393_, _35294_);
  or (_35395_, _35394_, _07017_);
  or (_35396_, _10334_, _07016_);
  and (_35397_, _35396_, _01778_);
  and (_35398_, _35397_, _35395_);
  or (_35399_, _35295_, _01778_);
  nand (_35401_, _35399_, _10527_);
  or (_35402_, _35401_, _35398_);
  or (_35403_, _10527_, _10334_);
  and (_35404_, _35403_, _07633_);
  and (_35405_, _35404_, _35402_);
  nand (_35406_, _10169_, _02218_);
  nand (_35407_, _35406_, _10534_);
  or (_35408_, _35407_, _35405_);
  or (_35409_, _10334_, _10534_);
  and (_35410_, _35409_, _02037_);
  and (_35412_, _35410_, _35408_);
  or (_35413_, _35412_, _35293_);
  and (_35414_, _35413_, _10542_);
  nor (_35415_, _35295_, _10542_);
  or (_35416_, _35415_, _10545_);
  or (_35417_, _35416_, _35414_);
  or (_35418_, _10544_, _10334_);
  and (_35419_, _35418_, _10551_);
  and (_35420_, _35419_, _35417_);
  and (_35421_, _35324_, _10550_);
  or (_35423_, _35421_, _04920_);
  or (_35424_, _35423_, _35420_);
  or (_35425_, _10334_, _04919_);
  and (_35426_, _35425_, _01995_);
  and (_35427_, _35426_, _35424_);
  and (_35428_, _10169_, _01994_);
  or (_35429_, _35428_, _07239_);
  or (_35430_, _35429_, _35427_);
  and (_35431_, _11982_, _07239_);
  nor (_35432_, _35431_, _10149_);
  and (_35434_, _35432_, _35430_);
  or (_35435_, _10593_, \oc8051_golden_model_1.DPH [5]);
  nor (_35436_, _10594_, _10150_);
  and (_35437_, _35436_, _35435_);
  or (_35438_, _35437_, _10601_);
  or (_35439_, _35438_, _35434_);
  or (_35440_, _10600_, _10334_);
  and (_35441_, _35440_, _10605_);
  and (_35442_, _35441_, _35439_);
  or (_35443_, _35324_, _07587_);
  or (_35445_, _10334_, _10611_);
  and (_35446_, _35445_, _10604_);
  and (_35447_, _35446_, _35443_);
  or (_35448_, _35447_, _10609_);
  or (_35449_, _35448_, _35442_);
  and (_35450_, _35449_, _35292_);
  or (_35451_, _35450_, _10619_);
  or (_35452_, _10618_, _10334_);
  and (_35453_, _35452_, _03059_);
  and (_35454_, _35453_, _35451_);
  nand (_35456_, _10169_, _02210_);
  nand (_35457_, _35456_, _10625_);
  or (_35458_, _35457_, _35454_);
  or (_35459_, _10625_, _10334_);
  and (_35460_, _35459_, _10630_);
  and (_35461_, _35460_, _35458_);
  or (_35462_, _35324_, _10611_);
  or (_35463_, _10334_, _07587_);
  and (_35464_, _35463_, _10629_);
  and (_35465_, _35464_, _35462_);
  or (_35467_, _35465_, _10634_);
  or (_35468_, _35467_, _35461_);
  and (_35469_, _35468_, _35291_);
  or (_35470_, _35469_, _10136_);
  or (_35471_, _10334_, _10135_);
  and (_35472_, _35471_, _02208_);
  and (_35473_, _35472_, _35470_);
  nand (_35474_, _10169_, _02206_);
  nand (_35475_, _35474_, _09561_);
  or (_35476_, _35475_, _35473_);
  nor (_35478_, _10649_, _11982_);
  or (_35479_, _35478_, _22844_);
  and (_35480_, _35479_, _35476_);
  or (_35481_, _35324_, \oc8051_golden_model_1.PSW [7]);
  or (_35482_, _10334_, _06707_);
  and (_35483_, _35482_, _10649_);
  and (_35484_, _35483_, _35481_);
  or (_35485_, _35484_, _10654_);
  or (_35486_, _35485_, _35480_);
  and (_35487_, _35486_, _35289_);
  or (_35490_, _35487_, _07340_);
  or (_35491_, _10334_, _07339_);
  and (_35492_, _35491_, _04953_);
  and (_35493_, _35492_, _35490_);
  nand (_35494_, _10169_, _02202_);
  nand (_35495_, _35494_, _10124_);
  or (_35496_, _35495_, _35493_);
  nor (_35497_, _11982_, _10122_);
  or (_35498_, _35497_, _22985_);
  and (_35499_, _35498_, _35496_);
  or (_35501_, _35324_, _06707_);
  or (_35502_, _10334_, \oc8051_golden_model_1.PSW [7]);
  and (_35503_, _35502_, _10122_);
  and (_35504_, _35503_, _35501_);
  or (_35505_, _35504_, _10671_);
  or (_35506_, _35505_, _35499_);
  and (_35507_, _35506_, _35288_);
  or (_35508_, _35507_, _07386_);
  or (_35509_, _10334_, _07385_);
  and (_35510_, _35509_, _07416_);
  and (_35512_, _35510_, _35508_);
  and (_35513_, _35286_, _07415_);
  or (_35514_, _35513_, _02350_);
  or (_35515_, _35514_, _35512_);
  nand (_35516_, _04057_, _02350_);
  and (_35517_, _35516_, _35515_);
  or (_35518_, _35517_, _01726_);
  nand (_35519_, _11982_, _01726_);
  and (_35520_, _35519_, _10689_);
  and (_35521_, _35520_, _35518_);
  or (_35523_, _35303_, _10694_);
  or (_35524_, _10169_, _08690_);
  and (_35525_, _35524_, _02200_);
  and (_35526_, _35525_, _35523_);
  or (_35527_, _35526_, _10693_);
  or (_35528_, _35527_, _35521_);
  and (_35529_, _35528_, _35287_);
  or (_35530_, _35529_, _07489_);
  or (_35531_, _10334_, _07488_);
  and (_35532_, _35531_, _07534_);
  and (_35534_, _35532_, _35530_);
  and (_35535_, _35286_, _07533_);
  or (_35536_, _35535_, _02083_);
  or (_35537_, _35536_, _35534_);
  nand (_35538_, _04057_, _02083_);
  and (_35539_, _35538_, _35537_);
  or (_35540_, _35539_, _01738_);
  nand (_35541_, _11982_, _01738_);
  and (_35542_, _35541_, _02367_);
  and (_35543_, _35542_, _35540_);
  or (_35545_, _10169_, _10694_);
  or (_35546_, _35303_, _08690_);
  and (_35547_, _35546_, _35545_);
  and (_35548_, _35547_, _02243_);
  or (_35549_, _35548_, _10723_);
  or (_35550_, _35549_, _35543_);
  or (_35551_, _35286_, _10722_);
  and (_35552_, _35551_, _02778_);
  and (_35553_, _35552_, _35550_);
  nand (_35554_, _10334_, _02366_);
  nand (_35556_, _35554_, _07581_);
  or (_35557_, _35556_, _35553_);
  or (_35558_, _35286_, _07581_);
  and (_35559_, _35558_, _05395_);
  and (_35560_, _35559_, _35557_);
  nor (_35561_, _02410_, _05395_);
  or (_35562_, _35561_, _01733_);
  or (_35563_, _35562_, _35560_);
  nand (_35564_, _11982_, _01733_);
  and (_35565_, _35564_, _01698_);
  and (_35567_, _35565_, _35563_);
  and (_35568_, _35547_, _01697_);
  or (_35569_, _35568_, _10744_);
  or (_35570_, _35569_, _35567_);
  nand (_35571_, _35295_, _10744_);
  and (_35572_, _35571_, _02082_);
  and (_35573_, _35572_, _35570_);
  nand (_35574_, _10334_, _02081_);
  nand (_35575_, _35574_, _10751_);
  or (_35576_, _35575_, _35573_);
  or (_35577_, _35286_, _10751_);
  and (_35578_, _35577_, _10755_);
  and (_35579_, _35578_, _35576_);
  nor (_35580_, _02410_, _10755_);
  or (_35581_, _35580_, _01732_);
  or (_35582_, _35581_, _35579_);
  nand (_35583_, _11982_, _01732_);
  and (_35584_, _35583_, _10763_);
  and (_35585_, _35584_, _35582_);
  and (_35586_, _35286_, _10762_);
  or (_35588_, _35586_, _35585_);
  or (_35589_, _35588_, _39633_);
  or (_35590_, _39632_, \oc8051_golden_model_1.PC [13]);
  and (_35591_, _35590_, _39026_);
  and (_41807_, _35591_, _35589_);
  nor (_35592_, _10113_, \oc8051_golden_model_1.PC [14]);
  nor (_35593_, _35592_, _10114_);
  not (_35594_, _35593_);
  and (_35595_, _35594_, _07533_);
  not (_35596_, _10328_);
  nor (_35598_, _35596_, _10124_);
  nor (_35599_, _35596_, _09561_);
  nor (_35600_, _10625_, _35596_);
  and (_35601_, _10163_, _02218_);
  nand (_35602_, _10162_, _08842_);
  and (_35603_, _10272_, _10167_);
  nor (_35604_, _35603_, _10273_);
  not (_35605_, _35604_);
  or (_35606_, _35605_, _08842_);
  and (_35607_, _35606_, _08790_);
  nand (_35609_, _35607_, _35602_);
  not (_35610_, _02230_);
  and (_35611_, _10163_, _08770_);
  nor (_35612_, _35604_, _08770_);
  nor (_35613_, _35612_, _35611_);
  and (_35614_, _35613_, _35610_);
  nor (_35615_, _35614_, _10471_);
  nor (_35616_, _35593_, _10452_);
  and (_35617_, _35593_, _02079_);
  and (_35618_, _10435_, _10328_);
  and (_35620_, _10423_, _10332_);
  nor (_35621_, _35620_, _10424_);
  and (_35622_, _35621_, _10437_);
  nor (_35623_, _35622_, _35618_);
  and (_35624_, _35623_, _04535_);
  and (_35625_, _35593_, _06845_);
  nor (_35626_, _35594_, _06859_);
  nor (_35627_, _35594_, _10312_);
  and (_35628_, _02063_, \oc8051_golden_model_1.PC [14]);
  and (_35629_, _35628_, _10299_);
  and (_35631_, _35629_, _10312_);
  and (_35632_, _35631_, _06859_);
  or (_35633_, _35632_, _35627_);
  and (_35634_, _35633_, _01747_);
  or (_35635_, _35634_, _35626_);
  and (_35636_, _35635_, _06847_);
  or (_35637_, _35636_, _35625_);
  and (_35638_, _35637_, _01752_);
  nor (_35639_, _34728_, _35596_);
  or (_35640_, _35639_, _04535_);
  nor (_35642_, _35640_, _35638_);
  or (_35643_, _35642_, _02079_);
  nor (_35644_, _35643_, _35624_);
  or (_35645_, _35644_, _35617_);
  and (_35646_, _35645_, _03006_);
  or (_35647_, _10295_, _10162_);
  or (_35648_, _35604_, _10293_);
  and (_35649_, _35648_, _35647_);
  and (_35650_, _35649_, _02158_);
  nor (_35651_, _35650_, _35646_);
  nand (_35653_, _35651_, _10287_);
  nor (_35654_, _35593_, _10287_);
  nor (_35655_, _35654_, _34737_);
  and (_35656_, _35655_, _35653_);
  nor (_35657_, _10447_, _35596_);
  nor (_35658_, _35657_, _35656_);
  and (_35659_, _35658_, _10452_);
  or (_35660_, _35659_, _35616_);
  nand (_35661_, _35660_, _02549_);
  and (_35662_, _35596_, _02153_);
  nor (_35664_, _35662_, _10462_);
  and (_35665_, _35664_, _35661_);
  nor (_35666_, _35594_, _10460_);
  or (_35667_, _35666_, _35665_);
  nand (_35668_, _35667_, _10466_);
  nor (_35669_, _10466_, _35596_);
  nor (_35670_, _35669_, _10470_);
  and (_35671_, _35670_, _35668_);
  nor (_35672_, _35671_, _35615_);
  and (_35673_, _35613_, _02230_);
  or (_35675_, _35673_, _08790_);
  or (_35676_, _35675_, _35672_);
  and (_35677_, _35676_, _35609_);
  and (_35678_, _35677_, _08692_);
  nor (_35679_, _35604_, _08877_);
  and (_35680_, _10163_, _08877_);
  or (_35681_, _35680_, _02547_);
  nor (_35682_, _35681_, _35679_);
  nor (_35683_, _35682_, _35678_);
  nand (_35684_, _10162_, _08922_);
  nand (_35686_, _35604_, _32011_);
  and (_35687_, _35686_, _35684_);
  or (_35688_, _35687_, _08917_);
  and (_35689_, _35688_, _35683_);
  or (_35690_, _35689_, _08881_);
  nand (_35691_, _35593_, _08881_);
  and (_35692_, _35691_, _35690_);
  and (_35693_, _35692_, _10506_);
  nor (_35694_, _10506_, _10328_);
  or (_35695_, _35694_, _35693_);
  nand (_35697_, _35695_, _10158_);
  nor (_35698_, _35593_, _10158_);
  nor (_35699_, _35698_, _34780_);
  nand (_35700_, _35699_, _35697_);
  nor (_35701_, _10515_, _35596_);
  nor (_35702_, _35701_, _10517_);
  nand (_35703_, _35702_, _35700_);
  nor (_35704_, _35593_, _10153_);
  nor (_35705_, _35704_, _07017_);
  nand (_35706_, _35705_, _35703_);
  nor (_35708_, _35596_, _07016_);
  nor (_35709_, _35708_, _01876_);
  nand (_35710_, _35709_, _35706_);
  nor (_35711_, _35593_, _01778_);
  nor (_35712_, _35711_, _10528_);
  nand (_35713_, _35712_, _35710_);
  nor (_35714_, _10527_, _35596_);
  nor (_35715_, _35714_, _02218_);
  nand (_35716_, _35715_, _35713_);
  nand (_35717_, _35716_, _10534_);
  or (_35719_, _35717_, _35601_);
  nor (_35720_, _35596_, _10534_);
  nor (_35721_, _35720_, _01765_);
  nand (_35722_, _35721_, _35719_);
  and (_35723_, _10163_, _01765_);
  nor (_35724_, _35723_, _10546_);
  nand (_35725_, _35724_, _35722_);
  nor (_35726_, _35594_, _10542_);
  nor (_35727_, _35726_, _10545_);
  nand (_35728_, _35727_, _35725_);
  nor (_35730_, _10544_, _10328_);
  nor (_35731_, _35730_, _10550_);
  and (_35732_, _35731_, _35728_);
  and (_35733_, _35621_, _10550_);
  nor (_35734_, _35733_, _35732_);
  or (_35735_, _35734_, _04920_);
  or (_35736_, _35596_, _04919_);
  and (_35737_, _35736_, _01995_);
  nand (_35738_, _35737_, _35735_);
  and (_35739_, _10163_, _01994_);
  nor (_35741_, _35739_, _07239_);
  nand (_35742_, _35741_, _35738_);
  and (_35743_, _10328_, _07239_);
  nor (_35744_, _35743_, _10149_);
  and (_35745_, _35744_, _35742_);
  nor (_35746_, _10594_, \oc8051_golden_model_1.DPH [6]);
  nor (_35747_, _35746_, _10595_);
  nor (_35748_, _35747_, _10150_);
  or (_35749_, _35748_, _35745_);
  nand (_35750_, _35749_, _10600_);
  nor (_35752_, _10600_, _10328_);
  nor (_35753_, _35752_, _10604_);
  nand (_35754_, _35753_, _35750_);
  and (_35755_, _10328_, _07587_);
  and (_35756_, _35621_, _10611_);
  or (_35757_, _35756_, _35755_);
  and (_35758_, _35757_, _10604_);
  nor (_35759_, _35758_, _10609_);
  nand (_35760_, _35759_, _35754_);
  nor (_35761_, _35593_, _10147_);
  nor (_35763_, _35761_, _10619_);
  nand (_35764_, _35763_, _35760_);
  nor (_35765_, _10618_, _35596_);
  nor (_35766_, _35765_, _02210_);
  nand (_35767_, _35766_, _35764_);
  and (_35768_, _10163_, _02210_);
  nor (_35769_, _35768_, _10626_);
  and (_35770_, _35769_, _35767_);
  or (_35771_, _35770_, _35600_);
  nand (_35772_, _35771_, _10630_);
  and (_35774_, _10328_, _10611_);
  and (_35775_, _35621_, _07587_);
  or (_35776_, _35775_, _35774_);
  and (_35777_, _35776_, _10629_);
  nor (_35778_, _35777_, _10634_);
  nand (_35779_, _35778_, _35772_);
  nor (_35780_, _35593_, _10139_);
  nor (_35781_, _35780_, _10136_);
  nand (_35782_, _35781_, _35779_);
  nor (_35783_, _35596_, _10135_);
  nor (_35785_, _35783_, _02206_);
  nand (_35786_, _35785_, _35782_);
  and (_35787_, _10163_, _02206_);
  nor (_35788_, _35787_, _09562_);
  and (_35789_, _35788_, _35786_);
  or (_35790_, _35789_, _35599_);
  nand (_35791_, _35790_, _10650_);
  or (_35792_, _35621_, \oc8051_golden_model_1.PSW [7]);
  or (_35793_, _10328_, _06707_);
  and (_35794_, _35793_, _10649_);
  and (_35796_, _35794_, _35792_);
  nor (_35797_, _35796_, _10654_);
  nand (_35798_, _35797_, _35791_);
  nor (_35799_, _35593_, _10133_);
  nor (_35800_, _35799_, _07340_);
  nand (_35801_, _35800_, _35798_);
  nor (_35802_, _35596_, _07339_);
  nor (_35803_, _35802_, _02202_);
  nand (_35804_, _35803_, _35801_);
  and (_35805_, _10163_, _02202_);
  nor (_35807_, _35805_, _10666_);
  and (_35808_, _35807_, _35804_);
  or (_35809_, _35808_, _35598_);
  nand (_35810_, _35809_, _10123_);
  nor (_35811_, _35621_, _06707_);
  nor (_35812_, _10328_, \oc8051_golden_model_1.PSW [7]);
  nor (_35813_, _35812_, _10123_);
  not (_35814_, _35813_);
  nor (_35815_, _35814_, _35811_);
  nor (_35816_, _35815_, _10671_);
  nand (_35818_, _35816_, _35810_);
  nor (_35819_, _35593_, _10120_);
  nor (_35820_, _35819_, _07386_);
  nand (_35821_, _35820_, _35818_);
  nor (_35822_, _35596_, _07385_);
  nor (_35823_, _35822_, _07415_);
  nand (_35824_, _35823_, _35821_);
  and (_35825_, _35594_, _07415_);
  nor (_35826_, _35825_, _02350_);
  and (_35827_, _35826_, _35824_);
  nor (_35829_, _03964_, _09472_);
  or (_35830_, _35829_, _01726_);
  or (_35831_, _35830_, _35827_);
  and (_35832_, _35596_, _01726_);
  nor (_35833_, _35832_, _02200_);
  nand (_35834_, _35833_, _35831_);
  and (_35835_, _35605_, _08690_);
  nor (_35836_, _10162_, _08690_);
  or (_35837_, _35836_, _10689_);
  nor (_35838_, _35837_, _35835_);
  nor (_35839_, _35838_, _10693_);
  nand (_35840_, _35839_, _35834_);
  nor (_35841_, _35593_, _10118_);
  nor (_35842_, _35841_, _07489_);
  nand (_35843_, _35842_, _35840_);
  nor (_35844_, _35596_, _07488_);
  nor (_35845_, _35844_, _07533_);
  and (_35846_, _35845_, _35843_);
  or (_35847_, _35846_, _35595_);
  nand (_35848_, _35847_, _02084_);
  and (_35850_, _03964_, _02083_);
  nor (_35851_, _35850_, _01738_);
  nand (_35852_, _35851_, _35848_);
  and (_35853_, _10328_, _01738_);
  nor (_35854_, _35853_, _02243_);
  nand (_35855_, _35854_, _35852_);
  and (_35856_, _10163_, _08690_);
  nor (_35857_, _35604_, _08690_);
  nor (_35858_, _35857_, _35856_);
  nor (_35859_, _35858_, _02367_);
  nor (_35861_, _35859_, _10723_);
  and (_35862_, _35861_, _35855_);
  nor (_35863_, _35594_, _10722_);
  or (_35864_, _35863_, _02366_);
  or (_35865_, _35864_, _35862_);
  nand (_35866_, _35596_, _02366_);
  and (_35867_, _35866_, _07581_);
  nand (_35868_, _35867_, _35865_);
  nor (_35869_, _35594_, _07581_);
  nor (_35870_, _35869_, _01989_);
  nand (_35872_, _35870_, _35868_);
  and (_35873_, _01989_, _02118_);
  nor (_35874_, _35873_, _01733_);
  nand (_35875_, _35874_, _35872_);
  and (_35876_, _10328_, _01733_);
  nor (_35877_, _35876_, _01697_);
  nand (_35878_, _35877_, _35875_);
  nor (_35879_, _35858_, _01698_);
  nor (_35880_, _35879_, _10744_);
  nand (_35881_, _35880_, _35878_);
  and (_35883_, _35593_, _10744_);
  nor (_35884_, _35883_, _02081_);
  nand (_35885_, _35884_, _35881_);
  and (_35886_, _35596_, _02081_);
  nor (_35887_, _35886_, _31497_);
  nand (_35888_, _35887_, _35885_);
  nor (_35889_, _35594_, _10751_);
  nor (_35890_, _35889_, _02198_);
  and (_35891_, _35890_, _35888_);
  and (_35892_, _02198_, _02118_);
  or (_35894_, _35892_, _35891_);
  nand (_35895_, _35894_, _10764_);
  and (_35896_, _35596_, _01732_);
  nor (_35897_, _35896_, _10762_);
  and (_35898_, _35897_, _35895_);
  and (_35899_, _35593_, _10762_);
  or (_35900_, _35899_, _35898_);
  or (_35901_, _35900_, _39633_);
  or (_35902_, _39632_, \oc8051_golden_model_1.PC [14]);
  and (_35903_, _35902_, _39026_);
  and (_41808_, _35903_, _35901_);
  and (_35905_, _39633_, \oc8051_golden_model_1.P0INREG [0]);
  or (_35906_, _35905_, _39993_);
  and (_41810_, _35906_, _39026_);
  and (_35907_, _39633_, \oc8051_golden_model_1.P0INREG [1]);
  or (_35908_, _35907_, _39978_);
  and (_41811_, _35908_, _39026_);
  and (_35909_, _39633_, \oc8051_golden_model_1.P0INREG [2]);
  or (_35910_, _35909_, _39971_);
  and (_41812_, _35910_, _39026_);
  and (_35912_, _39633_, \oc8051_golden_model_1.P0INREG [3]);
  or (_35913_, _35912_, _39986_);
  and (_41813_, _35913_, _39026_);
  and (_35914_, _39633_, \oc8051_golden_model_1.P0INREG [4]);
  or (_35915_, _35914_, _40050_);
  and (_41814_, _35915_, _39026_);
  and (_35916_, _39633_, \oc8051_golden_model_1.P0INREG [5]);
  or (_35917_, _35916_, _40020_);
  and (_41815_, _35917_, _39026_);
  and (_35918_, _39633_, \oc8051_golden_model_1.P0INREG [6]);
  or (_35920_, _35918_, _40006_);
  and (_41817_, _35920_, _39026_);
  and (_35921_, _39633_, \oc8051_golden_model_1.P1INREG [0]);
  or (_35922_, _35921_, _39644_);
  and (_41818_, _35922_, _39026_);
  and (_35923_, _39633_, \oc8051_golden_model_1.P1INREG [1]);
  or (_35924_, _35923_, _39635_);
  and (_41819_, _35924_, _39026_);
  and (_35925_, _39633_, \oc8051_golden_model_1.P1INREG [2]);
  or (_35926_, _35925_, _39653_);
  and (_41821_, _35926_, _39026_);
  and (_35928_, _39633_, \oc8051_golden_model_1.P1INREG [3]);
  or (_35929_, _35928_, _39661_);
  and (_41822_, _35929_, _39026_);
  and (_35930_, _39633_, \oc8051_golden_model_1.P1INREG [4]);
  or (_35931_, _35930_, _39679_);
  and (_41823_, _35931_, _39026_);
  and (_35932_, _39633_, \oc8051_golden_model_1.P1INREG [5]);
  or (_35933_, _35932_, _39672_);
  and (_41824_, _35933_, _39026_);
  and (_35935_, _39633_, \oc8051_golden_model_1.P1INREG [6]);
  or (_35936_, _35935_, _39687_);
  and (_41825_, _35936_, _39026_);
  and (_35937_, _39633_, \oc8051_golden_model_1.P2INREG [0]);
  or (_35938_, _35937_, _39795_);
  and (_41827_, _35938_, _39026_);
  and (_35939_, _39633_, \oc8051_golden_model_1.P2INREG [1]);
  or (_35940_, _35939_, _39844_);
  and (_41828_, _35940_, _39026_);
  and (_35941_, _39633_, \oc8051_golden_model_1.P2INREG [2]);
  or (_35943_, _35941_, _39828_);
  and (_41829_, _35943_, _39026_);
  and (_35944_, _39633_, \oc8051_golden_model_1.P2INREG [3]);
  or (_35945_, _35944_, _39811_);
  and (_41830_, _35945_, _39026_);
  and (_35946_, _39633_, \oc8051_golden_model_1.P2INREG [4]);
  or (_35947_, _35946_, _39802_);
  and (_41831_, _35947_, _39026_);
  and (_35948_, _39633_, \oc8051_golden_model_1.P2INREG [5]);
  or (_35949_, _35948_, _39851_);
  and (_41832_, _35949_, _39026_);
  and (_35951_, _39633_, \oc8051_golden_model_1.P2INREG [6]);
  or (_35952_, _35951_, _39835_);
  and (_41833_, _35952_, _39026_);
  and (_35953_, _39633_, \oc8051_golden_model_1.P3INREG [0]);
  or (_35954_, _35953_, _39727_);
  and (_41835_, _35954_, _39026_);
  and (_35955_, _39633_, \oc8051_golden_model_1.P3INREG [1]);
  or (_35956_, _35955_, _39776_);
  and (_41836_, _35956_, _39026_);
  and (_35958_, _39633_, \oc8051_golden_model_1.P3INREG [2]);
  or (_35959_, _35958_, _39760_);
  and (_41837_, _35959_, _39026_);
  and (_35960_, _39633_, \oc8051_golden_model_1.P3INREG [3]);
  or (_35961_, _35960_, _39743_);
  and (_41838_, _35961_, _39026_);
  and (_35962_, _39633_, \oc8051_golden_model_1.P3INREG [4]);
  or (_35963_, _35962_, _39734_);
  and (_41840_, _35963_, _39026_);
  and (_35964_, _39633_, \oc8051_golden_model_1.P3INREG [5]);
  or (_35966_, _35964_, _39783_);
  and (_41841_, _35966_, _39026_);
  and (_35967_, _39633_, \oc8051_golden_model_1.P3INREG [6]);
  or (_35968_, _35967_, _39767_);
  and (_41842_, _35968_, _39026_);
  and (_00006_[6], _39768_, _39026_);
  and (_00006_[5], _39784_, _39026_);
  and (_00006_[4], _39735_, _39026_);
  and (_00006_[3], _39744_, _39026_);
  and (_00006_[2], _39761_, _39026_);
  and (_00006_[1], _39777_, _39026_);
  and (_00006_[0], _39728_, _39026_);
  and (_00005_[6], _39836_, _39026_);
  and (_00005_[5], _39852_, _39026_);
  and (_00005_[4], _39803_, _39026_);
  and (_00005_[3], _39812_, _39026_);
  and (_00005_[2], _39829_, _39026_);
  and (_00005_[1], _39845_, _39026_);
  and (_00005_[0], _39796_, _39026_);
  and (_00004_[6], _39688_, _39026_);
  and (_00004_[5], _39673_, _39026_);
  and (_00004_[4], _39680_, _39026_);
  and (_00004_[3], _39662_, _39026_);
  and (_00004_[2], _39654_, _39026_);
  and (_00004_[1], _39636_, _39026_);
  and (_00004_[0], _39645_, _39026_);
  and (_00002_[6], _40008_, _39026_);
  and (_00002_[5], _40022_, _39026_);
  and (_00002_[4], _40052_, _39026_);
  and (_00002_[3], _39987_, _39026_);
  and (_00002_[2], _39972_, _39026_);
  and (_00002_[1], _39979_, _39026_);
  and (_00002_[0], _39994_, _39026_);
  and (_00004_[7], _39695_, _39026_);
  and (_00005_[7], _39819_, _39026_);
  and (_00006_[7], _39751_, _39026_);
  nor (_35972_, _08026_, _07919_);
  nor (_35973_, _09708_, _09461_);
  and (_35974_, _35973_, _35972_);
  nor (_35975_, _18119_, _17554_);
  nor (_35977_, _25628_, _18349_);
  and (_35978_, _35977_, _35975_);
  nor (_35979_, _28952_, _28435_);
  nor (_35980_, _28346_, _25409_);
  and (_35981_, _35980_, _35979_);
  nor (_35982_, _29563_, _29040_);
  nor (_35983_, _30165_, _29652_);
  and (_35984_, _35983_, _35982_);
  and (_35985_, _35984_, _35981_);
  or (_35986_, _30771_, _30252_);
  or (_35988_, _35986_, _30858_);
  nor (_35989_, _35988_, _17325_);
  and (_35990_, _35989_, _35985_);
  and (_35991_, _35990_, _35978_);
  not (_35992_, _25858_);
  nand (_35993_, _27255_, _35992_);
  or (_35994_, _35993_, _27485_);
  nor (_35995_, _35994_, _17785_);
  and (_35996_, _35995_, _35991_);
  or (_35997_, _25972_, _18464_);
  nor (_35999_, _35997_, _27599_);
  nor (_36000_, _09945_, _09866_);
  nor (_36001_, _10103_, _10024_);
  and (_36002_, _36001_, _36000_);
  or (_36003_, _30507_, _30420_);
  or (_36004_, _36003_, _30682_);
  nor (_36005_, _36004_, _09275_);
  nor (_36006_, _09787_, _09354_);
  and (_36007_, _36006_, _36005_);
  and (_36008_, _36007_, _36002_);
  nor (_36010_, _18234_, _17440_);
  and (_36011_, _36010_, _36008_);
  nor (_36012_, _25322_, _24808_);
  nor (_36013_, _24721_, _18008_);
  and (_36014_, _36013_, _36012_);
  nor (_36015_, _28086_, _27997_);
  nor (_36016_, _28603_, _28259_);
  and (_36017_, _36016_, _36015_);
  nor (_36018_, _24976_, _24634_);
  nor (_36019_, _25234_, _25062_);
  and (_36021_, _36019_, _36018_);
  and (_36022_, _36021_, _36017_);
  nor (_36023_, _29821_, _29473_);
  nor (_36024_, _30079_, _29907_);
  and (_36025_, _36024_, _36023_);
  nor (_36026_, _28864_, _28690_);
  nor (_36027_, _29298_, _29210_);
  and (_36028_, _36027_, _36026_);
  and (_36029_, _36028_, _36025_);
  and (_36030_, _36029_, _36022_);
  nor (_36032_, _29123_, _28517_);
  nor (_36033_, _30332_, _29735_);
  and (_36034_, _36033_, _36032_);
  nor (_36035_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_36036_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_36037_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_36038_, _36037_, _36036_);
  and (_36039_, _36038_, _36035_);
  nor (_36040_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_36041_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_36043_, _36041_, _36040_);
  nor (_36044_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_36045_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_36046_, _36045_, _36044_);
  and (_36047_, _36046_, _36043_);
  and (_36048_, _36047_, _36039_);
  nor (_36049_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_36050_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_36051_, _36050_, _36049_);
  nor (_36052_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_36054_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_36055_, _36054_, _36052_);
  and (_36056_, _36055_, _36051_);
  nor (_36057_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_36058_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_36059_, _36058_, _36057_);
  nor (_36060_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_36061_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_36062_, _36061_, _36060_);
  and (_36063_, _36062_, _36059_);
  and (_36065_, _36063_, _36056_);
  and (_36066_, _36065_, _36048_);
  nor (_36067_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_36068_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_36069_, _36068_, _36067_);
  nor (_36070_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_36071_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_36072_, _36071_, _36070_);
  and (_36073_, _36072_, _36069_);
  nor (_36074_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  nor (_36075_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  and (_36076_, _36075_, _36074_);
  nor (_36077_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_36078_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_36079_, _36078_, _36077_);
  and (_36080_, _36079_, _36076_);
  and (_36081_, _36080_, _36073_);
  nor (_36082_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_36083_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_36084_, _36083_, _36082_);
  nor (_36086_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  nor (_36087_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  and (_36088_, _36087_, _36086_);
  and (_36089_, _36088_, _36084_);
  nor (_36090_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_36091_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_36092_, _36091_, _36090_);
  nor (_36093_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_36094_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_36095_, _36094_, _36093_);
  and (_36097_, _36095_, _36092_);
  and (_36098_, _36097_, _36089_);
  and (_36099_, _36098_, _36081_);
  nor (_36100_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_36101_, _36100_, regs_always_zero);
  nor (_36102_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_36103_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_36104_, _36103_, _36102_);
  nor (_36105_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_36106_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_36108_, _36106_, _36105_);
  and (_36109_, _36108_, _36104_);
  and (_36110_, _36109_, _36101_);
  and (_36111_, \oc8051_golden_model_1.TCON [1], _27042_);
  nor (_36112_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_36113_, _36112_, _36111_);
  nor (_36114_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_36115_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_36116_, _36115_, _36114_);
  and (_36117_, _36116_, _36113_);
  nor (_36119_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_36120_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_36121_, _36120_, _36119_);
  nor (_36122_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_36123_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_36124_, _36123_, _36122_);
  and (_36125_, _36124_, _36121_);
  and (_36126_, _36125_, _36117_);
  and (_36127_, _36126_, _36110_);
  and (_36128_, _36127_, _36099_);
  nand (_36130_, _36128_, _36066_);
  nor (_36131_, _36130_, _24288_);
  nor (_36132_, _27911_, _24890_);
  and (_36133_, _36132_, _36131_);
  and (_36134_, _36133_, _36034_);
  nor (_36135_, _24462_, _24374_);
  and (_36136_, _36135_, _36134_);
  or (_36137_, _29994_, _29387_);
  nor (_36138_, _36137_, _30596_);
  nor (_36139_, _25149_, _24549_);
  nor (_36141_, _28778_, _28173_);
  and (_36142_, _36141_, _36139_);
  and (_36143_, _36142_, _36138_);
  nand (_36144_, _36143_, _36136_);
  nor (_36145_, _36144_, _17212_);
  and (_36146_, _36145_, _36030_);
  and (_36147_, _36146_, _36014_);
  and (_36148_, _36147_, _36011_);
  not (_36149_, _25516_);
  nor (_36150_, _25742_, _36149_);
  not (_36152_, _27144_);
  nor (_36153_, _27370_, _36152_);
  nand (_36154_, _36153_, _36150_);
  nor (_36155_, _36154_, _17670_);
  and (_36156_, _36155_, _36148_);
  and (_36157_, _36156_, _35999_);
  and (_36158_, _36157_, _35996_);
  or (_36159_, _27715_, _26202_);
  nor (_36160_, _36159_, _27830_);
  nor (_36161_, _18579_, _17900_);
  nor (_36163_, _26087_, _18694_);
  and (_36164_, _36163_, _36161_);
  and (_36165_, _36164_, _36160_);
  and (_36166_, _36165_, _36158_);
  and (_36167_, _36166_, _35974_);
  or (_00009_, _36167_, rst);
  or (_36168_, _09195_, _25218_);
  nand (_36169_, _23923_, _37436_);
  or (_36170_, _23923_, _37436_);
  or (_36171_, _23808_, _37312_);
  and (_36173_, _36171_, _39026_);
  and (_36174_, _36173_, _36170_);
  and (_36175_, _36174_, _36169_);
  not (_36176_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_36177_, _24038_, _36176_);
  nand (_36178_, _24038_, _36176_);
  not (_36179_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_36180_, _23468_, _36179_);
  or (_36181_, _23468_, _36179_);
  nand (_36182_, _23808_, _37312_);
  and (_36184_, _36182_, _36181_);
  and (_36185_, _36184_, _36180_);
  and (_36186_, _36185_, _36178_);
  and (_36187_, _36186_, _36177_);
  and (_36188_, _36187_, _36175_);
  nand (_36189_, _24206_, _25909_);
  or (_36190_, _24206_, _25909_);
  and (_36191_, _36190_, _36189_);
  and (_36192_, _36191_, _36188_);
  and (_36193_, _36192_, _36168_);
  nand (_36195_, _09195_, _25218_);
  nand (_36196_, _23695_, _25499_);
  or (_36197_, _23695_, _25499_);
  and (_36198_, _36197_, _36196_);
  and (_36199_, _36198_, _36195_);
  and (_00007_, _36199_, _36193_);
  or (_36200_, _09601_, _23389_);
  nand (_36201_, _26643_, _23713_);
  and (_36202_, _36201_, _36200_);
  nand (_36203_, _09601_, _23389_);
  or (_36205_, _26774_, _23789_);
  nand (_36206_, _26774_, _23789_);
  and (_36207_, _36206_, _36205_);
  and (_36208_, _36207_, _36203_);
  and (_36209_, _36208_, _36202_);
  or (_36210_, _27036_, _23939_);
  nand (_36211_, _27036_, _23939_);
  and (_36212_, _36211_, _36210_);
  nand (_36213_, _26524_, _23638_);
  and (_36214_, _36213_, _36212_);
  or (_36216_, _26905_, _23864_);
  or (_36217_, _26286_, _23486_);
  nand (_36218_, _26286_, _23486_);
  and (_36219_, _36218_, _36217_);
  and (_36220_, _36219_, _39026_);
  nand (_36221_, _26401_, _37499_);
  or (_36222_, _26401_, _37499_);
  and (_36223_, _36222_, _36221_);
  and (_36224_, _36223_, _36220_);
  and (_36225_, _36224_, _36216_);
  or (_36227_, _26524_, _23638_);
  nand (_36228_, _26905_, _23864_);
  or (_36229_, _26643_, _23713_);
  and (_36230_, _36229_, _36228_);
  and (_36231_, _36230_, _36227_);
  and (_36232_, _36231_, _36225_);
  and (_36233_, _36232_, _36214_);
  and (_00008_, _36233_, _36209_);
  nand (_36234_, _31510_, _41234_);
  or (_36235_, _31510_, _41234_);
  or (_36237_, _33323_, _41257_);
  nand (_36238_, _33323_, _41257_);
  nand (_36239_, _36238_, _36237_);
  nand (_36240_, _33691_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_36241_, _32245_, _41243_);
  or (_36242_, _33691_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_36243_, _36242_, _36241_);
  and (_36244_, _36243_, _36240_);
  or (_36245_, _32967_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_36246_, _34346_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_36248_, _34346_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_36249_, _10769_, _40434_);
  not (_36250_, _36249_);
  and (_36251_, _10769_, _40434_);
  nand (_36252_, _35900_, _41287_);
  or (_36253_, _35900_, _41287_);
  or (_36254_, _34670_, _40695_);
  nand (_36255_, _34670_, _40695_);
  nand (_36256_, _36255_, _36254_);
  or (_36257_, _35281_, _40693_);
  nand (_36259_, _35281_, _40693_);
  and (_36260_, _36259_, _36257_);
  nor (_36261_, _31121_, _41230_);
  and (_36262_, _31121_, _41230_);
  nor (_36263_, _36262_, _36261_);
  nor (_36264_, _36263_, _36260_);
  and (_36265_, _36264_, _36256_);
  and (_36266_, _36265_, _36253_);
  and (_36267_, _36266_, _36252_);
  and (_36268_, _35588_, _40691_);
  nor (_36270_, _35588_, _40691_);
  nor (_36271_, _36270_, _36268_);
  and (_36272_, _36271_, _36267_);
  or (_36273_, _34015_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_36274_, _34015_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_36275_, _36274_, _36273_);
  nand (_36276_, _36275_, _36272_);
  nor (_36277_, _36276_, _36251_);
  and (_36278_, _36277_, _36250_);
  and (_36279_, _34973_, _40694_);
  nor (_36281_, _34973_, _40694_);
  nor (_36282_, _36281_, _36279_);
  and (_36283_, _36282_, _36278_);
  nand (_36284_, _36283_, _36248_);
  nor (_36285_, _36284_, _36246_);
  and (_36286_, _36285_, _36245_);
  nand (_36287_, _32967_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_36288_, _32245_, _41243_);
  and (_36289_, _36288_, _36287_);
  and (_36290_, _36289_, _36286_);
  and (_36292_, _36290_, _36244_);
  or (_36293_, _32600_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_36294_, _32600_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_36295_, _36294_, _36293_);
  and (_36296_, _36295_, _36292_);
  and (_36297_, _36296_, _36239_);
  nand (_36298_, _31887_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_36299_, _31887_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_36300_, _36299_, _36298_);
  and (_36301_, _36300_, _36297_);
  and (_36303_, _36301_, _36235_);
  nand (_36304_, _36303_, _36234_);
  nand (_36305_, _36167_, _00001_);
  nor (_00003_, _36305_, _36304_);
  or (_36306_, _03948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_36307_, \oc8051_golden_model_1.P0 [0], _28142_);
  and (_36308_, _36307_, _36306_);
  or (_36309_, \oc8051_golden_model_1.IRAM[15] [0], _38194_);
  or (_36310_, _03950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_36311_, _36310_, _36309_);
  or (_36313_, \oc8051_golden_model_1.IRAM[14] [4], _38184_);
  or (_36314_, _03610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and (_36315_, _36314_, _36313_);
  and (_36316_, _36315_, _36311_);
  and (_36317_, \oc8051_golden_model_1.IRAM[13] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_36318_, \oc8051_golden_model_1.IRAM[13] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_36319_, _36318_, _36317_);
  and (_36320_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_36321_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_36322_, _36321_, _36320_);
  and (_36324_, _36322_, _36319_);
  or (_36325_, _04364_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_36326_, \oc8051_golden_model_1.IRAM[13] [6], _38167_);
  and (_36327_, _36326_, _36325_);
  or (_36328_, \oc8051_golden_model_1.IRAM[13] [4], _38162_);
  or (_36329_, _03616_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_36330_, _36329_, _36328_);
  and (_36331_, _36330_, _36327_);
  and (_36332_, _36331_, _36324_);
  and (_36333_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor (_36334_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_36335_, _36334_, _36333_);
  and (_36336_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_36337_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_36338_, _36337_, _36336_);
  or (_36339_, _02988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_36340_, \oc8051_golden_model_1.IRAM[14] [2], _38179_);
  and (_36341_, _36340_, _36339_);
  and (_36342_, _36341_, _36338_);
  and (_36343_, _36342_, _36335_);
  and (_36345_, _36343_, _36332_);
  and (_36346_, _36345_, _36316_);
  and (_36347_, _36346_, _36308_);
  and (_36348_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_36349_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_36350_, _36349_, _36348_);
  and (_36351_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_36352_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_36353_, _36352_, _36351_);
  and (_36354_, _36353_, _36350_);
  or (_36356_, _02994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_36357_, \oc8051_golden_model_1.IRAM[13] [2], _38157_);
  and (_36358_, _36357_, _36356_);
  or (_36359_, _03954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_36360_, \oc8051_golden_model_1.IRAM[13] [0], _38150_);
  and (_36361_, _36360_, _36359_);
  and (_36362_, _36361_, _36358_);
  and (_36363_, _36362_, _36354_);
  or (_36364_, _04342_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_36365_, \oc8051_golden_model_1.IRAM[11] [6], _38118_);
  and (_36366_, _36365_, _36364_);
  or (_36367_, _03594_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_36368_, \oc8051_golden_model_1.IRAM[11] [4], _38113_);
  and (_36369_, _36368_, _36367_);
  and (_36370_, _36369_, _36366_);
  and (_36371_, \oc8051_golden_model_1.IRAM[11] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_36372_, \oc8051_golden_model_1.IRAM[11] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_36373_, _36372_, _36371_);
  and (_36374_, \oc8051_golden_model_1.IRAM[12] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_36375_, \oc8051_golden_model_1.IRAM[12] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_36377_, _36375_, _36374_);
  and (_36378_, _36377_, _36373_);
  and (_36379_, _36378_, _36370_);
  nor (_36380_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_36381_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_36382_, _36381_, _36380_);
  nor (_36383_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_36384_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_36385_, _36384_, _36383_);
  and (_36386_, _36385_, _36382_);
  or (_36388_, _04362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_36389_, \oc8051_golden_model_1.IRAM[12] [6], _38144_);
  and (_36390_, _36389_, _36388_);
  or (_36391_, _03614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_36392_, \oc8051_golden_model_1.IRAM[12] [4], _38138_);
  and (_36393_, _36392_, _36391_);
  and (_36394_, _36393_, _36390_);
  and (_36395_, _36394_, _36386_);
  nor (_36396_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_36397_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_36398_, _36397_, _36396_);
  and (_36399_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_36400_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_36401_, _36400_, _36399_);
  and (_36402_, _36401_, _36398_);
  or (_36403_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_36404_, \oc8051_golden_model_1.IRAM[12] [2], _38132_);
  and (_36405_, _36404_, _36403_);
  or (_36406_, \oc8051_golden_model_1.IRAM[12] [0], _38124_);
  or (_36407_, _03934_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_36409_, _36407_, _36406_);
  and (_36410_, _36409_, _36405_);
  and (_36411_, _36410_, _36402_);
  and (_36412_, _36411_, _36395_);
  and (_36413_, _36412_, _36379_);
  and (_36414_, _36413_, _36363_);
  and (_36415_, _36414_, _36347_);
  or (_36416_, _20786_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_36417_, \oc8051_golden_model_1.P2 [6], _31143_);
  and (_36418_, _36417_, _36416_);
  or (_36420_, \oc8051_golden_model_1.P2 [4], _30817_);
  or (_36421_, _20563_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_36422_, _36421_, _36420_);
  and (_36423_, _36422_, _36418_);
  and (_36424_, \oc8051_golden_model_1.P2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_36425_, \oc8051_golden_model_1.P2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_36426_, _36425_, _36424_);
  and (_36427_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_36428_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_36429_, _36428_, _36427_);
  and (_36431_, _36429_, _36426_);
  and (_36432_, _36431_, _36423_);
  and (_36433_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_36434_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_36435_, _36434_, _36433_);
  and (_36436_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_36437_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_36438_, _36437_, _36436_);
  and (_36439_, _36438_, _36435_);
  or (_36440_, \oc8051_golden_model_1.P3 [2], _31634_);
  or (_36442_, _21119_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_36443_, _36442_, _36440_);
  or (_36444_, _21008_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_36445_, \oc8051_golden_model_1.P3 [0], _31307_);
  and (_36446_, _36445_, _36444_);
  and (_36447_, _36446_, _36443_);
  and (_36448_, _36447_, _36439_);
  and (_36449_, _36448_, _36432_);
  and (_36450_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_36451_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_36453_, _36451_, _36450_);
  and (_36454_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_36455_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_36456_, _36455_, _36454_);
  and (_36457_, _36456_, _36453_);
  or (_36458_, \oc8051_golden_model_1.P1 [6], _30061_);
  or (_36459_, _20014_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_36460_, _36459_, _36458_);
  or (_36461_, _19793_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_36462_, \oc8051_golden_model_1.P1 [4], _29758_);
  and (_36464_, _36462_, _36461_);
  and (_36465_, _36464_, _36460_);
  and (_36466_, _36465_, _36457_);
  and (_36467_, \oc8051_golden_model_1.P1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_36468_, \oc8051_golden_model_1.P1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_36469_, _36468_, _36467_);
  and (_36470_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_36471_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_36472_, _36471_, _36470_);
  or (_36473_, _20348_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_36475_, \oc8051_golden_model_1.P2 [2], _30493_);
  and (_36476_, _36475_, _36473_);
  and (_36477_, _36476_, _36472_);
  and (_36478_, _36477_, _36469_);
  and (_36479_, _36478_, _36466_);
  and (_36480_, _36479_, _36449_);
  and (_36481_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_36482_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_36483_, _36482_, _36481_);
  and (_36484_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_36486_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_36487_, _36486_, _36484_);
  and (_36488_, _36487_, _36483_);
  or (_36489_, \oc8051_golden_model_1.P3 [7], _27969_);
  or (_36490_, _21780_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_36491_, _08356_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_36492_, _36491_, _36490_);
  and (_36493_, _36492_, _36489_);
  or (_36494_, _21558_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_36495_, \oc8051_golden_model_1.P3 [6], _32288_);
  and (_36496_, _36495_, _36494_);
  or (_36497_, _21335_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_36498_, \oc8051_golden_model_1.P3 [4], _31961_);
  and (_36499_, _36498_, _36497_);
  and (_36500_, _36499_, _36496_);
  and (_36501_, _36500_, _36493_);
  and (_36502_, _36501_, _36488_);
  or (_36503_, \oc8051_golden_model_1.P2 [0], _30169_);
  or (_36504_, _20236_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_36505_, _36504_, _36503_);
  and (_36507_, _36505_, _36502_);
  and (_36508_, _36507_, _36480_);
  or (_36509_, _03936_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_36510_, \oc8051_golden_model_1.IRAM[11] [0], _38099_);
  and (_36511_, _36510_, _36509_);
  or (_36512_, \oc8051_golden_model_1.IRAM[9] [6], _38067_);
  or (_36513_, _04350_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_36514_, _36513_, _36512_);
  or (_36515_, _03602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_36516_, \oc8051_golden_model_1.IRAM[9] [4], _38062_);
  and (_36518_, _36516_, _36515_);
  and (_36519_, _36518_, _36514_);
  and (_36520_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_36521_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_36522_, _36521_, _36520_);
  and (_36523_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_36524_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_36525_, _36524_, _36523_);
  and (_36526_, _36525_, _36522_);
  and (_36527_, _36526_, _36519_);
  nor (_36529_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_36530_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_36531_, _36530_, _36529_);
  nor (_36532_, \oc8051_golden_model_1.IRAM[9] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_36533_, \oc8051_golden_model_1.IRAM[9] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_36534_, _36533_, _36532_);
  and (_36535_, _36534_, _36531_);
  or (_36536_, \oc8051_golden_model_1.IRAM[10] [2], _38080_);
  or (_36537_, _02974_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_36538_, _36537_, _36536_);
  or (_36540_, \oc8051_golden_model_1.IRAM[10] [0], _38072_);
  or (_36541_, _03942_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_36542_, _36541_, _36540_);
  and (_36543_, _36542_, _36538_);
  and (_36544_, _36543_, _36535_);
  and (_36545_, _36544_, _36527_);
  nor (_36546_, \oc8051_golden_model_1.IRAM[10] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and (_36547_, \oc8051_golden_model_1.IRAM[10] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_36548_, _36547_, _36546_);
  and (_36549_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_36551_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_36552_, _36551_, _36549_);
  and (_36553_, _36552_, _36548_);
  or (_36554_, \oc8051_golden_model_1.IRAM[10] [6], _38093_);
  or (_36555_, _04344_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_36556_, _36555_, _36554_);
  or (_36557_, \oc8051_golden_model_1.IRAM[10] [4], _38087_);
  or (_36558_, _03596_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_36559_, _36558_, _36557_);
  and (_36560_, _36559_, _36556_);
  and (_36562_, _36560_, _36553_);
  and (_36563_, \oc8051_golden_model_1.IRAM[10] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor (_36564_, \oc8051_golden_model_1.IRAM[10] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_36565_, _36564_, _36563_);
  and (_36566_, \oc8051_golden_model_1.IRAM[11] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_36567_, \oc8051_golden_model_1.IRAM[11] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_36568_, _36567_, _36566_);
  or (_36569_, \oc8051_golden_model_1.IRAM[11] [2], _38107_);
  or (_36570_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_36571_, _36570_, _36569_);
  and (_36573_, _36571_, _36568_);
  and (_36574_, _36573_, _36565_);
  and (_36575_, _36574_, _36562_);
  and (_36576_, _36575_, _36545_);
  and (_36577_, _36576_, _36511_);
  or (_36578_, _03956_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_36579_, \oc8051_golden_model_1.IRAM[14] [0], _38172_);
  and (_36580_, _36579_, _36578_);
  and (_36581_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_36582_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_36584_, _36582_, _36581_);
  and (_36585_, \oc8051_golden_model_1.IRAM[14] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_36586_, \oc8051_golden_model_1.IRAM[14] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_36587_, _36586_, _36585_);
  or (_36588_, _04358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_36589_, \oc8051_golden_model_1.IRAM[14] [6], _38189_);
  and (_36590_, _36589_, _36588_);
  and (_36591_, _36590_, _36587_);
  and (_36592_, _36591_, _36584_);
  and (_36593_, \oc8051_golden_model_1.IRAM[14] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor (_36594_, \oc8051_golden_model_1.IRAM[14] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_36595_, _36594_, _36593_);
  and (_36596_, \oc8051_golden_model_1.IRAM[15] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_36597_, \oc8051_golden_model_1.IRAM[15] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_36598_, _36597_, _36596_);
  or (_36599_, _02986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_36600_, \oc8051_golden_model_1.IRAM[15] [2], _38199_);
  and (_36601_, _36600_, _36599_);
  and (_36602_, _36601_, _36598_);
  and (_36603_, _36602_, _36595_);
  and (_36605_, _36603_, _36592_);
  and (_36606_, _36605_, _36580_);
  or (_36607_, \oc8051_golden_model_1.P0 [6], _29039_);
  or (_36608_, _19189_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_36609_, _36608_, _36607_);
  or (_36610_, \oc8051_golden_model_1.P0 [4], _28736_);
  or (_36611_, _18941_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_36612_, _36611_, _36610_);
  and (_36613_, _36612_, _36609_);
  and (_36614_, \oc8051_golden_model_1.P0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_36616_, \oc8051_golden_model_1.P0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_36617_, _36616_, _36614_);
  and (_36618_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_36619_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_36620_, _36619_, _36618_);
  and (_36621_, _36620_, _36617_);
  and (_36622_, _36621_, _36613_);
  and (_36623_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_36624_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_36625_, _36624_, _36623_);
  and (_36627_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_36628_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_36629_, _36628_, _36627_);
  and (_36630_, _36629_, _36625_);
  or (_36631_, _19577_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_36632_, \oc8051_golden_model_1.P1 [2], _29464_);
  and (_36633_, _36632_, _36631_);
  or (_36634_, _19451_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_36635_, \oc8051_golden_model_1.P1 [0], _29181_);
  and (_36636_, _36635_, _36634_);
  and (_36638_, _36636_, _36633_);
  and (_36639_, _36638_, _36630_);
  and (_36640_, _36639_, _36622_);
  and (_36641_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_36642_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_36643_, _36642_, _36641_);
  and (_36644_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_36645_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_36646_, _36645_, _36644_);
  and (_36647_, _36646_, _36643_);
  or (_36649_, _04356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_36650_, \oc8051_golden_model_1.IRAM[15] [6], _38210_);
  and (_36651_, _36650_, _36649_);
  or (_36652_, \oc8051_golden_model_1.IRAM[15] [4], _38204_);
  or (_36653_, _03608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_36654_, _36653_, _36652_);
  and (_36655_, _36654_, _36651_);
  and (_36656_, _36655_, _36647_);
  and (_36657_, \oc8051_golden_model_1.IRAM[15] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_36658_, \oc8051_golden_model_1.IRAM[15] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_36660_, _36658_, _36657_);
  and (_36661_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_36662_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_36663_, _36662_, _36661_);
  or (_36664_, _18699_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_36665_, \oc8051_golden_model_1.P0 [2], _28401_);
  and (_36666_, _36665_, _36664_);
  and (_36667_, _36666_, _36663_);
  and (_36668_, _36667_, _36660_);
  and (_36669_, _36668_, _36656_);
  and (_36671_, _36669_, _36640_);
  and (_36672_, _36671_, _36606_);
  and (_36673_, _36672_, _36577_);
  and (_36674_, _36673_, _36508_);
  or (_36675_, _06224_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_36676_, \oc8051_golden_model_1.B [6], _18490_);
  and (_36677_, _36676_, _36675_);
  or (_36678_, _06222_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_36679_, \oc8051_golden_model_1.B [4], _18143_);
  and (_36680_, _36679_, _36678_);
  and (_36682_, _36680_, _36677_);
  and (_36683_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_36684_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_36685_, _36684_, _36683_);
  and (_36686_, \oc8051_golden_model_1.B [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_36687_, \oc8051_golden_model_1.B [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_36688_, _36687_, _36686_);
  and (_36689_, _36688_, _36685_);
  and (_36690_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_36691_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_36692_, _36691_, _36690_);
  and (_36693_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_36694_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_36695_, _36694_, _36693_);
  and (_36696_, _36695_, _36692_);
  nand (_36697_, _15995_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_36698_, _15813_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_36699_, _36698_, _36697_);
  or (_36700_, _06475_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_36701_, _15813_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_36703_, _36701_, _36700_);
  and (_36704_, _36703_, _36699_);
  and (_36705_, _36704_, _36696_);
  and (_36706_, _36705_, _36689_);
  and (_36707_, _36706_, _36682_);
  and (_36708_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_36709_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_36710_, _36709_, _36708_);
  and (_36711_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_36712_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_36714_, _36712_, _36711_);
  and (_36715_, _36714_, _36710_);
  or (_36716_, _06283_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_36717_, \oc8051_golden_model_1.ACC [6], _27275_);
  and (_36718_, _36717_, _36716_);
  or (_36719_, \oc8051_golden_model_1.ACC [4], _26994_);
  or (_36720_, _06383_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_36721_, _36720_, _36719_);
  and (_36722_, _36721_, _36718_);
  nor (_36723_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_36725_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_36726_, _36725_, _36723_);
  or (_36727_, _01887_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_36728_, \oc8051_golden_model_1.ACC [2], _26690_);
  and (_36729_, _36728_, _36727_);
  and (_36730_, _36729_, _36726_);
  or (_36731_, \oc8051_golden_model_1.ACC [0], _26452_);
  and (_36732_, inst_finished_r, p1_valid_r);
  and (_36733_, _36732_, _36731_);
  and (_36734_, _36733_, _36730_);
  nor (_36736_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_36737_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_36738_, _36737_, _36736_);
  nor (_36739_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_36740_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_36741_, _36740_, _36739_);
  and (_36742_, _36741_, _36738_);
  or (_36743_, _06214_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_36744_, \oc8051_golden_model_1.B [2], _17796_);
  and (_36745_, _36744_, _36743_);
  or (_36747_, \oc8051_golden_model_1.B [0], _17373_);
  or (_36748_, _06231_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_36749_, _36748_, _36747_);
  and (_36750_, _36749_, _36745_);
  and (_36751_, _36750_, _36742_);
  and (_36752_, _36751_, _36734_);
  and (_36753_, _36752_, _36722_);
  and (_36754_, _36753_, _36715_);
  and (_36755_, _36754_, _36707_);
  or (_36756_, \oc8051_golden_model_1.IRAM[2] [6], _37906_);
  or (_36758_, _04320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_36759_, _36758_, _36756_);
  or (_36760_, \oc8051_golden_model_1.IRAM[2] [4], _37901_);
  or (_36761_, _03572_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_36762_, _36761_, _36760_);
  and (_36763_, _36762_, _36759_);
  and (_36764_, \oc8051_golden_model_1.IRAM[2] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_36765_, \oc8051_golden_model_1.IRAM[2] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_36766_, _36765_, _36764_);
  nor (_36767_, \oc8051_golden_model_1.IRAM[3] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_36769_, \oc8051_golden_model_1.IRAM[3] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_36770_, _36769_, _36767_);
  and (_36771_, _36770_, _36766_);
  and (_36772_, _36771_, _36763_);
  and (_36773_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_36774_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_36775_, _36774_, _36773_);
  and (_36776_, \oc8051_golden_model_1.IRAM[1] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_36777_, \oc8051_golden_model_1.IRAM[1] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_36778_, _36777_, _36776_);
  and (_36779_, _36778_, _36775_);
  or (_36780_, _03906_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_36781_, \oc8051_golden_model_1.IRAM[2] [0], _37888_);
  and (_36782_, _36781_, _36780_);
  or (_36783_, \oc8051_golden_model_1.IRAM[2] [2], _37896_);
  or (_36784_, _02948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_36785_, _36784_, _36783_);
  and (_36786_, _36785_, _36782_);
  and (_36787_, _36786_, _36779_);
  and (_36788_, _36787_, _36772_);
  and (_36790_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_36791_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_36792_, _36791_, _36790_);
  or (_36793_, \oc8051_golden_model_1.IRAM[4] [6], _37952_);
  or (_36794_, _04332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_36795_, _36794_, _36793_);
  and (_36796_, _36795_, _36792_);
  and (_36797_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_36798_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_36799_, _36798_, _36797_);
  or (_36801_, \oc8051_golden_model_1.IRAM[4] [4], _37947_);
  or (_36802_, _03584_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_36803_, _36802_, _36801_);
  and (_36804_, _36803_, _36799_);
  and (_36805_, _36804_, _36796_);
  and (_36806_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_36807_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_36808_, _36807_, _36806_);
  or (_36809_, _04318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_36810_, \oc8051_golden_model_1.IRAM[3] [6], _37929_);
  and (_36812_, _36810_, _36809_);
  and (_36813_, _36812_, _36808_);
  and (_36814_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_36815_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_36816_, _36815_, _36814_);
  or (_36817_, \oc8051_golden_model_1.IRAM[3] [4], _37924_);
  or (_36818_, _03570_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  and (_36819_, _36818_, _36817_);
  and (_36820_, _36819_, _36816_);
  and (_36821_, _36820_, _36813_);
  and (_36823_, _36821_, _36805_);
  and (_36824_, \oc8051_golden_model_1.IRAM[2] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_36825_, \oc8051_golden_model_1.IRAM[2] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_36826_, _36825_, _36824_);
  nor (_36827_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_36828_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_36829_, _36828_, _36827_);
  and (_36830_, _36829_, _36826_);
  or (_36831_, _02945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_36832_, \oc8051_golden_model_1.IRAM[3] [2], _37918_);
  and (_36834_, _36832_, _36831_);
  or (_36835_, _03912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_36836_, \oc8051_golden_model_1.IRAM[3] [0], _37911_);
  and (_36837_, _36836_, _36835_);
  and (_36838_, _36837_, _36834_);
  and (_36839_, _36838_, _36830_);
  or (_36840_, \oc8051_golden_model_1.IRAM[1] [6], _37883_);
  or (_36841_, _04314_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_36842_, _36841_, _36840_);
  or (_36843_, _03566_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_36845_, \oc8051_golden_model_1.IRAM[1] [4], _37877_);
  and (_36846_, _36845_, _36843_);
  and (_36847_, _36846_, _36842_);
  nor (_36848_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_36849_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_36850_, _36849_, _36848_);
  nor (_36851_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_36852_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_36853_, _36852_, _36851_);
  and (_36854_, _36853_, _36850_);
  and (_36856_, _36854_, _36847_);
  and (_36857_, _36856_, _36839_);
  nor (_36858_, \oc8051_golden_model_1.IRAM[4] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_36859_, \oc8051_golden_model_1.IRAM[4] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_36860_, _36859_, _36858_);
  and (_36861_, \oc8051_golden_model_1.IRAM[3] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_36862_, \oc8051_golden_model_1.IRAM[3] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_36863_, _36862_, _36861_);
  and (_36864_, _36863_, _36860_);
  or (_36865_, _02961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_36866_, \oc8051_golden_model_1.IRAM[4] [2], _37942_);
  and (_36867_, _36866_, _36865_);
  or (_36868_, \oc8051_golden_model_1.IRAM[4] [0], _37934_);
  or (_36869_, _03910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_36870_, _36869_, _36868_);
  and (_36871_, _36870_, _36867_);
  and (_36872_, _36871_, _36864_);
  and (_36873_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_36874_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_36875_, _36874_, _36873_);
  and (_36877_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor (_36878_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_36879_, _36878_, _36877_);
  and (_36880_, _36879_, _36875_);
  or (_36881_, \oc8051_golden_model_1.IRAM[5] [2], _37964_);
  or (_36882_, _02963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_36883_, _36882_, _36881_);
  or (_36884_, \oc8051_golden_model_1.IRAM[5] [0], _37957_);
  or (_36885_, _03924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_36886_, _36885_, _36884_);
  and (_36888_, _36886_, _36883_);
  and (_36889_, _36888_, _36880_);
  and (_36890_, _36889_, _36872_);
  and (_36891_, _36890_, _36857_);
  and (_36892_, _36891_, _36823_);
  and (_36893_, _36892_, _36788_);
  and (_36894_, _36893_, _36755_);
  and (_36895_, _36894_, _36674_);
  and (_36896_, _36895_, _36415_);
  or (_36897_, _23389_, \oc8051_golden_model_1.SP [7]);
  nand (_36899_, _23389_, \oc8051_golden_model_1.SP [7]);
  and (_36900_, _36899_, _36897_);
  or (_36901_, _23939_, \oc8051_golden_model_1.SP [6]);
  nand (_36902_, _23939_, \oc8051_golden_model_1.SP [6]);
  and (_36903_, _36902_, _36901_);
  nand (_36904_, _23864_, \oc8051_golden_model_1.SP [5]);
  or (_36905_, _23864_, \oc8051_golden_model_1.SP [5]);
  and (_36906_, _36905_, _36904_);
  nand (_36907_, _23713_, \oc8051_golden_model_1.SP [3]);
  or (_36908_, _23713_, \oc8051_golden_model_1.SP [3]);
  and (_36910_, _36908_, _36907_);
  or (_36911_, _23562_, \oc8051_golden_model_1.SP [1]);
  or (_36912_, _23486_, \oc8051_golden_model_1.SP [0]);
  nand (_36913_, _23486_, \oc8051_golden_model_1.SP [0]);
  and (_36914_, _36913_, _36912_);
  nand (_36915_, _23562_, \oc8051_golden_model_1.SP [1]);
  and (_36916_, _36915_, _36914_);
  and (_36917_, _36916_, _36911_);
  or (_36918_, _23638_, \oc8051_golden_model_1.SP [2]);
  nand (_36919_, _23638_, \oc8051_golden_model_1.SP [2]);
  and (_36921_, _36919_, _36918_);
  and (_36922_, _36921_, _36917_);
  and (_36923_, _36922_, _36910_);
  or (_36924_, _23789_, \oc8051_golden_model_1.SP [4]);
  nand (_36925_, _23789_, \oc8051_golden_model_1.SP [4]);
  and (_36926_, _36925_, _36924_);
  and (_36927_, _36926_, _36923_);
  and (_36928_, _36927_, _36906_);
  and (_36929_, _36928_, _36903_);
  and (_36930_, _36929_, _36900_);
  or (_36932_, _36930_, property_valid_sp_1_r);
  or (_36933_, \oc8051_golden_model_1.IRAM[7] [0], _38002_);
  or (_36934_, _03920_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_36935_, _36934_, _36933_);
  and (_36936_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_36937_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_36938_, _36937_, _36936_);
  and (_36939_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_36940_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_36941_, _36940_, _36939_);
  and (_36943_, _36941_, _36938_);
  or (_36944_, _02980_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_36945_, \oc8051_golden_model_1.IRAM[9] [2], _38057_);
  and (_36946_, _36945_, _36944_);
  or (_36947_, _03940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_36948_, \oc8051_golden_model_1.IRAM[9] [0], _38050_);
  and (_36949_, _36948_, _36947_);
  and (_36950_, _36949_, _36946_);
  and (_36951_, _36950_, _36943_);
  and (_36952_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_36953_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_36954_, _36953_, _36952_);
  or (_36955_, \oc8051_golden_model_1.IRAM[7] [6], _38020_);
  or (_36956_, _04326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_36957_, _36956_, _36955_);
  and (_36958_, _36957_, _36954_);
  and (_36959_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_36960_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_36961_, _36960_, _36959_);
  or (_36962_, _03578_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_36964_, \oc8051_golden_model_1.IRAM[7] [4], _38014_);
  and (_36965_, _36964_, _36962_);
  and (_36966_, _36965_, _36961_);
  and (_36967_, _36966_, _36958_);
  and (_36968_, _36967_, _36951_);
  and (_36969_, \oc8051_golden_model_1.IRAM[8] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_36970_, \oc8051_golden_model_1.IRAM[8] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_36971_, _36970_, _36969_);
  and (_36972_, \oc8051_golden_model_1.IRAM[7] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_36973_, \oc8051_golden_model_1.IRAM[7] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_36975_, _36973_, _36972_);
  and (_36976_, _36975_, _36971_);
  or (_36977_, \oc8051_golden_model_1.IRAM[8] [2], _38033_);
  or (_36978_, _02978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_36979_, _36978_, _36977_);
  or (_36980_, _03918_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_36981_, \oc8051_golden_model_1.IRAM[8] [0], _38025_);
  and (_36982_, _36981_, _36980_);
  and (_36983_, _36982_, _36979_);
  and (_36984_, _36983_, _36976_);
  or (_36986_, \oc8051_golden_model_1.IRAM[8] [6], _38045_);
  or (_36987_, _04348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_36988_, _36987_, _36986_);
  or (_36989_, \oc8051_golden_model_1.IRAM[8] [4], _38039_);
  or (_36990_, _03600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_36991_, _36990_, _36989_);
  and (_36992_, _36991_, _36988_);
  and (_36993_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_36994_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_36995_, _36994_, _36993_);
  and (_36997_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_36998_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_36999_, _36998_, _36997_);
  and (_37000_, _36999_, _36995_);
  and (_37001_, _37000_, _36992_);
  and (_37002_, _37001_, _36984_);
  and (_37003_, _37002_, _36968_);
  or (_37004_, \oc8051_golden_model_1.IRAM[5] [6], _37975_);
  or (_37005_, _04334_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_37006_, _37005_, _37004_);
  or (_37008_, \oc8051_golden_model_1.IRAM[5] [4], _37969_);
  or (_37009_, _03586_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_37010_, _37009_, _37008_);
  and (_37011_, _37010_, _37006_);
  and (_37012_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_37013_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_37014_, _37013_, _37012_);
  and (_37015_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_37016_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_37017_, _37016_, _37015_);
  and (_37019_, _37017_, _37014_);
  and (_37020_, _37019_, _37011_);
  and (_37021_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_37022_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_37023_, _37022_, _37021_);
  and (_37024_, \oc8051_golden_model_1.IRAM[5] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_37025_, \oc8051_golden_model_1.IRAM[5] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_37026_, _37025_, _37024_);
  and (_37027_, _37026_, _37023_);
  or (_37028_, _02957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_37030_, \oc8051_golden_model_1.IRAM[6] [2], _37987_);
  and (_37031_, _37030_, _37028_);
  or (_37032_, \oc8051_golden_model_1.IRAM[6] [0], _37980_);
  or (_37033_, _03926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_37034_, _37033_, _37032_);
  and (_37035_, _37034_, _37031_);
  and (_37036_, _37035_, _37027_);
  and (_37037_, _37036_, _37020_);
  nor (_37038_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_37039_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_37040_, _37039_, _37038_);
  and (_37041_, \oc8051_golden_model_1.IRAM[6] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_37042_, \oc8051_golden_model_1.IRAM[6] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_37043_, _37042_, _37041_);
  and (_37044_, _37043_, _37040_);
  or (_37045_, _04328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_37046_, \oc8051_golden_model_1.IRAM[6] [6], _37997_);
  and (_37047_, _37046_, _37045_);
  or (_37048_, _03580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_37049_, \oc8051_golden_model_1.IRAM[6] [4], _37992_);
  and (_37051_, _37049_, _37048_);
  and (_37052_, _37051_, _37047_);
  and (_37053_, _37052_, _37044_);
  and (_37054_, \oc8051_golden_model_1.IRAM[6] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_37055_, \oc8051_golden_model_1.IRAM[6] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_37056_, _37055_, _37054_);
  nor (_37057_, \oc8051_golden_model_1.IRAM[7] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_37058_, \oc8051_golden_model_1.IRAM[7] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_37059_, _37058_, _37057_);
  or (_37060_, _02955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_37062_, \oc8051_golden_model_1.IRAM[7] [2], _38009_);
  and (_37063_, _37062_, _37060_);
  and (_37064_, _37063_, _37059_);
  and (_37065_, _37064_, _37056_);
  and (_37066_, _37065_, _37053_);
  and (_37067_, _37066_, _37037_);
  and (_37068_, _37067_, _37003_);
  and (_37069_, _37068_, _36935_);
  and (_37070_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_37071_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_37073_, _37071_, _37070_);
  or (_37074_, \oc8051_golden_model_1.PSW [1], _36179_);
  or (_37075_, _23361_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_37076_, _37075_, _37074_);
  and (_37077_, _37076_, _37073_);
  or (_37078_, \oc8051_golden_model_1.PSW [4], _37436_);
  or (_37079_, _23813_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_37080_, _37079_, _37078_);
  or (_37081_, \oc8051_golden_model_1.PSW [3], _37312_);
  or (_37082_, _23699_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_37084_, _37082_, _37081_);
  and (_37085_, _37084_, _37080_);
  and (_37086_, _37085_, _37077_);
  or (_37087_, _06707_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_37088_, \oc8051_golden_model_1.PSW [7], _25218_);
  and (_37089_, _37088_, _37087_);
  and (_37090_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_37091_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_37092_, _37091_, _37090_);
  or (_37093_, \oc8051_golden_model_1.PSW [5], _36176_);
  or (_37095_, _23927_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_37096_, _37095_, _37093_);
  and (_37097_, _37096_, _37092_);
  and (_37098_, _37097_, _37089_);
  and (_37099_, _37098_, _37086_);
  or (_37100_, _37099_, property_valid_psw_1_r);
  or (_37101_, _16368_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand (_37102_, _16462_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_37103_, _37102_, _37101_);
  nor (_37104_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_37106_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_37107_, _37106_, _37104_);
  and (_37108_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_37109_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_37110_, _37109_, _37108_);
  and (_37111_, _37110_, _37107_);
  or (_37112_, _16182_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_37113_, _16368_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_37114_, _37113_, _37112_);
  or (_37115_, _15995_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_37117_, _16182_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_37118_, _37117_, _37115_);
  and (_37119_, _37118_, _37114_);
  and (_37120_, _37119_, _37111_);
  and (_37121_, \oc8051_golden_model_1.DPL [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_37122_, \oc8051_golden_model_1.DPL [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_37123_, _37122_, _37121_);
  and (_37124_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_37125_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_37126_, _37125_, _37124_);
  nand (_37127_, _07747_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_37128_, _16462_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_37129_, _37128_, _37127_);
  and (_37130_, _37129_, _37126_);
  and (_37131_, _37130_, _37123_);
  and (_37132_, _37131_, _37120_);
  and (_37133_, _37132_, _37103_);
  and (_37134_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_37135_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_37136_, _37135_, _37134_);
  and (_37138_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_37139_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_37140_, _37139_, _37138_);
  and (_37141_, _37140_, _37136_);
  or (_37142_, \oc8051_golden_model_1.IRAM[1] [2], _37871_);
  or (_37143_, _02940_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_37144_, _37143_, _37142_);
  or (_37145_, _03904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_37146_, \oc8051_golden_model_1.IRAM[1] [0], _37863_);
  and (_37147_, _37146_, _37145_);
  and (_37149_, _37147_, _37144_);
  and (_37150_, _37149_, _37141_);
  and (_37151_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nor (_37152_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_37153_, _37152_, _37151_);
  or (_37154_, _16830_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_37155_, _17016_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_37156_, _37155_, _37154_);
  and (_37157_, _37156_, _37153_);
  and (_37158_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor (_37160_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_37161_, _37160_, _37158_);
  nand (_37162_, _16830_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_37163_, _07747_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_37164_, _37163_, _37162_);
  and (_37165_, _37164_, _37161_);
  and (_37166_, _37165_, _37157_);
  and (_37167_, _37166_, _37150_);
  nor (_37168_, \oc8051_golden_model_1.DPH [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_37169_, \oc8051_golden_model_1.DPH [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_37171_, _37169_, _37168_);
  and (_37172_, \oc8051_golden_model_1.IRAM[0] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_37173_, \oc8051_golden_model_1.IRAM[0] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_37174_, _37173_, _37172_);
  and (_37175_, _37174_, _37171_);
  or (_37176_, \oc8051_golden_model_1.IRAM[0] [2], _37786_);
  or (_37177_, _02543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and (_37178_, _37177_, _37176_);
  or (_37179_, _17016_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_37180_, \oc8051_golden_model_1.IRAM[0] [0], _37747_);
  and (_37182_, _37180_, _37179_);
  and (_37183_, _37182_, _37178_);
  and (_37184_, _37183_, _37175_);
  or (_37185_, _04312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_37186_, \oc8051_golden_model_1.IRAM[0] [6], _37846_);
  and (_37187_, _37186_, _37185_);
  or (_37188_, _03564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_37189_, \oc8051_golden_model_1.IRAM[0] [4], _37817_);
  and (_37190_, _37189_, _37188_);
  and (_37191_, _37190_, _37187_);
  nor (_37193_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_37194_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_37195_, _37194_, _37193_);
  nor (_37196_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_37197_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_37198_, _37197_, _37196_);
  and (_37199_, _37198_, _37195_);
  and (_37200_, _37199_, _37191_);
  and (_37201_, _37200_, _37184_);
  and (_37202_, _37201_, _37167_);
  and (_37204_, _37202_, _37133_);
  and (_37205_, _37204_, _37100_);
  and (_37206_, _37205_, _37069_);
  and (_37207_, _37206_, _36932_);
  and (_37208_, _37207_, _36896_);
  or (_37209_, _37208_, rst);
  and (_00000_, _37209_, _00009_);
  and (_00002_[7], _40038_, _39026_);
  and (_37210_, _39632_, eq_state);
  and (_37211_, _37210_, _07599_);
  and (property_invalid_pc, _37211_, _36304_);
  buf (_00070_, _39026_);
  buf (_00120_, _39026_);
  buf (_00173_, _39026_);
  buf (_00225_, _39026_);
  buf (_00277_, _39026_);
  buf (_00329_, _39026_);
  buf (_00381_, _39026_);
  buf (_00433_, _39026_);
  buf (_00485_, _39026_);
  buf (_00537_, _39026_);
  buf (_00589_, _39026_);
  buf (_00641_, _39026_);
  buf (_00693_, _39026_);
  buf (_00745_, _39026_);
  buf (_00796_, _39026_);
  buf (_00848_, _39026_);
  buf (_03169_, _00924_);
  buf (_03172_, _00928_);
  buf (_03206_, _00924_);
  buf (_03209_, _00928_);
  buf (_05681_, _01069_);
  buf (_05683_, _01072_);
  buf (_05685_, _01075_);
  buf (_05687_, _01078_);
  buf (_05689_, _01081_);
  buf (_05691_, _01084_);
  buf (_05693_, _01087_);
  buf (_05695_, _01090_);
  buf (_05697_, _01093_);
  buf (_05699_, _01096_);
  buf (_05701_, _01099_);
  buf (_05703_, _01102_);
  buf (_05705_, _01105_);
  buf (_05707_, _01107_);
  buf (_05801_, _01069_);
  buf (_05803_, _01072_);
  buf (_05805_, _01075_);
  buf (_05807_, _01078_);
  buf (_05809_, _01081_);
  buf (_05811_, _01084_);
  buf (_05813_, _01087_);
  buf (_05815_, _01090_);
  buf (_05817_, _01093_);
  buf (_05819_, _01096_);
  buf (_05821_, _01099_);
  buf (_05823_, _01102_);
  buf (_05825_, _01105_);
  buf (_05827_, _01107_);
  buf (_08210_, _01529_);
  buf (_08313_, _01529_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00004_[0]);
  dff (p1in_reg[1], _00004_[1]);
  dff (p1in_reg[2], _00004_[2]);
  dff (p1in_reg[3], _00004_[3]);
  dff (p1in_reg[4], _00004_[4]);
  dff (p1in_reg[5], _00004_[5]);
  dff (p1in_reg[6], _00004_[6]);
  dff (p1in_reg[7], _00004_[7]);
  dff (p2in_reg[0], _00005_[0]);
  dff (p2in_reg[1], _00005_[1]);
  dff (p2in_reg[2], _00005_[2]);
  dff (p2in_reg[3], _00005_[3]);
  dff (p2in_reg[4], _00005_[4]);
  dff (p2in_reg[5], _00005_[5]);
  dff (p2in_reg[6], _00005_[6]);
  dff (p2in_reg[7], _00005_[7]);
  dff (p3in_reg[0], _00006_[0]);
  dff (p3in_reg[1], _00006_[1]);
  dff (p3in_reg[2], _00006_[2]);
  dff (p3in_reg[3], _00006_[3]);
  dff (p3in_reg[4], _00006_[4]);
  dff (p3in_reg[5], _00006_[5]);
  dff (p3in_reg[6], _00006_[6]);
  dff (p3in_reg[7], _00006_[7]);
  dff (inst_finished_r, _00001_);
  dff (regs_always_zero, _00009_);
  dff (property_valid_psw_1_r, _00007_);
  dff (property_valid_sp_1_r, _00008_);
  dff (p1_valid_r, _00003_);
  dff (eq_state, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _00098_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _00100_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _00102_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _00104_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _00106_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _00108_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _00110_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _00067_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _00070_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _00150_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _00152_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _00154_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _00156_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _00158_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _00160_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _00162_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _00117_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _00120_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00618_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00620_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00622_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00624_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00626_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00628_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00630_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00586_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00589_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00670_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00672_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00674_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00676_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00678_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00680_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00682_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00638_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00641_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00722_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00724_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00726_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00728_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00730_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00732_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00734_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00690_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00693_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00774_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00776_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00778_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00780_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00782_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00784_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00786_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00742_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00745_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _00826_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _00828_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _00829_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _00831_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _00833_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _00835_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _00837_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _00794_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00796_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _00877_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _00879_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _00881_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _00883_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _00885_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _00887_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _00889_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _00845_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _00848_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _00203_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _00205_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _00207_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00209_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00211_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00213_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00215_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _00170_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _00173_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00255_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00257_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00258_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00260_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00262_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00264_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00266_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00223_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00225_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00306_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00308_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00310_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00312_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00314_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00316_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00318_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00274_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00277_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00358_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00360_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00362_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00364_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00366_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00368_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00370_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00326_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00329_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00410_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00412_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00414_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00416_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00418_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00420_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00422_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00378_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00381_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00462_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00464_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00466_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00468_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00470_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00472_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00474_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00430_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00433_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00514_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00516_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00518_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00520_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00522_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00524_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00526_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00482_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00485_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00566_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00568_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00570_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00572_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00574_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00576_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00578_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00534_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00537_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _38817_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _38819_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _38820_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _38821_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _38822_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _38823_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _38825_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _38581_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _38806_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _38808_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _38809_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _38810_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _38811_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _38812_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _38814_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _38815_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _38795_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _38797_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _38798_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _38799_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _38800_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _38801_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _38802_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _38803_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _38783_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _38784_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _38786_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _38787_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _38788_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _38789_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _38790_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _38792_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _38772_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _38773_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _38774_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _38776_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _38777_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _38778_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _38779_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _38780_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _38761_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _38762_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _38763_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _38764_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _38765_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _38766_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _38767_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _38768_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _38749_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _38750_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _38751_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _38752_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _38754_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _38755_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _38756_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _38757_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _38738_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _38739_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _38740_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _38741_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _38742_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _38744_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _38745_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _38746_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _38726_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _38727_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _38728_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _38730_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _38731_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _38732_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _38733_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _38734_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _38714_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _38715_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _38716_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _38717_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _38719_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _38720_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _38721_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _38722_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _38703_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _38704_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _38705_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _38706_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _38708_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _38709_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _38710_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _38711_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _38692_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _38693_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _38694_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _38695_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _38696_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _38698_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _38699_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _38700_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _38680_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _38681_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _38682_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _38683_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _38684_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _38685_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _38686_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _38687_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _38668_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _38669_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _38670_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _38671_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _38672_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _38674_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _38675_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _38676_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _38656_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _38657_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _38658_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _38660_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _38661_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _38662_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _38663_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _38664_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _38643_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _38644_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _38646_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _38647_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _38649_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _38650_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _38651_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _38652_);
  dff (\oc8051_golden_model_1.B [0], _41617_);
  dff (\oc8051_golden_model_1.B [1], _41618_);
  dff (\oc8051_golden_model_1.B [2], _41619_);
  dff (\oc8051_golden_model_1.B [3], _41620_);
  dff (\oc8051_golden_model_1.B [4], _41621_);
  dff (\oc8051_golden_model_1.B [5], _41622_);
  dff (\oc8051_golden_model_1.B [6], _41623_);
  dff (\oc8051_golden_model_1.B [7], _38582_);
  dff (\oc8051_golden_model_1.ACC [0], _41625_);
  dff (\oc8051_golden_model_1.ACC [1], _41626_);
  dff (\oc8051_golden_model_1.ACC [2], _41627_);
  dff (\oc8051_golden_model_1.ACC [3], _41628_);
  dff (\oc8051_golden_model_1.ACC [4], _41629_);
  dff (\oc8051_golden_model_1.ACC [5], _41630_);
  dff (\oc8051_golden_model_1.ACC [6], _41632_);
  dff (\oc8051_golden_model_1.ACC [7], _38583_);
  dff (\oc8051_golden_model_1.DPL [0], _41633_);
  dff (\oc8051_golden_model_1.DPL [1], _41634_);
  dff (\oc8051_golden_model_1.DPL [2], _41636_);
  dff (\oc8051_golden_model_1.DPL [3], _41637_);
  dff (\oc8051_golden_model_1.DPL [4], _41638_);
  dff (\oc8051_golden_model_1.DPL [5], _41639_);
  dff (\oc8051_golden_model_1.DPL [6], _41640_);
  dff (\oc8051_golden_model_1.DPL [7], _38584_);
  dff (\oc8051_golden_model_1.DPH [0], _41642_);
  dff (\oc8051_golden_model_1.DPH [1], _41643_);
  dff (\oc8051_golden_model_1.DPH [2], _41644_);
  dff (\oc8051_golden_model_1.DPH [3], _41645_);
  dff (\oc8051_golden_model_1.DPH [4], _41646_);
  dff (\oc8051_golden_model_1.DPH [5], _41647_);
  dff (\oc8051_golden_model_1.DPH [6], _41648_);
  dff (\oc8051_golden_model_1.DPH [7], _38586_);
  dff (\oc8051_golden_model_1.IE [0], _41650_);
  dff (\oc8051_golden_model_1.IE [1], _41651_);
  dff (\oc8051_golden_model_1.IE [2], _41652_);
  dff (\oc8051_golden_model_1.IE [3], _41653_);
  dff (\oc8051_golden_model_1.IE [4], _41655_);
  dff (\oc8051_golden_model_1.IE [5], _41656_);
  dff (\oc8051_golden_model_1.IE [6], _41657_);
  dff (\oc8051_golden_model_1.IE [7], _38587_);
  dff (\oc8051_golden_model_1.IP [0], _41659_);
  dff (\oc8051_golden_model_1.IP [1], _41660_);
  dff (\oc8051_golden_model_1.IP [2], _41661_);
  dff (\oc8051_golden_model_1.IP [3], _41662_);
  dff (\oc8051_golden_model_1.IP [4], _41663_);
  dff (\oc8051_golden_model_1.IP [5], _41664_);
  dff (\oc8051_golden_model_1.IP [6], _41665_);
  dff (\oc8051_golden_model_1.IP [7], _38588_);
  dff (\oc8051_golden_model_1.P0 [0], _41667_);
  dff (\oc8051_golden_model_1.P0 [1], _41668_);
  dff (\oc8051_golden_model_1.P0 [2], _41669_);
  dff (\oc8051_golden_model_1.P0 [3], _41670_);
  dff (\oc8051_golden_model_1.P0 [4], _41671_);
  dff (\oc8051_golden_model_1.P0 [5], _41672_);
  dff (\oc8051_golden_model_1.P0 [6], _41674_);
  dff (\oc8051_golden_model_1.P0 [7], _38589_);
  dff (\oc8051_golden_model_1.P1 [0], _41675_);
  dff (\oc8051_golden_model_1.P1 [1], _41676_);
  dff (\oc8051_golden_model_1.P1 [2], _41678_);
  dff (\oc8051_golden_model_1.P1 [3], _41679_);
  dff (\oc8051_golden_model_1.P1 [4], _41680_);
  dff (\oc8051_golden_model_1.P1 [5], _41681_);
  dff (\oc8051_golden_model_1.P1 [6], _41682_);
  dff (\oc8051_golden_model_1.P1 [7], _38590_);
  dff (\oc8051_golden_model_1.P2 [0], _41684_);
  dff (\oc8051_golden_model_1.P2 [1], _41685_);
  dff (\oc8051_golden_model_1.P2 [2], _41686_);
  dff (\oc8051_golden_model_1.P2 [3], _41687_);
  dff (\oc8051_golden_model_1.P2 [4], _41688_);
  dff (\oc8051_golden_model_1.P2 [5], _41689_);
  dff (\oc8051_golden_model_1.P2 [6], _41690_);
  dff (\oc8051_golden_model_1.P2 [7], _38592_);
  dff (\oc8051_golden_model_1.P3 [0], _41692_);
  dff (\oc8051_golden_model_1.P3 [1], _41693_);
  dff (\oc8051_golden_model_1.P3 [2], _41694_);
  dff (\oc8051_golden_model_1.P3 [3], _41695_);
  dff (\oc8051_golden_model_1.P3 [4], _41697_);
  dff (\oc8051_golden_model_1.P3 [5], _41698_);
  dff (\oc8051_golden_model_1.P3 [6], _41699_);
  dff (\oc8051_golden_model_1.P3 [7], _38593_);
  dff (\oc8051_golden_model_1.PSW [0], _41701_);
  dff (\oc8051_golden_model_1.PSW [1], _41702_);
  dff (\oc8051_golden_model_1.PSW [2], _41703_);
  dff (\oc8051_golden_model_1.PSW [3], _41704_);
  dff (\oc8051_golden_model_1.PSW [4], _41705_);
  dff (\oc8051_golden_model_1.PSW [5], _41706_);
  dff (\oc8051_golden_model_1.PSW [6], _41707_);
  dff (\oc8051_golden_model_1.PSW [7], _38594_);
  dff (\oc8051_golden_model_1.PCON [0], _41709_);
  dff (\oc8051_golden_model_1.PCON [1], _41710_);
  dff (\oc8051_golden_model_1.PCON [2], _41711_);
  dff (\oc8051_golden_model_1.PCON [3], _41712_);
  dff (\oc8051_golden_model_1.PCON [4], _41713_);
  dff (\oc8051_golden_model_1.PCON [5], _41714_);
  dff (\oc8051_golden_model_1.PCON [6], _41715_);
  dff (\oc8051_golden_model_1.PCON [7], _38595_);
  dff (\oc8051_golden_model_1.SBUF [0], _41716_);
  dff (\oc8051_golden_model_1.SBUF [1], _41717_);
  dff (\oc8051_golden_model_1.SBUF [2], _41719_);
  dff (\oc8051_golden_model_1.SBUF [3], _41720_);
  dff (\oc8051_golden_model_1.SBUF [4], _41721_);
  dff (\oc8051_golden_model_1.SBUF [5], _41722_);
  dff (\oc8051_golden_model_1.SBUF [6], _41723_);
  dff (\oc8051_golden_model_1.SBUF [7], _38596_);
  dff (\oc8051_golden_model_1.SCON [0], _41725_);
  dff (\oc8051_golden_model_1.SCON [1], _41726_);
  dff (\oc8051_golden_model_1.SCON [2], _41727_);
  dff (\oc8051_golden_model_1.SCON [3], _41728_);
  dff (\oc8051_golden_model_1.SCON [4], _41729_);
  dff (\oc8051_golden_model_1.SCON [5], _41730_);
  dff (\oc8051_golden_model_1.SCON [6], _41731_);
  dff (\oc8051_golden_model_1.SCON [7], _38597_);
  dff (\oc8051_golden_model_1.SP [0], _41733_);
  dff (\oc8051_golden_model_1.SP [1], _41734_);
  dff (\oc8051_golden_model_1.SP [2], _41735_);
  dff (\oc8051_golden_model_1.SP [3], _41736_);
  dff (\oc8051_golden_model_1.SP [4], _41738_);
  dff (\oc8051_golden_model_1.SP [5], _41739_);
  dff (\oc8051_golden_model_1.SP [6], _41740_);
  dff (\oc8051_golden_model_1.SP [7], _38598_);
  dff (\oc8051_golden_model_1.TCON [0], _41742_);
  dff (\oc8051_golden_model_1.TCON [1], _41743_);
  dff (\oc8051_golden_model_1.TCON [2], _41744_);
  dff (\oc8051_golden_model_1.TCON [3], _41745_);
  dff (\oc8051_golden_model_1.TCON [4], _41746_);
  dff (\oc8051_golden_model_1.TCON [5], _41747_);
  dff (\oc8051_golden_model_1.TCON [6], _41748_);
  dff (\oc8051_golden_model_1.TCON [7], _38599_);
  dff (\oc8051_golden_model_1.TH0 [0], _41750_);
  dff (\oc8051_golden_model_1.TH0 [1], _41751_);
  dff (\oc8051_golden_model_1.TH0 [2], _41752_);
  dff (\oc8051_golden_model_1.TH0 [3], _41753_);
  dff (\oc8051_golden_model_1.TH0 [4], _41754_);
  dff (\oc8051_golden_model_1.TH0 [5], _41755_);
  dff (\oc8051_golden_model_1.TH0 [6], _41757_);
  dff (\oc8051_golden_model_1.TH0 [7], _38600_);
  dff (\oc8051_golden_model_1.TH1 [0], _41758_);
  dff (\oc8051_golden_model_1.TH1 [1], _41759_);
  dff (\oc8051_golden_model_1.TH1 [2], _41761_);
  dff (\oc8051_golden_model_1.TH1 [3], _41762_);
  dff (\oc8051_golden_model_1.TH1 [4], _41763_);
  dff (\oc8051_golden_model_1.TH1 [5], _41764_);
  dff (\oc8051_golden_model_1.TH1 [6], _41765_);
  dff (\oc8051_golden_model_1.TH1 [7], _38601_);
  dff (\oc8051_golden_model_1.TL0 [0], _41767_);
  dff (\oc8051_golden_model_1.TL0 [1], _41768_);
  dff (\oc8051_golden_model_1.TL0 [2], _41769_);
  dff (\oc8051_golden_model_1.TL0 [3], _41770_);
  dff (\oc8051_golden_model_1.TL0 [4], _41771_);
  dff (\oc8051_golden_model_1.TL0 [5], _41772_);
  dff (\oc8051_golden_model_1.TL0 [6], _41773_);
  dff (\oc8051_golden_model_1.TL0 [7], _38603_);
  dff (\oc8051_golden_model_1.TL1 [0], _41775_);
  dff (\oc8051_golden_model_1.TL1 [1], _41776_);
  dff (\oc8051_golden_model_1.TL1 [2], _41777_);
  dff (\oc8051_golden_model_1.TL1 [3], _41778_);
  dff (\oc8051_golden_model_1.TL1 [4], _41780_);
  dff (\oc8051_golden_model_1.TL1 [5], _41781_);
  dff (\oc8051_golden_model_1.TL1 [6], _41782_);
  dff (\oc8051_golden_model_1.TL1 [7], _38604_);
  dff (\oc8051_golden_model_1.TMOD [0], _41784_);
  dff (\oc8051_golden_model_1.TMOD [1], _41785_);
  dff (\oc8051_golden_model_1.TMOD [2], _41786_);
  dff (\oc8051_golden_model_1.TMOD [3], _41787_);
  dff (\oc8051_golden_model_1.TMOD [4], _41788_);
  dff (\oc8051_golden_model_1.TMOD [5], _41789_);
  dff (\oc8051_golden_model_1.TMOD [6], _41790_);
  dff (\oc8051_golden_model_1.TMOD [7], _38605_);
  dff (\oc8051_golden_model_1.PC [0], _41793_);
  dff (\oc8051_golden_model_1.PC [1], _41794_);
  dff (\oc8051_golden_model_1.PC [2], _41795_);
  dff (\oc8051_golden_model_1.PC [3], _41796_);
  dff (\oc8051_golden_model_1.PC [4], _41797_);
  dff (\oc8051_golden_model_1.PC [5], _41798_);
  dff (\oc8051_golden_model_1.PC [6], _41799_);
  dff (\oc8051_golden_model_1.PC [7], _41800_);
  dff (\oc8051_golden_model_1.PC [8], _41802_);
  dff (\oc8051_golden_model_1.PC [9], _41803_);
  dff (\oc8051_golden_model_1.PC [10], _41804_);
  dff (\oc8051_golden_model_1.PC [11], _41805_);
  dff (\oc8051_golden_model_1.PC [12], _41806_);
  dff (\oc8051_golden_model_1.PC [13], _41807_);
  dff (\oc8051_golden_model_1.PC [14], _41808_);
  dff (\oc8051_golden_model_1.PC [15], _38606_);
  dff (\oc8051_golden_model_1.P0INREG [0], _41810_);
  dff (\oc8051_golden_model_1.P0INREG [1], _41811_);
  dff (\oc8051_golden_model_1.P0INREG [2], _41812_);
  dff (\oc8051_golden_model_1.P0INREG [3], _41813_);
  dff (\oc8051_golden_model_1.P0INREG [4], _41814_);
  dff (\oc8051_golden_model_1.P0INREG [5], _41815_);
  dff (\oc8051_golden_model_1.P0INREG [6], _41817_);
  dff (\oc8051_golden_model_1.P0INREG [7], _38607_);
  dff (\oc8051_golden_model_1.P1INREG [0], _41818_);
  dff (\oc8051_golden_model_1.P1INREG [1], _41819_);
  dff (\oc8051_golden_model_1.P1INREG [2], _41821_);
  dff (\oc8051_golden_model_1.P1INREG [3], _41822_);
  dff (\oc8051_golden_model_1.P1INREG [4], _41823_);
  dff (\oc8051_golden_model_1.P1INREG [5], _41824_);
  dff (\oc8051_golden_model_1.P1INREG [6], _41825_);
  dff (\oc8051_golden_model_1.P1INREG [7], _38609_);
  dff (\oc8051_golden_model_1.P2INREG [0], _41827_);
  dff (\oc8051_golden_model_1.P2INREG [1], _41828_);
  dff (\oc8051_golden_model_1.P2INREG [2], _41829_);
  dff (\oc8051_golden_model_1.P2INREG [3], _41830_);
  dff (\oc8051_golden_model_1.P2INREG [4], _41831_);
  dff (\oc8051_golden_model_1.P2INREG [5], _41832_);
  dff (\oc8051_golden_model_1.P2INREG [6], _41833_);
  dff (\oc8051_golden_model_1.P2INREG [7], _38610_);
  dff (\oc8051_golden_model_1.P3INREG [0], _41835_);
  dff (\oc8051_golden_model_1.P3INREG [1], _41836_);
  dff (\oc8051_golden_model_1.P3INREG [2], _41837_);
  dff (\oc8051_golden_model_1.P3INREG [3], _41838_);
  dff (\oc8051_golden_model_1.P3INREG [4], _41840_);
  dff (\oc8051_golden_model_1.P3INREG [5], _41841_);
  dff (\oc8051_golden_model_1.P3INREG [6], _41842_);
  dff (\oc8051_golden_model_1.P3INREG [7], _38611_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _01049_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _01052_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _01055_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _01058_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _01060_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _01063_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _01066_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _00920_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _01069_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _01072_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _01075_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _01078_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _01081_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _01084_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _01087_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _00924_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _01090_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _01093_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _01096_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _01099_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _01102_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _01105_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _01107_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00928_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _37213_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _12321_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _37214_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _12324_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _37215_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _37216_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _12327_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _37217_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _37218_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _12329_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _37219_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _12332_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _37220_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _37221_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _37222_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _12335_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _37224_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _12337_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _12340_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12382_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12384_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _12308_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12387_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _12389_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _12311_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _12392_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _12313_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _12395_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _12397_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _12400_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _12403_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _12405_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _12408_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _12411_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _12316_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _12319_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _08210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _03627_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _03629_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _03631_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _03633_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _03635_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _03637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _03639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _03641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _03643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _03645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _03647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _03649_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _03651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _03653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _03655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _02773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _03687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _03689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _03691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _03693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _03695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _03697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _03699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _03701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _03703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _03705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _03707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _03709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _03711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _03713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _03715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _02777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _05587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _05589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _05591_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _05593_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _05595_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _05597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _05599_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _05601_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _05603_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _05605_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _05607_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _05609_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _05611_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _05613_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _05615_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _05617_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _05619_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _05621_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _05623_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _05625_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _05627_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _05629_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _05631_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _05633_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _05635_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _05637_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _05639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _05641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _05643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _05645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _05647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _03155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _05650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _05653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _05656_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _05658_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _05661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _05664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _05667_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _05670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _05673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _05676_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _05679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _05681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _05683_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _05685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _05687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _05689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _05691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _05693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _05695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _05697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _05699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _05701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _05703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _05705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _05707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _03172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _03175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _05709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _05711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _05713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _05715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _05717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _05719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _05721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _03182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _05723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _05725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _05727_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _05729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _05731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _05733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _05735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _05737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _05739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _05741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _05743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _05745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _05747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _05749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _05751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _05753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _05755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _05757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _05759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _05761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _05763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _05765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _05767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _05769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _05771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _05773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _05775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _05777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _05779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _05781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _03193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _05783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _05785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _05789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _05791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _05793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _05797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _05799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _05801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _05803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _05805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _05807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _05809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _05811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _05813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _03206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _05815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _05817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _05819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _05821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _05823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _05825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _05827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _03209_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _03212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _05829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _05831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _05833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _05835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _05837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _05839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _05841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03217_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _05843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _05845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _05847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03223_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _05849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _05851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _05853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _05855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _05857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _05859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _05861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _05863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _05865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _05867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _05869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _05871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _05873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _05875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _05877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _05879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _05881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _05883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _05885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _05887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _05889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _05891_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _05893_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _05895_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _05897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _05899_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _05901_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _05903_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _05905_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _05907_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _05909_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _03228_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _05911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _05913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _05915_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _05917_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _05919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _05921_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _05923_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _03230_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _03232_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _03234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _05925_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _05927_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _05929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _05931_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _05933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _05935_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _05937_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _05939_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _05941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _05943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _05945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _05947_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _05949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _05951_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _05953_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _03236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03238_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03240_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _05955_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _05957_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _05959_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _05961_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _05963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _05965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _05967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _05969_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _05971_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _05973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _05975_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _05977_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _05979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _05981_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _05983_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _03244_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _03246_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _08307_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _08467_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _08469_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _08471_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _08473_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _08475_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _08477_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _08479_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _08310_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _08313_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _08481_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _08483_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _08316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _40438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _40441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _40445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _40451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _40457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _40463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _40469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _40472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _40515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _40519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _40523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _40527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _40531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _40535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _40539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _40542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _40711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _40715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _40719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _40723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _40727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _40731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _40735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _40738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _40676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _40680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _40684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _40688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _40692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _40696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _40700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _40703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _40644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _40648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _40652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _40656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _40660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _40664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _40668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _40671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _40612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _40616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _40620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _40624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _40628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _40632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _40636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _40639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _40580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _40584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _40588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _40592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _40596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _40600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _40604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _40607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _40548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _40552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _40556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _40560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _40564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _40568_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _40572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _40574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _40480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _40484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _40488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _40492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _40496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _40500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _40504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _40507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _40743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _40747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _40751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _40755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _40759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _40763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _40767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _40770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _40903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _40907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _40911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _40915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _40919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _40923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _40927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _40930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _40871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _40875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _40879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _40883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _40887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _40891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _40895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _40898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _40839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _40843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _40847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _40851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _40855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _40859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _40863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _40866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _40806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _40810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _40814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _40818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _40822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _40826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _40830_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _40833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _40775_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _40779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _40783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _40787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _40791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _40795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _40799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _40801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _40935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _40939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _40943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _40947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _40951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _40955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _40959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _40157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _00048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _00050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _00052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _00053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _00055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _00057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _00059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _40145_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _01522_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _01524_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _02205_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _02207_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _02209_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _02211_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _02213_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _02215_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _02217_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _01526_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _01529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _08869_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _08880_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _08891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _08902_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _08913_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _08924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _08935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _07163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _29071_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _29180_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _29289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _29398_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _29507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _29616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _29725_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _41219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _41228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _41236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _41245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _41254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _41263_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _41272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _40187_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _41280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _41289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _41297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _41306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _41314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _41323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _41331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _40208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _39026_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _40001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _40003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _40005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _40007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _40009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _40011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _40013_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _38993_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _40015_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _39028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _38995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _39030_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _38997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _40025_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _39031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _39033_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _39017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _39019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _39020_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _39022_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _40029_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _40031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _40033_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _40035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _40037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _40039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _40041_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _40043_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _40045_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _40047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _38937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _40049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _40051_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _40053_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _40055_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _40057_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _40059_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _40061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _38973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _38290_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _38292_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _38294_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _38296_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _38298_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _38300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _38302_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _19308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _38304_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _38306_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _38308_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _38310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _38312_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _38314_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _38316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _19330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _38318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _38320_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _38322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _38324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _38326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _38328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _38329_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _19353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _38331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _38333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _38335_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _38337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _38339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _38341_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _38343_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _19376_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06399_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _06410_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _06432_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _06443_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _01572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _38077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _38086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _38094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _38103_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _38111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _38119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _38128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _35488_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _35268_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [8], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [9], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [10], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [11], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [12], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [13], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [14], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [15], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_data_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_comp1.des [0], ABINPUT[27]);
  buf(\oc8051_top_1.oc8051_comp1.des [1], ABINPUT[28]);
  buf(\oc8051_top_1.oc8051_comp1.des [2], ABINPUT[29]);
  buf(\oc8051_top_1.oc8051_comp1.des [3], ABINPUT[30]);
  buf(\oc8051_top_1.oc8051_comp1.des [4], ABINPUT[31]);
  buf(\oc8051_top_1.oc8051_comp1.des [5], ABINPUT[32]);
  buf(\oc8051_top_1.oc8051_comp1.des [6], ABINPUT[33]);
  buf(\oc8051_top_1.oc8051_comp1.des [7], ABINPUT[34]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1046 , \oc8051_golden_model_1.n1047 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1063 , \oc8051_golden_model_1.n1064 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1157 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1157 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1157 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1157 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1159 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1167 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1214 , \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1265 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1276 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1284 [0]);
  buf(\oc8051_golden_model_1.n1284 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1284 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1284 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1284 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1284 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1284 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1284 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1300 , \oc8051_golden_model_1.n1301 [0]);
  buf(\oc8051_golden_model_1.n1301 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1301 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1301 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1301 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1301 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1301 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1360 , \oc8051_golden_model_1.n1361 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1367 [8], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1374 [4], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1375 , \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1384 , \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.n1402 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.n1402 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.n1402 [7]);
  buf(\oc8051_golden_model_1.n1401 , \oc8051_golden_model_1.n1402 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1424 [8], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1425 , \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1430 [4], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1431 , \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1439 , \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1440 [2], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1440 [6], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1440 [7], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.n1457 [2]);
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.n1457 [6]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.n1457 [7]);
  buf(\oc8051_golden_model_1.n1456 , \oc8051_golden_model_1.n1457 [0]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1459 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1459 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1461 [8], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1462 , \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1463 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1463 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1463 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1463 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1464 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1464 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1464 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1464 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1466 [4], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1467 , \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1468 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n1468 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n1468 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n1468 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n1468 [4], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n1468 [5], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n1468 [6], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n1468 [7], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1468 [8], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n1475 , \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1477 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1477 [1], \oc8051_golden_model_1.n1493 [2]);
  buf(\oc8051_golden_model_1.n1477 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1477 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1477 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1477 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1477 [6], \oc8051_golden_model_1.n1493 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.n1507 [0]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1496 [8], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1497 , \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1504 , \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.n1507 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.n1507 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.n1507 [7]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1509 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1511 [8], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1513 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1516 , \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1517 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1517 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1517 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1517 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1517 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1517 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1517 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1517 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1524 , \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1525 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1525 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1525 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1546 [7], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.n1548 [2]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.n1548 [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1559 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1559 [6], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1559 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1560 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1560 [5], \oc8051_golden_model_1.n1561 [6]);
  buf(\oc8051_golden_model_1.n1560 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1561 [0], \oc8051_golden_model_1.n1564 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1562 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1562 [2], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1562 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1562 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1562 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1562 [6], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1562 [7], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1563 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1563 [1], \oc8051_golden_model_1.n1564 [2]);
  buf(\oc8051_golden_model_1.n1563 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1563 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1563 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1563 [5], \oc8051_golden_model_1.n1564 [6]);
  buf(\oc8051_golden_model_1.n1563 [6], \oc8051_golden_model_1.n1564 [7]);
  buf(\oc8051_golden_model_1.n1564 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1564 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1564 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1564 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1567 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1568 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1568 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1568 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1568 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1568 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1568 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1568 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1573 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1575 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1577 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1586 , \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1587 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1588 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1591 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1593 [8], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1594 , \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1595 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1595 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1597 [4], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1598 , \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1605 , \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1606 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1606 [2], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1606 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1606 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1606 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1606 [6], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1606 [7], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1607 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1607 [1], \oc8051_golden_model_1.n1623 [2]);
  buf(\oc8051_golden_model_1.n1607 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1607 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1607 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [5], \oc8051_golden_model_1.n1623 [6]);
  buf(\oc8051_golden_model_1.n1607 [6], \oc8051_golden_model_1.n1623 [7]);
  buf(\oc8051_golden_model_1.n1622 , \oc8051_golden_model_1.n1623 [0]);
  buf(\oc8051_golden_model_1.n1623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1627 [8], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1628 , \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1630 [4], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1631 , \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1638 , \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1639 [2], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1639 [6], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1639 [7], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1640 [1], \oc8051_golden_model_1.n1656 [2]);
  buf(\oc8051_golden_model_1.n1640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [5], \oc8051_golden_model_1.n1656 [6]);
  buf(\oc8051_golden_model_1.n1640 [6], \oc8051_golden_model_1.n1656 [7]);
  buf(\oc8051_golden_model_1.n1655 , \oc8051_golden_model_1.n1656 [0]);
  buf(\oc8051_golden_model_1.n1656 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1656 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1656 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1656 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1660 [8], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1664 , \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1672 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1672 [2], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1672 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1672 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1672 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1672 [6], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1672 [7], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1673 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1673 [1], \oc8051_golden_model_1.n1689 [2]);
  buf(\oc8051_golden_model_1.n1673 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1673 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1673 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [5], \oc8051_golden_model_1.n1689 [6]);
  buf(\oc8051_golden_model_1.n1673 [6], \oc8051_golden_model_1.n1689 [7]);
  buf(\oc8051_golden_model_1.n1688 , \oc8051_golden_model_1.n1689 [0]);
  buf(\oc8051_golden_model_1.n1689 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1689 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1689 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1689 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1693 [8], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1694 , \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1697 , \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [2], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1705 [6], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1705 [7], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1706 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1706 [1], \oc8051_golden_model_1.n1722 [2]);
  buf(\oc8051_golden_model_1.n1706 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1706 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1706 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1706 [5], \oc8051_golden_model_1.n1722 [6]);
  buf(\oc8051_golden_model_1.n1706 [6], \oc8051_golden_model_1.n1722 [7]);
  buf(\oc8051_golden_model_1.n1721 , \oc8051_golden_model_1.n1722 [0]);
  buf(\oc8051_golden_model_1.n1722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1747 [2], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1747 [6], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1747 [7], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1748 [0], \oc8051_golden_model_1.n1749 [1]);
  buf(\oc8051_golden_model_1.n1748 [1], \oc8051_golden_model_1.n1749 [2]);
  buf(\oc8051_golden_model_1.n1748 [2], \oc8051_golden_model_1.n1749 [3]);
  buf(\oc8051_golden_model_1.n1748 [3], \oc8051_golden_model_1.n1749 [4]);
  buf(\oc8051_golden_model_1.n1748 [4], \oc8051_golden_model_1.n1749 [5]);
  buf(\oc8051_golden_model_1.n1748 [5], \oc8051_golden_model_1.n1749 [6]);
  buf(\oc8051_golden_model_1.n1748 [6], \oc8051_golden_model_1.n1749 [7]);
  buf(\oc8051_golden_model_1.n1749 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1805 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1821 , \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.n1822 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1822 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1822 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1822 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1822 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1822 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1822 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1838 , \oc8051_golden_model_1.n1839 [0]);
  buf(\oc8051_golden_model_1.n1839 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1839 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1839 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1839 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1839 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1839 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1839 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1855 , \oc8051_golden_model_1.n1856 [0]);
  buf(\oc8051_golden_model_1.n1856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1879 [1], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1879 [2], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1879 [3], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1879 [4], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1879 [5], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1879 [6], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1879 [7], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1880 [0], \oc8051_golden_model_1.n1881 [1]);
  buf(\oc8051_golden_model_1.n1880 [1], \oc8051_golden_model_1.n1881 [2]);
  buf(\oc8051_golden_model_1.n1880 [2], \oc8051_golden_model_1.n1881 [3]);
  buf(\oc8051_golden_model_1.n1880 [3], \oc8051_golden_model_1.n1881 [4]);
  buf(\oc8051_golden_model_1.n1880 [4], \oc8051_golden_model_1.n1881 [5]);
  buf(\oc8051_golden_model_1.n1880 [5], \oc8051_golden_model_1.n1881 [6]);
  buf(\oc8051_golden_model_1.n1880 [6], \oc8051_golden_model_1.n1881 [7]);
  buf(\oc8051_golden_model_1.n1881 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n1936 , \oc8051_golden_model_1.n1937 [0]);
  buf(\oc8051_golden_model_1.n1937 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1937 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1937 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1937 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1937 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1937 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1937 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1953 , \oc8051_golden_model_1.n1954 [0]);
  buf(\oc8051_golden_model_1.n1954 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1954 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1954 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1954 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1954 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1954 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1954 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1970 , \oc8051_golden_model_1.n1971 [0]);
  buf(\oc8051_golden_model_1.n1971 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1971 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1971 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1971 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1971 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1971 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1971 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1987 , \oc8051_golden_model_1.n1988 [0]);
  buf(\oc8051_golden_model_1.n1988 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1988 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1988 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1988 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1988 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1988 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1988 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2085 , \oc8051_golden_model_1.n2086 [0]);
  buf(\oc8051_golden_model_1.n2086 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2086 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2086 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2086 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2086 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2086 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2102 , \oc8051_golden_model_1.n2103 [0]);
  buf(\oc8051_golden_model_1.n2103 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2103 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2103 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2103 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2103 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2103 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2119 , \oc8051_golden_model_1.n2120 [0]);
  buf(\oc8051_golden_model_1.n2120 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2120 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2120 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2120 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2120 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2136 , \oc8051_golden_model_1.n2137 [0]);
  buf(\oc8051_golden_model_1.n2137 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2137 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2137 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2137 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2137 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2137 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2137 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2141 , \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2142 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2142 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2142 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2142 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2142 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2142 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2143 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2143 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2143 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2143 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2143 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [7], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2144 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2144 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2144 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2144 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2144 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2144 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2144 [6], \oc8051_golden_model_1.n2145 [7]);
  buf(\oc8051_golden_model_1.n2145 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2145 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2145 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2145 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2145 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2145 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2160 , \oc8051_golden_model_1.n2161 [0]);
  buf(\oc8051_golden_model_1.n2161 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2161 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2161 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2161 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2161 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2161 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2200 , \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2201 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2201 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2201 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2201 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2201 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2201 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2201 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2201 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2202 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2202 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2202 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2202 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2202 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2202 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2202 [6], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2203 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2203 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2203 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2203 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2203 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2203 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2203 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2210 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2210 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2210 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2210 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2211 , \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2212 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2212 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2212 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2212 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2212 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2212 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2213 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2213 [1], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2213 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2213 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2213 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2213 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2213 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2228 , \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.n2229 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2229 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2229 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2229 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2229 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2229 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2444 , \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2446 , \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2452 , \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2453 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2453 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2453 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2453 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2453 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2453 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2454 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2454 [1], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2454 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2454 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2454 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 [5], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2454 [6], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2474 , \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2476 , \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2482 , \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2483 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2483 [2], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2483 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2483 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2483 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2483 [6], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2483 [7], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2484 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2484 [1], \oc8051_golden_model_1.n2500 [2]);
  buf(\oc8051_golden_model_1.n2484 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2484 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2484 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2484 [5], \oc8051_golden_model_1.n2500 [6]);
  buf(\oc8051_golden_model_1.n2484 [6], \oc8051_golden_model_1.n2500 [7]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2504 , \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2512 , \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2513 [2], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2513 [6], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2513 [7], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2514 [1], \oc8051_golden_model_1.n2530 [2]);
  buf(\oc8051_golden_model_1.n2514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 [5], \oc8051_golden_model_1.n2530 [6]);
  buf(\oc8051_golden_model_1.n2514 [6], \oc8051_golden_model_1.n2530 [7]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.n2530 [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2534 , \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.n2560 [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.n2560 [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.n2560 [7]);
  buf(\oc8051_golden_model_1.n2559 , \oc8051_golden_model_1.n2560 [0]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2564 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2564 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2564 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2564 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2564 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2564 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2564 [6], \oc8051_golden_model_1.n2565 [7]);
  buf(\oc8051_golden_model_1.n2565 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2565 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2565 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2565 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2565 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2565 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2565 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], \oc8051_golden_model_1.n2568 [7]);
  buf(\oc8051_golden_model_1.n2568 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2568 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2568 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2568 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2568 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2568 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2568 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2572 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2572 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2572 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2572 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2572 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2572 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2572 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2572 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2572 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.n2596 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2596 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2596 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2596 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2596 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2596 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2600 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2600 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2600 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2600 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2600 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2600 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2600 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2600 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2601 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2601 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2601 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2601 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2601 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2601 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2601 [6], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2602 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2602 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2602 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2602 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2602 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2602 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2602 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2666 , \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2667 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2667 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2667 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2667 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2667 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2667 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2667 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2667 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2669 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2696 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2696 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2698 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2698 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2698 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2698 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2698 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2698 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2702 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2703 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2705 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2706 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2713 , \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2734 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2734 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2734 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2734 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2734 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2734 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2734 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2735 [0], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2735 [1], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2735 [2], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2735 [3], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2735 [4], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2735 [5], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2735 [6], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2750 , \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.n2751 [1], \oc8051_golden_model_1.n2914 [1]);
  buf(\oc8051_golden_model_1.n2751 [2], \oc8051_golden_model_1.n2914 [2]);
  buf(\oc8051_golden_model_1.n2751 [3], \oc8051_golden_model_1.n2914 [3]);
  buf(\oc8051_golden_model_1.n2751 [4], \oc8051_golden_model_1.n2914 [4]);
  buf(\oc8051_golden_model_1.n2751 [5], \oc8051_golden_model_1.n2914 [5]);
  buf(\oc8051_golden_model_1.n2751 [6], \oc8051_golden_model_1.n2914 [6]);
  buf(\oc8051_golden_model_1.n2751 [7], \oc8051_golden_model_1.n2914 [7]);
  buf(\oc8051_golden_model_1.n2752 , \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2753 , \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2754 , \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2755 , \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2756 , \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2757 , \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2758 , \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2759 , \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2766 , \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.n2767 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2767 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2767 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2767 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2767 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2767 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2767 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2782 , \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.n2783 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2783 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2783 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2783 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2783 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2783 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2783 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2815 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2815 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2815 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2815 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2815 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2815 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2815 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2815 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2816 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2816 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2816 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2816 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2816 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2816 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.n2914 [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2836 , \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2837 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2837 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2837 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2837 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2837 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2837 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2837 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2837 [7], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.n2854 [7]);
  buf(\oc8051_golden_model_1.n2853 , \oc8051_golden_model_1.n2854 [0]);
  buf(\oc8051_golden_model_1.n2854 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2854 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2854 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2854 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2854 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2854 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2858 [0], \oc8051_golden_model_1.n2868 );
  buf(\oc8051_golden_model_1.n2858 [1], \oc8051_golden_model_1.n2867 );
  buf(\oc8051_golden_model_1.n2858 [2], \oc8051_golden_model_1.n2866 );
  buf(\oc8051_golden_model_1.n2858 [3], \oc8051_golden_model_1.n2865 );
  buf(\oc8051_golden_model_1.n2858 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2858 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2858 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2858 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2859 [0], \oc8051_golden_model_1.n2860 [4]);
  buf(\oc8051_golden_model_1.n2859 [1], \oc8051_golden_model_1.n2860 [5]);
  buf(\oc8051_golden_model_1.n2859 [2], \oc8051_golden_model_1.n2860 [6]);
  buf(\oc8051_golden_model_1.n2859 [3], \oc8051_golden_model_1.n2860 [7]);
  buf(\oc8051_golden_model_1.n2860 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2860 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2860 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2860 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2861 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2862 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2864 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2875 , \oc8051_golden_model_1.n2876 [0]);
  buf(\oc8051_golden_model_1.n2876 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2876 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2876 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2876 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2876 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2876 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2876 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2894 , \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.n2895 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2895 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2895 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2895 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2895 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2895 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2895 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2896 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2896 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2896 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2896 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2896 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2896 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2896 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2912 , \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.n2913 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2913 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2913 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2913 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2913 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2913 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2913 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.sub_result [0], ABINPUT[27]);
  buf(\oc8051_top_1.sub_result [1], ABINPUT[28]);
  buf(\oc8051_top_1.sub_result [2], ABINPUT[29]);
  buf(\oc8051_top_1.sub_result [3], ABINPUT[30]);
  buf(\oc8051_top_1.sub_result [4], ABINPUT[31]);
  buf(\oc8051_top_1.sub_result [5], ABINPUT[32]);
  buf(\oc8051_top_1.sub_result [6], ABINPUT[33]);
  buf(\oc8051_top_1.sub_result [7], ABINPUT[34]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_top_1.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_top_1.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_top_1.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_top_1.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_top_1.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_top_1.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_top_1.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_top_1.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_top_1.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_top_1.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_top_1.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_top_1.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_top_1.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_top_1.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_top_1.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_top_1.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_top_1.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_top_1.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_top_1.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_top_1.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_top_1.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_top_1.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_top_1.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_top_1.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_top_1.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.desCy , ABINPUT[0]);
  buf(\oc8051_top_1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
